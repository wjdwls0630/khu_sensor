
module converter_i2f ( i_A, i_A_STB, o_A_ACK, o_Z, o_Z_STB, i_Z_ACK, i_CLK, 
        i_RST );
  input [31:0] i_A;
  output [31:0] o_Z;
  input i_A_STB, i_Z_ACK, i_CLK, i_RST;
  output o_A_ACK, o_Z_STB;
  wire   z_s, N53, N117, guard, round_bit, N165, N166, N167, N168, N169, N170,
         N171, N172, N232, n1, n13, n15, n78, n124, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584;
  wire   [2:0] state;
  wire   [30:1] a;
  wire   [31:0] value;
  wire   [7:0] z_e;
  wire   [23:0] z_m;
  wire   [7:0] z_r;
  wire   [31:0] z;

  ivd1_hd U229 ( .A(i_RST), .Y(N232) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n233), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n233), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n233), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n233), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n233), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n233), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n233), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n233), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n233), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n233), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n233), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n233), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n233), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n233), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n233), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n233), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n233), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n233), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n233), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n233), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n233), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n228), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n228), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n228), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n228), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n228), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n233), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n233), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n233), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n233), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n233), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n233), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd z_reg_23_ ( .D(N165), .E(n234), .CK(i_CLK), .Q(z[23]) );
  fd1eqd1_hd z_reg_24_ ( .D(N166), .E(n234), .CK(i_CLK), .Q(z[24]) );
  fd1eqd1_hd z_reg_25_ ( .D(N167), .E(n234), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd z_reg_26_ ( .D(N168), .E(n234), .CK(i_CLK), .Q(z[26]) );
  fd1eqd1_hd z_reg_27_ ( .D(N169), .E(n234), .CK(i_CLK), .Q(z[27]) );
  fd1eqd1_hd z_reg_28_ ( .D(N170), .E(n234), .CK(i_CLK), .Q(z[28]) );
  fd1eqd1_hd z_reg_29_ ( .D(N171), .E(n234), .CK(i_CLK), .Q(z[29]) );
  fd1eqd1_hd z_reg_30_ ( .D(N172), .E(n234), .CK(i_CLK), .Q(z[30]) );
  fd1eqd1_hd z_s_reg ( .D(N117), .E(n15), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd z_reg_31_ ( .D(z_s), .E(n234), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd z_reg_0_ ( .D(z_m[0]), .E(n234), .CK(i_CLK), .Q(z[0]) );
  fd1eqd1_hd z_reg_1_ ( .D(z_m[1]), .E(n227), .CK(i_CLK), .Q(z[1]) );
  fd1eqd1_hd z_reg_2_ ( .D(z_m[2]), .E(n227), .CK(i_CLK), .Q(z[2]) );
  fd1eqd1_hd z_reg_3_ ( .D(z_m[3]), .E(n227), .CK(i_CLK), .Q(z[3]) );
  fd1eqd1_hd z_reg_4_ ( .D(z_m[4]), .E(n227), .CK(i_CLK), .Q(z[4]) );
  fd1eqd1_hd z_reg_5_ ( .D(z_m[5]), .E(n227), .CK(i_CLK), .Q(z[5]) );
  fd1eqd1_hd z_reg_6_ ( .D(z_m[6]), .E(n227), .CK(i_CLK), .Q(z[6]) );
  fd1eqd1_hd z_reg_7_ ( .D(z_m[7]), .E(n234), .CK(i_CLK), .Q(z[7]) );
  fd1eqd1_hd z_reg_8_ ( .D(z_m[8]), .E(n234), .CK(i_CLK), .Q(z[8]) );
  fd1eqd1_hd z_reg_9_ ( .D(z_m[9]), .E(n234), .CK(i_CLK), .Q(z[9]) );
  fd1eqd1_hd z_reg_10_ ( .D(z_m[10]), .E(n234), .CK(i_CLK), .Q(z[10]) );
  fd1eqd1_hd z_reg_11_ ( .D(z_m[11]), .E(n234), .CK(i_CLK), .Q(z[11]) );
  fd1eqd1_hd z_reg_12_ ( .D(z_m[12]), .E(n234), .CK(i_CLK), .Q(z[12]) );
  fd1eqd1_hd z_reg_13_ ( .D(z_m[13]), .E(n234), .CK(i_CLK), .Q(z[13]) );
  fd1eqd1_hd z_reg_14_ ( .D(z_m[14]), .E(n234), .CK(i_CLK), .Q(z[14]) );
  fd1eqd1_hd z_reg_15_ ( .D(z_m[15]), .E(n234), .CK(i_CLK), .Q(z[15]) );
  fd1eqd1_hd z_reg_16_ ( .D(z_m[16]), .E(n234), .CK(i_CLK), .Q(z[16]) );
  fd1eqd1_hd z_reg_17_ ( .D(z_m[17]), .E(n234), .CK(i_CLK), .Q(z[17]) );
  fd1eqd1_hd z_reg_18_ ( .D(z_m[18]), .E(n234), .CK(i_CLK), .Q(z[18]) );
  fd1eqd1_hd z_reg_19_ ( .D(z_m[19]), .E(n234), .CK(i_CLK), .Q(z[19]) );
  fd1eqd1_hd z_reg_20_ ( .D(z_m[20]), .E(n234), .CK(i_CLK), .Q(z[20]) );
  fd1eqd1_hd z_reg_21_ ( .D(z_m[21]), .E(n234), .CK(i_CLK), .Q(z[21]) );
  fd1eqd1_hd z_reg_22_ ( .D(z_m[22]), .E(n234), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd value_reg_0_ ( .D(n221), .CK(i_CLK), .Q(value[0]) );
  fd1qd1_hd value_reg_30_ ( .D(n191), .CK(i_CLK), .Q(value[30]) );
  fd1qd1_hd value_reg_10_ ( .D(n211), .CK(i_CLK), .Q(value[10]) );
  fd1qd1_hd value_reg_31_ ( .D(n190), .CK(i_CLK), .Q(value[31]) );
  fd1qd1_hd z_r_reg_1_ ( .D(n186), .CK(i_CLK), .Q(z_r[1]) );
  fd1qd1_hd z_r_reg_2_ ( .D(n185), .CK(i_CLK), .Q(z_r[2]) );
  fd1qd1_hd z_r_reg_3_ ( .D(n184), .CK(i_CLK), .Q(z_r[3]) );
  fd1qd1_hd value_reg_2_ ( .D(n219), .CK(i_CLK), .Q(value[2]) );
  fd1qd1_hd value_reg_4_ ( .D(n217), .CK(i_CLK), .Q(value[4]) );
  fd1qd1_hd value_reg_6_ ( .D(n215), .CK(i_CLK), .Q(value[6]) );
  fd1qd1_hd value_reg_8_ ( .D(n213), .CK(i_CLK), .Q(value[8]) );
  fd1qd1_hd value_reg_12_ ( .D(n209), .CK(i_CLK), .Q(value[12]) );
  fd1qd1_hd value_reg_14_ ( .D(n207), .CK(i_CLK), .Q(value[14]) );
  fd1qd1_hd value_reg_16_ ( .D(n205), .CK(i_CLK), .Q(value[16]) );
  fd1qd1_hd value_reg_18_ ( .D(n203), .CK(i_CLK), .Q(value[18]) );
  fd1qd1_hd value_reg_20_ ( .D(n201), .CK(i_CLK), .Q(value[20]) );
  fd1qd1_hd value_reg_22_ ( .D(n199), .CK(i_CLK), .Q(value[22]) );
  fd1qd1_hd value_reg_24_ ( .D(n197), .CK(i_CLK), .Q(value[24]) );
  fd1qd1_hd value_reg_26_ ( .D(n195), .CK(i_CLK), .Q(value[26]) );
  fd1qd1_hd value_reg_28_ ( .D(n193), .CK(i_CLK), .Q(value[28]) );
  fd1qd1_hd value_reg_1_ ( .D(n220), .CK(i_CLK), .Q(value[1]) );
  fd1qd1_hd value_reg_3_ ( .D(n218), .CK(i_CLK), .Q(value[3]) );
  fd1qd1_hd value_reg_5_ ( .D(n216), .CK(i_CLK), .Q(value[5]) );
  fd1qd1_hd value_reg_7_ ( .D(n214), .CK(i_CLK), .Q(value[7]) );
  fd1qd1_hd value_reg_9_ ( .D(n212), .CK(i_CLK), .Q(value[9]) );
  fd1qd1_hd value_reg_11_ ( .D(n210), .CK(i_CLK), .Q(value[11]) );
  fd1qd1_hd value_reg_13_ ( .D(n208), .CK(i_CLK), .Q(value[13]) );
  fd1qd1_hd value_reg_15_ ( .D(n206), .CK(i_CLK), .Q(value[15]) );
  fd1qd1_hd value_reg_17_ ( .D(n204), .CK(i_CLK), .Q(value[17]) );
  fd1qd1_hd value_reg_19_ ( .D(n202), .CK(i_CLK), .Q(value[19]) );
  fd1qd1_hd value_reg_21_ ( .D(n200), .CK(i_CLK), .Q(value[21]) );
  fd1qd1_hd value_reg_23_ ( .D(n198), .CK(i_CLK), .Q(value[23]) );
  fd1qd1_hd value_reg_25_ ( .D(n196), .CK(i_CLK), .Q(value[25]) );
  fd1qd1_hd value_reg_27_ ( .D(n194), .CK(i_CLK), .Q(value[27]) );
  fd1qd1_hd value_reg_29_ ( .D(n192), .CK(i_CLK), .Q(value[29]) );
  fd1qd1_hd z_r_reg_6_ ( .D(n188), .CK(i_CLK), .Q(z_r[6]) );
  fd1qd1_hd z_r_reg_0_ ( .D(n187), .CK(i_CLK), .Q(z_r[0]) );
  fd1qd1_hd z_r_reg_7_ ( .D(n181), .CK(i_CLK), .Q(z_r[7]) );
  fd1qd1_hd z_r_reg_4_ ( .D(n183), .CK(i_CLK), .Q(z_r[4]) );
  fd1qd1_hd z_r_reg_5_ ( .D(n182), .CK(i_CLK), .Q(z_r[5]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n189), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_e_reg_4_ ( .D(n150), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n157), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n155), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n156), .CK(i_CLK), .Q(z_e[5]) );
  fd1eqd1_hd sticky_reg ( .D(n78), .E(n13), .CK(i_CLK), .Q(n1) );
  fd1qd1_hd z_e_reg_0_ ( .D(n154), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd o_A_ACK_reg ( .D(n222), .CK(i_CLK), .Q(o_A_ACK) );
  fd1qd1_hd z_e_reg_3_ ( .D(n151), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n153), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n152), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n163), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n162), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n158), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd guard_reg ( .D(z_r[7]), .E(n13), .CK(i_CLK), .Q(guard) );
  fd1eqd1_hd round_bit_reg ( .D(z_r[6]), .E(n13), .CK(i_CLK), .Q(round_bit) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n124), .CK(i_CLK), .Q(N117) );
  fd1qd1_hd z_m_reg_9_ ( .D(n171), .CK(i_CLK), .Q(z_m[9]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n124), .CK(i_CLK), .Q(a[30]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n226), .CK(i_CLK), .Q(z_m[23]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n124), .CK(i_CLK), .Q(a[29]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n175), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n167), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n170), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n172), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n168), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n164), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n160), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n173), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n169), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n165), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n161), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n174), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n166), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n159), .CK(i_CLK), .Q(z_m[21]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n124), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n124), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n124), .CK(i_CLK), .Q(a[24]) );
  fd1qd1_hd state_reg_2_ ( .D(n225), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_0_ ( .D(n224), .CK(i_CLK), .Q(state[0]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n124), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n124), .CK(i_CLK), .Q(a[25]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n180), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd state_reg_1_ ( .D(n223), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n176), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n177), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n179), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n178), .CK(i_CLK), .Q(z_m[2]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n124), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n124), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n124), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n124), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n124), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n124), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n124), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n124), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n124), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n124), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n124), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n124), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n124), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n124), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n124), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n124), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n124), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n124), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n124), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n124), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n124), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n124), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n124), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n124), .CK(i_CLK), .Q(N53) );
  clknd2d1_hd U231 ( .A(z_m[2]), .B(z_m[1]), .Y(n531) );
  clknd2d1_hd U232 ( .A(z_m[14]), .B(z_m[13]), .Y(n532) );
  clknd2d1_hd U233 ( .A(n530), .B(n502), .Y(n244) );
  clknd2d1_hd U234 ( .A(n526), .B(n459), .Y(n469) );
  clknd2d1_hd U235 ( .A(n527), .B(n419), .Y(n429) );
  clknd2d1_hd U236 ( .A(n525), .B(n439), .Y(n449) );
  clknd2d1_hd U237 ( .A(n529), .B(n479), .Y(n490) );
  clknd2d1_hd U238 ( .A(z_m[18]), .B(z_m[17]), .Y(n540) );
  clknd2d1_hd U239 ( .A(n407), .B(n255), .Y(n541) );
  clknd2d1_hd U240 ( .A(n570), .B(guard), .Y(n241) );
  clknd2d1_hd U241 ( .A(z_m[6]), .B(z_m[5]), .Y(n539) );
  clknd2d1_hd U242 ( .A(z_e[4]), .B(n576), .Y(n545) );
  clknd2d1_hd U243 ( .A(n520), .B(n265), .Y(n559) );
  clknd2d1_hd U244 ( .A(n501), .B(n411), .Y(n414) );
  clknd2d1_hd U245 ( .A(n507), .B(n419), .Y(n424) );
  clknd2d1_hd U246 ( .A(n507), .B(n534), .Y(n411) );
  clknd2d1_hd U247 ( .A(n252), .B(n258), .Y(n254) );
  clknd2d1_hd U248 ( .A(n15), .B(n259), .Y(n255) );
  clknd2d1_hd U249 ( .A(n507), .B(n502), .Y(n509) );
  clknd2d1_hd U250 ( .A(n507), .B(n479), .Y(n484) );
  clknd2d1_hd U251 ( .A(n507), .B(n459), .Y(n464) );
  clknd2d1_hd U252 ( .A(n507), .B(n439), .Y(n444) );
  clknd2d1_hd U253 ( .A(z_m[21]), .B(n514), .Y(n524) );
  clknd2d1_hd U254 ( .A(n258), .B(n250), .Y(n564) );
  clknd2d1_hd U255 ( .A(n526), .B(n525), .Y(n538) );
  clknd2d1_hd U256 ( .A(n565), .B(z_e[2]), .Y(n572) );
  clknd2d1_hd U257 ( .A(state[1]), .B(n243), .Y(n544) );
  clknd2d1_hd U258 ( .A(z_e[5]), .B(n551), .Y(n555) );
  clknd2d1_hd U259 ( .A(n15), .B(n563), .Y(n557) );
  clknd2d1_hd U260 ( .A(n570), .B(n563), .Y(n583) );
  clknd2d1_hd U261 ( .A(n571), .B(n573), .Y(n577) );
  clknd2d1_hd U262 ( .A(n563), .B(n559), .Y(n581) );
  clknd2d1_hd U263 ( .A(n375), .B(n378), .Y(n383) );
  clknd2d1_hd U264 ( .A(n366), .B(n369), .Y(n373) );
  clknd2d1_hd U265 ( .A(n358), .B(n361), .Y(n365) );
  clknd2d1_hd U266 ( .A(n350), .B(n353), .Y(n357) );
  clknd2d1_hd U267 ( .A(n342), .B(n345), .Y(n349) );
  clknd2d1_hd U268 ( .A(n334), .B(n337), .Y(n341) );
  clknd2d1_hd U269 ( .A(n326), .B(n329), .Y(n333) );
  clknd2d1_hd U270 ( .A(n318), .B(n321), .Y(n325) );
  clknd2d1_hd U271 ( .A(n310), .B(n313), .Y(n317) );
  clknd2d1_hd U272 ( .A(n302), .B(n305), .Y(n309) );
  clknd2d1_hd U273 ( .A(n294), .B(n297), .Y(n301) );
  clknd2d1_hd U274 ( .A(n286), .B(n289), .Y(n293) );
  clknd2d1_hd U275 ( .A(n278), .B(n281), .Y(n285) );
  clknd2d1_hd U276 ( .A(n270), .B(n273), .Y(n277) );
  clknd2d1_hd U277 ( .A(n261), .B(n243), .Y(n265) );
  clknd2d1_hd U278 ( .A(n239), .B(n554), .Y(n240) );
  clknd2d1_hd U279 ( .A(n237), .B(n575), .Y(n238) );
  clknd2d1_hd U280 ( .A(n235), .B(n562), .Y(n236) );
  clknd2d1_hd U281 ( .A(n413), .B(n412), .Y(n179) );
  clknd2d1_hd U282 ( .A(z_m[3]), .B(n422), .Y(n420) );
  clknd2d1_hd U283 ( .A(n256), .B(n260), .Y(n257) );
  clknd2d1_hd U284 ( .A(n255), .B(n544), .Y(n251) );
  clknd2d1_hd U285 ( .A(n514), .B(n517), .Y(n515) );
  clknd2d1_hd U286 ( .A(z_m[19]), .B(n505), .Y(n503) );
  clknd2d1_hd U287 ( .A(z_m[15]), .B(n482), .Y(n480) );
  clknd2d1_hd U288 ( .A(z_m[11]), .B(n462), .Y(n460) );
  clknd2d1_hd U289 ( .A(z_m[7]), .B(n442), .Y(n440) );
  clknd2d1_hd U290 ( .A(n473), .B(n477), .Y(n470) );
  clknd2d1_hd U291 ( .A(n433), .B(n437), .Y(n430) );
  clknd2d1_hd U292 ( .A(n453), .B(n457), .Y(n450) );
  clknd2d1_hd U293 ( .A(z_m[22]), .B(n521), .Y(n522) );
  clknd2d1_hd U294 ( .A(n494), .B(n499), .Y(n491) );
  clknd2d1_hd U295 ( .A(n565), .B(n562), .Y(n568) );
  clknd2d1_hd U296 ( .A(n576), .B(n575), .Y(n584) );
  clknd2d1_hd U297 ( .A(n578), .B(n577), .Y(n580) );
  clknd2d1_hd U298 ( .A(N53), .B(n384), .Y(n269) );
  clknd2d1_hd U299 ( .A(a[30]), .B(n388), .Y(n387) );
  nid2_hd U300 ( .A(n228), .Y(n233) );
  xo2d1_hd U301 ( .A(z_e[7]), .B(n240), .Y(N172) );
  ivd3_hd U302 ( .A(n248), .Y(n124) );
  scg10d1_hd U303 ( .A(n390), .B(N53), .C(value[0]), .D(n266), .Y(n221) );
  ivd2_hd U304 ( .A(n266), .Y(n390) );
  scg2d1_hd U305 ( .A(n232), .B(value[0]), .C(n407), .D(z_r[0]), .Y(n187) );
  or2d1_hd U306 ( .A(n261), .B(n254), .Y(n520) );
  or2d1_hd U307 ( .A(n565), .B(n235), .Y(N166) );
  ad4d1_hd U308 ( .A(n530), .B(n529), .C(n528), .D(n527), .Y(n536) );
  nr2d2_hd U309 ( .A(n544), .B(n489), .Y(n519) );
  nr2ad1_hd U310 ( .A(n489), .B(n564), .Y(n507) );
  ivd1_hd U311 ( .A(n380), .Y(n374) );
  ivd1_hd U312 ( .A(n507), .Y(n496) );
  nr2d1_hd U313 ( .A(n543), .B(n541), .Y(n489) );
  nd2d1_hd U314 ( .A(n266), .B(n385), .Y(n380) );
  nr2d1_hd U315 ( .A(n259), .B(n265), .Y(n266) );
  ivd1_hd U316 ( .A(n489), .Y(n501) );
  ivd1_hd U317 ( .A(n569), .Y(n563) );
  nr2d1_hd U318 ( .A(N117), .B(n391), .Y(n259) );
  nd2bd1_hd U319 ( .AN(a[30]), .B(n386), .Y(n391) );
  nr2d1_hd U320 ( .A(a[29]), .B(n383), .Y(n386) );
  nr2d1_hd U321 ( .A(a[27]), .B(n373), .Y(n375) );
  nr2d1_hd U322 ( .A(a[25]), .B(n365), .Y(n366) );
  nr2d1_hd U323 ( .A(a[23]), .B(n357), .Y(n358) );
  nr2d1_hd U324 ( .A(a[21]), .B(n349), .Y(n350) );
  nr2d1_hd U325 ( .A(a[19]), .B(n341), .Y(n342) );
  nr2d1_hd U326 ( .A(a[17]), .B(n333), .Y(n334) );
  nr2d1_hd U327 ( .A(a[15]), .B(n325), .Y(n326) );
  nr2d1_hd U328 ( .A(a[13]), .B(n317), .Y(n318) );
  nr2d1_hd U329 ( .A(a[11]), .B(n309), .Y(n310) );
  nr2d1_hd U330 ( .A(a[9]), .B(n301), .Y(n302) );
  nr2d1_hd U331 ( .A(a[7]), .B(n293), .Y(n294) );
  nr2d1_hd U332 ( .A(a[5]), .B(n285), .Y(n286) );
  nr2d1_hd U333 ( .A(a[3]), .B(n277), .Y(n278) );
  ivd1_hd U334 ( .A(a[2]), .Y(n273) );
  nr2d1_hd U335 ( .A(a[1]), .B(N53), .Y(n270) );
  ivd1_hd U336 ( .A(n564), .Y(n570) );
  nid2_hd U337 ( .A(n384), .Y(n231) );
  nr2d1_hd U338 ( .A(n265), .B(n385), .Y(n384) );
  ivd1_hd U339 ( .A(n519), .Y(n508) );
  nr2d1_hd U340 ( .A(n544), .B(n569), .Y(n579) );
  ao21d1_hd U341 ( .A(n543), .B(n542), .C(n541), .Y(n569) );
  ivd1_hd U342 ( .A(a[6]), .Y(n289) );
  ivd1_hd U343 ( .A(a[4]), .Y(n281) );
  ivd1_hd U344 ( .A(n401), .Y(n407) );
  ivd1_hd U345 ( .A(n409), .Y(n399) );
  nid2_hd U346 ( .A(n227), .Y(n234) );
  nr2bd1_hd U347 ( .AN(n250), .B(n258), .Y(n227) );
  ivd2_hd U348 ( .A(n231), .Y(n230) );
  ivd1_hd U349 ( .A(N117), .Y(n385) );
  ivd2_hd U350 ( .A(n520), .Y(n232) );
  nr2bd1_hd U351 ( .AN(n528), .B(n449), .Y(n459) );
  scg17d1_hd U352 ( .A(n579), .B(N168), .C(n574), .D(n581), .Y(n151) );
  nr2bd1_hd U353 ( .AN(z_e[1]), .B(N165), .Y(n565) );
  ivd1_hd U354 ( .A(a[28]), .Y(n378) );
  ivd1_hd U355 ( .A(a[26]), .Y(n369) );
  ivd1_hd U356 ( .A(a[24]), .Y(n361) );
  ivd1_hd U357 ( .A(a[22]), .Y(n353) );
  ivd1_hd U358 ( .A(a[20]), .Y(n345) );
  ivd1_hd U359 ( .A(a[18]), .Y(n337) );
  ivd1_hd U360 ( .A(a[16]), .Y(n329) );
  ivd1_hd U361 ( .A(a[14]), .Y(n321) );
  ivd1_hd U362 ( .A(a[12]), .Y(n313) );
  ivd1_hd U363 ( .A(a[10]), .Y(n305) );
  ivd1_hd U364 ( .A(a[8]), .Y(n297) );
  ivd1_hd U365 ( .A(n265), .Y(n15) );
  ivd1_hd U366 ( .A(state[1]), .Y(n261) );
  ao21d1_hd U367 ( .A(n1), .B(n242), .C(n241), .Y(n543) );
  ivd1_hd U368 ( .A(state[2]), .Y(n252) );
  ivd1_hd U369 ( .A(state[0]), .Y(n258) );
  ivd1_hd U370 ( .A(z_r[2]), .Y(n403) );
  ivd1_hd U371 ( .A(z_r[3]), .Y(n402) );
  ivd1_hd U372 ( .A(z_r[1]), .Y(n404) );
  ivd1_hd U373 ( .A(z_r[5]), .Y(n405) );
  nd3d1_hd U374 ( .A(n264), .B(i_A_STB), .C(o_A_ACK), .Y(n248) );
  nr3d1_hd U375 ( .A(state[0]), .B(n252), .C(n261), .Y(n228) );
  ivd1_hd U376 ( .A(z_m[21]), .Y(n517) );
  scg14d1_hd U377 ( .A(value[30]), .B(n390), .C(n389), .Y(n191) );
  ivd1_hd U378 ( .A(z_m[13]), .Y(n477) );
  ivd1_hd U379 ( .A(z_m[17]), .Y(n499) );
  ivd1_hd U380 ( .A(z_m[5]), .Y(n437) );
  scg6d1_hd U381 ( .A(z_e[5]), .B(n238), .C(n239), .Y(N170) );
  scg6d1_hd U382 ( .A(z_e[3]), .B(n236), .C(n237), .Y(N168) );
  ivd1_hd U383 ( .A(z_e[0]), .Y(N165) );
  ivd1_hd U384 ( .A(z_e[6]), .Y(n554) );
  ivd1_hd U385 ( .A(z_e[4]), .Y(n575) );
  ivd1_hd U386 ( .A(z_e[2]), .Y(n562) );
  ivd1_hd U387 ( .A(z_m[23]), .Y(n533) );
  ivd1_hd U388 ( .A(z_m[0]), .Y(n534) );
  ivd1_hd U389 ( .A(z_m[4]), .Y(n427) );
  ivd1_hd U390 ( .A(z_m[9]), .Y(n457) );
  ivd1_hd U391 ( .A(z_m[16]), .Y(n487) );
  ivd1_hd U392 ( .A(z_m[20]), .Y(n512) );
  ivd1_hd U393 ( .A(z_m[8]), .Y(n447) );
  ivd1_hd U394 ( .A(z_m[12]), .Y(n467) );
  nr2d1_hd U395 ( .A(n258), .B(state[2]), .Y(n243) );
  nr2d1_hd U396 ( .A(n544), .B(n407), .Y(n409) );
  nr2d1_hd U397 ( .A(state[1]), .B(n254), .Y(n264) );
  nr2d1_hd U398 ( .A(z_e[3]), .B(n236), .Y(n237) );
  nr2d1_hd U399 ( .A(z_e[0]), .B(z_e[1]), .Y(n235) );
  oa21d1_hd U400 ( .A(n544), .B(z_m[23]), .C(n520), .Y(n401) );
  nr2d1_hd U401 ( .A(n252), .B(state[1]), .Y(n250) );
  oa21d1_hd U402 ( .A(n235), .B(n562), .C(n236), .Y(N167) );
  oa21d1_hd U403 ( .A(n237), .B(n575), .C(n238), .Y(N169) );
  nr2d1_hd U404 ( .A(z_e[5]), .B(n238), .Y(n239) );
  oa21d1_hd U405 ( .A(n239), .B(n554), .C(n240), .Y(N171) );
  nr2d1_hd U406 ( .A(z_m[0]), .B(round_bit), .Y(n242) );
  ivd1_hd U407 ( .A(z_m[19]), .Y(n506) );
  nr2d1_hd U408 ( .A(n512), .B(n506), .Y(n530) );
  ivd1_hd U409 ( .A(z_m[15]), .Y(n483) );
  nr2d1_hd U410 ( .A(n487), .B(n483), .Y(n529) );
  ivd1_hd U411 ( .A(z_m[11]), .Y(n463) );
  nr2d1_hd U412 ( .A(n467), .B(n463), .Y(n526) );
  ivd1_hd U413 ( .A(z_m[10]), .Y(n452) );
  nr2d1_hd U414 ( .A(n452), .B(n457), .Y(n528) );
  ivd1_hd U415 ( .A(z_m[7]), .Y(n443) );
  nr2d1_hd U416 ( .A(n447), .B(n443), .Y(n525) );
  ivd1_hd U417 ( .A(z_m[3]), .Y(n423) );
  nr2d1_hd U418 ( .A(n427), .B(n423), .Y(n527) );
  nr2d1_hd U419 ( .A(n534), .B(n531), .Y(n419) );
  nr2d1_hd U420 ( .A(n539), .B(n429), .Y(n439) );
  nr2d1_hd U421 ( .A(n532), .B(n469), .Y(n479) );
  nr2d1_hd U422 ( .A(n540), .B(n490), .Y(n502) );
  ao21d1_hd U423 ( .A(n507), .B(n244), .C(n489), .Y(n518) );
  oa21d1_hd U424 ( .A(z_m[21]), .B(n496), .C(n518), .Y(n521) );
  scg20d1_hd U425 ( .A(n496), .B(z_m[22]), .C(n521), .Y(n247) );
  nr2d1_hd U426 ( .A(n496), .B(n244), .Y(n514) );
  oa21d1_hd U427 ( .A(z_m[23]), .B(n524), .C(n508), .Y(n245) );
  ao22d1_hd U428 ( .A(n232), .B(value[31]), .C(z_m[22]), .D(n245), .Y(n246) );
  oa21d1_hd U429 ( .A(n247), .B(n533), .C(n246), .Y(n226) );
  nr2d1_hd U430 ( .A(n544), .B(n533), .Y(n13) );
  nr4d1_hd U431 ( .A(n250), .B(n13), .C(i_RST), .D(n559), .Y(n249) );
  nd3d1_hd U432 ( .A(n233), .B(i_Z_ACK), .C(o_Z_STB), .Y(n392) );
  nd3d1_hd U433 ( .A(n249), .B(n392), .C(n248), .Y(n260) );
  ao21d1_hd U434 ( .A(n251), .B(n260), .C(n250), .Y(n253) );
  ivd1_hd U435 ( .A(N232), .Y(n262) );
  oa22d1_hd U436 ( .A(n253), .B(n262), .C(n252), .D(n260), .Y(n225) );
  nd3d1_hd U437 ( .A(n564), .B(n255), .C(n254), .Y(n256) );
  oa22d1_hd U438 ( .A(n258), .B(n260), .C(n262), .D(n257), .Y(n224) );
  nr3d1_hd U439 ( .A(n232), .B(n266), .C(n234), .Y(n263) );
  oa22d1_hd U440 ( .A(n263), .B(n262), .C(n261), .D(n260), .Y(n223) );
  scg21d1_hd U441 ( .A(n264), .B(o_A_ACK), .C(i_RST), .D(n124), .Y(n222) );
  oa21d1_hd U442 ( .A(N53), .B(n230), .C(n380), .Y(n267) );
  ao22d1_hd U443 ( .A(a[1]), .B(n267), .C(value[1]), .D(n390), .Y(n268) );
  oa21d1_hd U444 ( .A(a[1]), .B(n269), .C(n268), .Y(n220) );
  ao21d1_hd U445 ( .A(n270), .B(n231), .C(n374), .Y(n274) );
  nr2d1_hd U446 ( .A(n270), .B(n230), .Y(n271) );
  ao22d1_hd U447 ( .A(value[2]), .B(n390), .C(n271), .D(n273), .Y(n272) );
  oa21d1_hd U448 ( .A(n274), .B(n273), .C(n272), .Y(n219) );
  oa21d1_hd U449 ( .A(n277), .B(n230), .C(n380), .Y(n275) );
  ao22d1_hd U450 ( .A(a[3]), .B(n275), .C(value[3]), .D(n390), .Y(n276) );
  scg22d1_hd U451 ( .A(n231), .B(n277), .C(a[3]), .D(n276), .Y(n218) );
  ao21d1_hd U452 ( .A(n278), .B(n231), .C(n374), .Y(n282) );
  nr2d1_hd U453 ( .A(n278), .B(n230), .Y(n279) );
  ao22d1_hd U454 ( .A(value[4]), .B(n390), .C(n279), .D(n281), .Y(n280) );
  oa21d1_hd U455 ( .A(n282), .B(n281), .C(n280), .Y(n217) );
  oa21d1_hd U456 ( .A(n285), .B(n230), .C(n380), .Y(n283) );
  ao22d1_hd U457 ( .A(a[5]), .B(n283), .C(value[5]), .D(n390), .Y(n284) );
  scg22d1_hd U458 ( .A(n231), .B(n285), .C(a[5]), .D(n284), .Y(n216) );
  ao21d1_hd U459 ( .A(n286), .B(n231), .C(n374), .Y(n290) );
  nr2d1_hd U460 ( .A(n286), .B(n230), .Y(n287) );
  ao22d1_hd U461 ( .A(value[6]), .B(n390), .C(n287), .D(n289), .Y(n288) );
  oa21d1_hd U462 ( .A(n290), .B(n289), .C(n288), .Y(n215) );
  oa21d1_hd U463 ( .A(n293), .B(n230), .C(n380), .Y(n291) );
  ao22d1_hd U464 ( .A(a[7]), .B(n291), .C(value[7]), .D(n390), .Y(n292) );
  scg22d1_hd U465 ( .A(n231), .B(n293), .C(a[7]), .D(n292), .Y(n214) );
  ao21d1_hd U466 ( .A(n294), .B(n231), .C(n374), .Y(n298) );
  nr2d1_hd U467 ( .A(n294), .B(n230), .Y(n295) );
  ao22d1_hd U468 ( .A(value[8]), .B(n390), .C(n295), .D(n297), .Y(n296) );
  oa21d1_hd U469 ( .A(n298), .B(n297), .C(n296), .Y(n213) );
  oa21d1_hd U470 ( .A(n301), .B(n230), .C(n380), .Y(n299) );
  ao22d1_hd U471 ( .A(a[9]), .B(n299), .C(value[9]), .D(n390), .Y(n300) );
  scg22d1_hd U472 ( .A(n231), .B(n301), .C(a[9]), .D(n300), .Y(n212) );
  ao21d1_hd U473 ( .A(n302), .B(n384), .C(n374), .Y(n306) );
  nr2d1_hd U474 ( .A(n302), .B(n230), .Y(n303) );
  ao22d1_hd U475 ( .A(value[10]), .B(n390), .C(n303), .D(n305), .Y(n304) );
  oa21d1_hd U476 ( .A(n306), .B(n305), .C(n304), .Y(n211) );
  oa21d1_hd U477 ( .A(n309), .B(n230), .C(n380), .Y(n307) );
  ao22d1_hd U478 ( .A(a[11]), .B(n307), .C(value[11]), .D(n390), .Y(n308) );
  scg22d1_hd U479 ( .A(n231), .B(n309), .C(a[11]), .D(n308), .Y(n210) );
  ao21d1_hd U480 ( .A(n310), .B(n384), .C(n374), .Y(n314) );
  nr2d1_hd U481 ( .A(n310), .B(n230), .Y(n311) );
  ao22d1_hd U482 ( .A(value[12]), .B(n390), .C(n311), .D(n313), .Y(n312) );
  oa21d1_hd U483 ( .A(n314), .B(n313), .C(n312), .Y(n209) );
  oa21d1_hd U484 ( .A(n317), .B(n230), .C(n380), .Y(n315) );
  ao22d1_hd U485 ( .A(a[13]), .B(n315), .C(value[13]), .D(n390), .Y(n316) );
  scg22d1_hd U486 ( .A(n231), .B(n317), .C(a[13]), .D(n316), .Y(n208) );
  ao21d1_hd U487 ( .A(n318), .B(n384), .C(n374), .Y(n322) );
  nr2d1_hd U488 ( .A(n318), .B(n230), .Y(n319) );
  ao22d1_hd U489 ( .A(value[14]), .B(n390), .C(n319), .D(n321), .Y(n320) );
  oa21d1_hd U490 ( .A(n322), .B(n321), .C(n320), .Y(n207) );
  oa21d1_hd U491 ( .A(n325), .B(n230), .C(n380), .Y(n323) );
  ao22d1_hd U492 ( .A(a[15]), .B(n323), .C(value[15]), .D(n390), .Y(n324) );
  scg22d1_hd U493 ( .A(n231), .B(n325), .C(a[15]), .D(n324), .Y(n206) );
  ao21d1_hd U494 ( .A(n326), .B(n384), .C(n374), .Y(n330) );
  nr2d1_hd U495 ( .A(n326), .B(n230), .Y(n327) );
  ao22d1_hd U496 ( .A(value[16]), .B(n390), .C(n327), .D(n329), .Y(n328) );
  oa21d1_hd U497 ( .A(n330), .B(n329), .C(n328), .Y(n205) );
  oa21d1_hd U498 ( .A(n333), .B(n230), .C(n380), .Y(n331) );
  ao22d1_hd U499 ( .A(a[17]), .B(n331), .C(value[17]), .D(n390), .Y(n332) );
  scg22d1_hd U500 ( .A(n231), .B(n333), .C(a[17]), .D(n332), .Y(n204) );
  ao21d1_hd U501 ( .A(n334), .B(n231), .C(n374), .Y(n338) );
  nr2d1_hd U502 ( .A(n334), .B(n230), .Y(n335) );
  ao22d1_hd U503 ( .A(value[18]), .B(n390), .C(n335), .D(n337), .Y(n336) );
  oa21d1_hd U504 ( .A(n338), .B(n337), .C(n336), .Y(n203) );
  oa21d1_hd U505 ( .A(n341), .B(n230), .C(n380), .Y(n339) );
  ao22d1_hd U506 ( .A(a[19]), .B(n339), .C(value[19]), .D(n390), .Y(n340) );
  scg22d1_hd U507 ( .A(n231), .B(n341), .C(a[19]), .D(n340), .Y(n202) );
  ao21d1_hd U508 ( .A(n342), .B(n231), .C(n374), .Y(n346) );
  nr2d1_hd U509 ( .A(n342), .B(n230), .Y(n343) );
  ao22d1_hd U510 ( .A(value[20]), .B(n390), .C(n343), .D(n345), .Y(n344) );
  oa21d1_hd U511 ( .A(n346), .B(n345), .C(n344), .Y(n201) );
  oa21d1_hd U512 ( .A(n349), .B(n230), .C(n380), .Y(n347) );
  ao22d1_hd U513 ( .A(a[21]), .B(n347), .C(value[21]), .D(n390), .Y(n348) );
  scg22d1_hd U514 ( .A(n231), .B(n349), .C(a[21]), .D(n348), .Y(n200) );
  ao21d1_hd U515 ( .A(n350), .B(n384), .C(n374), .Y(n354) );
  nr2d1_hd U516 ( .A(n350), .B(n230), .Y(n351) );
  ao22d1_hd U517 ( .A(value[22]), .B(n390), .C(n351), .D(n353), .Y(n352) );
  oa21d1_hd U518 ( .A(n354), .B(n353), .C(n352), .Y(n199) );
  oa21d1_hd U519 ( .A(n357), .B(n230), .C(n380), .Y(n355) );
  ao22d1_hd U520 ( .A(a[23]), .B(n355), .C(value[23]), .D(n390), .Y(n356) );
  scg22d1_hd U521 ( .A(n231), .B(n357), .C(a[23]), .D(n356), .Y(n198) );
  ao21d1_hd U522 ( .A(n358), .B(n384), .C(n374), .Y(n362) );
  nr2d1_hd U523 ( .A(n358), .B(n230), .Y(n359) );
  ao22d1_hd U524 ( .A(value[24]), .B(n390), .C(n359), .D(n361), .Y(n360) );
  oa21d1_hd U525 ( .A(n362), .B(n361), .C(n360), .Y(n197) );
  oa21d1_hd U526 ( .A(n365), .B(n230), .C(n380), .Y(n363) );
  ao22d1_hd U527 ( .A(a[25]), .B(n363), .C(value[25]), .D(n390), .Y(n364) );
  scg22d1_hd U528 ( .A(n231), .B(n365), .C(a[25]), .D(n364), .Y(n196) );
  ao21d1_hd U529 ( .A(n366), .B(n384), .C(n374), .Y(n370) );
  nr2d1_hd U530 ( .A(n366), .B(n230), .Y(n367) );
  ao22d1_hd U531 ( .A(value[26]), .B(n390), .C(n367), .D(n369), .Y(n368) );
  oa21d1_hd U532 ( .A(n370), .B(n369), .C(n368), .Y(n195) );
  oa21d1_hd U533 ( .A(n373), .B(n230), .C(n380), .Y(n371) );
  ao22d1_hd U534 ( .A(a[27]), .B(n371), .C(value[27]), .D(n390), .Y(n372) );
  scg22d1_hd U535 ( .A(n231), .B(n373), .C(a[27]), .D(n372), .Y(n194) );
  ao21d1_hd U536 ( .A(n375), .B(n231), .C(n374), .Y(n379) );
  nr2d1_hd U537 ( .A(n375), .B(n230), .Y(n376) );
  ao22d1_hd U538 ( .A(value[28]), .B(n390), .C(n376), .D(n378), .Y(n377) );
  oa21d1_hd U539 ( .A(n379), .B(n378), .C(n377), .Y(n193) );
  oa21d1_hd U540 ( .A(n383), .B(n230), .C(n380), .Y(n381) );
  ao22d1_hd U541 ( .A(a[29]), .B(n381), .C(value[29]), .D(n390), .Y(n382) );
  scg22d1_hd U542 ( .A(n231), .B(n383), .C(a[29]), .D(n382), .Y(n192) );
  nr2d1_hd U543 ( .A(n386), .B(n385), .Y(n388) );
  oa211d1_hd U544 ( .A(a[30]), .B(n388), .C(n15), .D(n387), .Y(n389) );
  oa22ad1_hd U545 ( .A(n391), .B(n230), .C(n390), .D(value[31]), .Y(n190) );
  ivd1_hd U546 ( .A(n392), .Y(n393) );
  scg21d1_hd U547 ( .A(n233), .B(o_Z_STB), .C(i_RST), .D(n393), .Y(n189) );
  ao22d1_hd U548 ( .A(n232), .B(value[6]), .C(n407), .D(z_r[6]), .Y(n394) );
  oa21d1_hd U549 ( .A(n399), .B(n405), .C(n394), .Y(n188) );
  ao22d1_hd U550 ( .A(n232), .B(value[1]), .C(n407), .D(z_r[1]), .Y(n395) );
  scg14d1_hd U551 ( .A(n409), .B(z_r[0]), .C(n395), .Y(n186) );
  ao22d1_hd U552 ( .A(n232), .B(value[2]), .C(n407), .D(z_r[2]), .Y(n396) );
  oa21d1_hd U553 ( .A(n399), .B(n404), .C(n396), .Y(n185) );
  ao22d1_hd U554 ( .A(n232), .B(value[3]), .C(n407), .D(z_r[3]), .Y(n397) );
  oa21d1_hd U555 ( .A(n399), .B(n403), .C(n397), .Y(n184) );
  ao22d1_hd U556 ( .A(n232), .B(value[4]), .C(n407), .D(z_r[4]), .Y(n398) );
  oa21d1_hd U557 ( .A(n399), .B(n402), .C(n398), .Y(n183) );
  ao22d1_hd U558 ( .A(n232), .B(value[5]), .C(n409), .D(z_r[4]), .Y(n400) );
  oa21d1_hd U559 ( .A(n401), .B(n405), .C(n400), .Y(n182) );
  nd4d1_hd U560 ( .A(n405), .B(n404), .C(n403), .D(n402), .Y(n406) );
  nr3d1_hd U561 ( .A(z_r[0]), .B(z_r[4]), .C(n406), .Y(n78) );
  ao22d1_hd U562 ( .A(n232), .B(value[7]), .C(n407), .D(z_r[7]), .Y(n408) );
  scg14d1_hd U563 ( .A(n409), .B(z_r[6]), .C(n408), .Y(n181) );
  ao22d1_hd U564 ( .A(n232), .B(value[8]), .C(n519), .D(z_r[7]), .Y(n410) );
  oa211d1_hd U565 ( .A(n501), .B(n534), .C(n410), .D(n411), .Y(n180) );
  ao22d1_hd U566 ( .A(n232), .B(value[9]), .C(z_m[1]), .D(n414), .Y(n413) );
  nr2d1_hd U567 ( .A(z_m[1]), .B(n496), .Y(n415) );
  oa21d1_hd U568 ( .A(n519), .B(n415), .C(z_m[0]), .Y(n412) );
  oa21d1_hd U569 ( .A(n415), .B(n414), .C(z_m[2]), .Y(n418) );
  nr3d1_hd U570 ( .A(z_m[2]), .B(n496), .C(n534), .Y(n416) );
  oa21d1_hd U571 ( .A(n519), .B(n416), .C(z_m[1]), .Y(n417) );
  scg15d1_hd U572 ( .A(n232), .B(value[10]), .C(n418), .D(n417), .Y(n178) );
  ao22d1_hd U573 ( .A(n232), .B(value[11]), .C(n519), .D(z_m[2]), .Y(n421) );
  oa21d1_hd U574 ( .A(n419), .B(n564), .C(n501), .Y(n422) );
  oa211d1_hd U575 ( .A(z_m[3]), .B(n424), .C(n421), .D(n420), .Y(n177) );
  ao21d1_hd U576 ( .A(n507), .B(n423), .C(n422), .Y(n428) );
  oa21d1_hd U577 ( .A(z_m[4]), .B(n424), .C(n508), .Y(n425) );
  ao22d1_hd U578 ( .A(n232), .B(value[12]), .C(z_m[3]), .D(n425), .Y(n426) );
  oa21d1_hd U579 ( .A(n428), .B(n427), .C(n426), .Y(n176) );
  ao21d1_hd U580 ( .A(n570), .B(n429), .C(n489), .Y(n434) );
  ao22d1_hd U581 ( .A(n232), .B(value[13]), .C(n519), .D(z_m[4]), .Y(n431) );
  nr2d1_hd U582 ( .A(n496), .B(n429), .Y(n433) );
  oa211d1_hd U583 ( .A(n434), .B(n437), .C(n431), .D(n430), .Y(n175) );
  ivd1_hd U584 ( .A(z_m[6]), .Y(n432) );
  ao21d1_hd U585 ( .A(n433), .B(n432), .C(n519), .Y(n438) );
  oa21d1_hd U586 ( .A(z_m[5]), .B(n496), .C(n434), .Y(n435) );
  ao22d1_hd U587 ( .A(n232), .B(value[14]), .C(z_m[6]), .D(n435), .Y(n436) );
  oa21d1_hd U588 ( .A(n438), .B(n437), .C(n436), .Y(n174) );
  ao22d1_hd U589 ( .A(n232), .B(value[15]), .C(n519), .D(z_m[6]), .Y(n441) );
  oa21d1_hd U590 ( .A(n439), .B(n564), .C(n501), .Y(n442) );
  oa211d1_hd U591 ( .A(z_m[7]), .B(n444), .C(n441), .D(n440), .Y(n173) );
  ao21d1_hd U592 ( .A(n507), .B(n443), .C(n442), .Y(n448) );
  oa21d1_hd U593 ( .A(z_m[8]), .B(n444), .C(n508), .Y(n445) );
  ao22d1_hd U594 ( .A(n232), .B(value[16]), .C(z_m[7]), .D(n445), .Y(n446) );
  oa21d1_hd U595 ( .A(n448), .B(n447), .C(n446), .Y(n172) );
  ao21d1_hd U596 ( .A(n570), .B(n449), .C(n489), .Y(n454) );
  ao22d1_hd U597 ( .A(n232), .B(value[17]), .C(n519), .D(z_m[8]), .Y(n451) );
  nr2d1_hd U598 ( .A(n496), .B(n449), .Y(n453) );
  oa211d1_hd U599 ( .A(n454), .B(n457), .C(n451), .D(n450), .Y(n171) );
  ao21d1_hd U600 ( .A(n453), .B(n452), .C(n519), .Y(n458) );
  oa21d1_hd U601 ( .A(z_m[9]), .B(n496), .C(n454), .Y(n455) );
  ao22d1_hd U602 ( .A(n232), .B(value[18]), .C(z_m[10]), .D(n455), .Y(n456) );
  oa21d1_hd U603 ( .A(n458), .B(n457), .C(n456), .Y(n170) );
  ao22d1_hd U604 ( .A(n232), .B(value[19]), .C(n519), .D(z_m[10]), .Y(n461) );
  oa21d1_hd U605 ( .A(n459), .B(n564), .C(n501), .Y(n462) );
  oa211d1_hd U606 ( .A(z_m[11]), .B(n464), .C(n461), .D(n460), .Y(n169) );
  ao21d1_hd U607 ( .A(n507), .B(n463), .C(n462), .Y(n468) );
  oa21d1_hd U608 ( .A(z_m[12]), .B(n464), .C(n508), .Y(n465) );
  ao22d1_hd U609 ( .A(n232), .B(value[20]), .C(z_m[11]), .D(n465), .Y(n466) );
  oa21d1_hd U610 ( .A(n468), .B(n467), .C(n466), .Y(n168) );
  ao21d1_hd U611 ( .A(n570), .B(n469), .C(n489), .Y(n474) );
  ao22d1_hd U612 ( .A(n232), .B(value[21]), .C(n519), .D(z_m[12]), .Y(n471) );
  nr2d1_hd U613 ( .A(n496), .B(n469), .Y(n473) );
  oa211d1_hd U614 ( .A(n474), .B(n477), .C(n471), .D(n470), .Y(n167) );
  ivd1_hd U615 ( .A(z_m[14]), .Y(n472) );
  ao21d1_hd U616 ( .A(n473), .B(n472), .C(n519), .Y(n478) );
  oa21d1_hd U617 ( .A(z_m[13]), .B(n496), .C(n474), .Y(n475) );
  ao22d1_hd U618 ( .A(n232), .B(value[22]), .C(z_m[14]), .D(n475), .Y(n476) );
  oa21d1_hd U619 ( .A(n478), .B(n477), .C(n476), .Y(n166) );
  ao22d1_hd U620 ( .A(n232), .B(value[23]), .C(n519), .D(z_m[14]), .Y(n481) );
  oa21d1_hd U621 ( .A(n479), .B(n564), .C(n501), .Y(n482) );
  oa211d1_hd U622 ( .A(z_m[15]), .B(n484), .C(n481), .D(n480), .Y(n165) );
  ao21d1_hd U623 ( .A(n507), .B(n483), .C(n482), .Y(n488) );
  oa21d1_hd U624 ( .A(z_m[16]), .B(n484), .C(n508), .Y(n485) );
  ao22d1_hd U625 ( .A(n232), .B(value[24]), .C(z_m[15]), .D(n485), .Y(n486) );
  oa21d1_hd U626 ( .A(n488), .B(n487), .C(n486), .Y(n164) );
  ao21d1_hd U627 ( .A(n570), .B(n490), .C(n489), .Y(n495) );
  ao22d1_hd U628 ( .A(n232), .B(value[25]), .C(n519), .D(z_m[16]), .Y(n492) );
  nr2d1_hd U629 ( .A(n496), .B(n490), .Y(n494) );
  oa211d1_hd U630 ( .A(n495), .B(n499), .C(n492), .D(n491), .Y(n163) );
  ivd1_hd U631 ( .A(z_m[18]), .Y(n493) );
  ao21d1_hd U632 ( .A(n494), .B(n493), .C(n519), .Y(n500) );
  oa21d1_hd U633 ( .A(z_m[17]), .B(n496), .C(n495), .Y(n497) );
  ao22d1_hd U634 ( .A(n232), .B(value[26]), .C(z_m[18]), .D(n497), .Y(n498) );
  oa21d1_hd U635 ( .A(n500), .B(n499), .C(n498), .Y(n162) );
  ao22d1_hd U636 ( .A(n232), .B(value[27]), .C(n519), .D(z_m[18]), .Y(n504) );
  oa21d1_hd U637 ( .A(n502), .B(n564), .C(n501), .Y(n505) );
  oa211d1_hd U638 ( .A(z_m[19]), .B(n509), .C(n504), .D(n503), .Y(n161) );
  ao21d1_hd U639 ( .A(n507), .B(n506), .C(n505), .Y(n513) );
  oa21d1_hd U640 ( .A(z_m[20]), .B(n509), .C(n508), .Y(n510) );
  ao22d1_hd U641 ( .A(n232), .B(value[28]), .C(z_m[19]), .D(n510), .Y(n511) );
  oa21d1_hd U642 ( .A(n513), .B(n512), .C(n511), .Y(n160) );
  ao22d1_hd U643 ( .A(n232), .B(value[29]), .C(n519), .D(z_m[20]), .Y(n516) );
  oa211d1_hd U644 ( .A(n518), .B(n517), .C(n516), .D(n515), .Y(n159) );
  ao22d1_hd U645 ( .A(n232), .B(value[30]), .C(n519), .D(z_m[21]), .Y(n523) );
  oa211d1_hd U646 ( .A(z_m[22]), .B(n524), .C(n523), .D(n522), .Y(n158) );
  nr4d1_hd U647 ( .A(n534), .B(n533), .C(n532), .D(n531), .Y(n535) );
  nd4d1_hd U648 ( .A(z_m[22]), .B(z_m[21]), .C(n536), .D(n535), .Y(n537) );
  nr4d1_hd U649 ( .A(n540), .B(n539), .C(n538), .D(n537), .Y(n542) );
  ivd1_hd U650 ( .A(n579), .Y(n549) );
  ivd1_hd U651 ( .A(z_e[3]), .Y(n573) );
  nr2d1_hd U652 ( .A(n573), .B(n572), .Y(n576) );
  nr2d1_hd U653 ( .A(n583), .B(n545), .Y(n551) );
  nr2d1_hd U654 ( .A(z_e[7]), .B(n555), .Y(n547) );
  ivd1_hd U655 ( .A(n583), .Y(n571) );
  ivd1_hd U656 ( .A(z_e[5]), .Y(n550) );
  scg6d1_hd U657 ( .A(n545), .B(n570), .C(n569), .Y(n553) );
  ao21d1_hd U658 ( .A(n571), .B(n550), .C(n553), .Y(n556) );
  oa21d1_hd U659 ( .A(z_e[6]), .B(n583), .C(n556), .Y(n546) );
  ao22d1_hd U660 ( .A(z_e[6]), .B(n547), .C(z_e[7]), .D(n546), .Y(n548) );
  oa211d1_hd U661 ( .A(n549), .B(N172), .C(n548), .D(n557), .Y(n157) );
  ao22d1_hd U662 ( .A(n579), .B(N170), .C(n551), .D(n550), .Y(n552) );
  scg15d1_hd U663 ( .A(z_e[5]), .B(n553), .C(n552), .D(n557), .Y(n156) );
  ao22d1_hd U664 ( .A(z_e[6]), .B(n556), .C(n555), .D(n554), .Y(n558) );
  scg17d1_hd U665 ( .A(n579), .B(N171), .C(n558), .D(n557), .Y(n155) );
  oa21d1_hd U666 ( .A(n571), .B(n579), .C(N165), .Y(n560) );
  oa211d1_hd U667 ( .A(N165), .B(n563), .C(n581), .D(n560), .Y(n154) );
  ao22d1_hd U668 ( .A(n569), .B(z_e[1]), .C(n579), .D(N166), .Y(n561) );
  oa211d1_hd U669 ( .A(n583), .B(N166), .C(n561), .D(n581), .Y(n153) );
  oa21d1_hd U670 ( .A(n565), .B(n564), .C(n563), .Y(n566) );
  ao22d1_hd U671 ( .A(z_e[2]), .B(n566), .C(n579), .D(N167), .Y(n567) );
  oa211d1_hd U672 ( .A(n583), .B(n568), .C(n567), .D(n581), .Y(n152) );
  ao21d1_hd U673 ( .A(n570), .B(n572), .C(n569), .Y(n578) );
  oa22d1_hd U674 ( .A(n578), .B(n573), .C(n572), .D(n577), .Y(n574) );
  ao22d1_hd U675 ( .A(z_e[4]), .B(n580), .C(n579), .D(N169), .Y(n582) );
  oa211d1_hd U676 ( .A(n584), .B(n583), .C(n582), .D(n581), .Y(n150) );
endmodule

