
module float_adder ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N394, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3,
         C91_DATA2_4, C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8,
         C91_DATA2_9, RSOP_150_C1_CONTROL1, n1, n2, n18, n28, n29, n93, n103,
         n104, n105, n106, n107, n108, n110, n111, n112, n124, n125, n127,
         n128, n129, n130, n131, n132, n136, n265, n266, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n509, n511, C1_Z_0, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23, C2_Z_22,
         C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16, C2_Z_15,
         C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8, C2_Z_7,
         C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0, C3_Z_26,
         C3_Z_25, C3_Z_24, C3_Z_23, C3_Z_22, C3_Z_21, C3_Z_20, C3_Z_19,
         C3_Z_18, C3_Z_17, C3_Z_16, C3_Z_15, C3_Z_14, C3_Z_13, C3_Z_12,
         C3_Z_11, C3_Z_10, C3_Z_9, C3_Z_8, C3_Z_7, C3_Z_6, C3_Z_5, C3_Z_4,
         C3_Z_3, C3_Z_2, C3_Z_1, C3_Z_0, DP_OP_43J1_124_6938_n58,
         DP_OP_43J1_124_6938_n57, DP_OP_43J1_124_6938_n56,
         DP_OP_43J1_124_6938_n55, DP_OP_43J1_124_6938_n54,
         DP_OP_43J1_124_6938_n53, DP_OP_43J1_124_6938_n52,
         DP_OP_43J1_124_6938_n51, DP_OP_43J1_124_6938_n50,
         DP_OP_43J1_124_6938_n49, DP_OP_43J1_124_6938_n48,
         DP_OP_43J1_124_6938_n47, DP_OP_43J1_124_6938_n46,
         DP_OP_43J1_124_6938_n45, DP_OP_43J1_124_6938_n44,
         DP_OP_43J1_124_6938_n43, DP_OP_43J1_124_6938_n42,
         DP_OP_43J1_124_6938_n41, DP_OP_43J1_124_6938_n40,
         DP_OP_43J1_124_6938_n39, DP_OP_43J1_124_6938_n38,
         DP_OP_43J1_124_6938_n37, DP_OP_43J1_124_6938_n36,
         DP_OP_43J1_124_6938_n35, DP_OP_43J1_124_6938_n34,
         DP_OP_43J1_124_6938_n33, DP_OP_43J1_124_6938_n32,
         DP_OP_43J1_124_6938_n27, DP_OP_43J1_124_6938_n26,
         DP_OP_43J1_124_6938_n25, DP_OP_43J1_124_6938_n24,
         DP_OP_43J1_124_6938_n23, DP_OP_43J1_124_6938_n22,
         DP_OP_43J1_124_6938_n21, DP_OP_43J1_124_6938_n20,
         DP_OP_43J1_124_6938_n19, DP_OP_43J1_124_6938_n18,
         DP_OP_43J1_124_6938_n17, DP_OP_43J1_124_6938_n16,
         DP_OP_43J1_124_6938_n15, DP_OP_43J1_124_6938_n14,
         DP_OP_43J1_124_6938_n13, DP_OP_43J1_124_6938_n12,
         DP_OP_43J1_124_6938_n11, DP_OP_43J1_124_6938_n10,
         DP_OP_43J1_124_6938_n9, DP_OP_43J1_124_6938_n8,
         DP_OP_43J1_124_6938_n7, DP_OP_43J1_124_6938_n6,
         DP_OP_43J1_124_6938_n5, DP_OP_43J1_124_6938_n4,
         DP_OP_43J1_124_6938_n3, DP_OP_43J1_124_6938_n2,
         DP_OP_43J1_124_6938_n1, DP_OP_154J1_137_6175_n25,
         DP_OP_154J1_137_6175_n9, DP_OP_154J1_137_6175_n8,
         DP_OP_154J1_137_6175_n7, DP_OP_154J1_137_6175_n6,
         DP_OP_154J1_137_6175_n5, DP_OP_154J1_137_6175_n4,
         DP_OP_154J1_137_6175_n3, DP_OP_154J1_137_6175_n2,
         DP_OP_154J1_137_6175_n1, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  scg21d1_hd U117 ( .A(o_AB_ACK), .B(n104), .C(n730), .D(i_RST), .Y(n499) );
  oa22d1_hd U119 ( .A(n106), .B(n107), .C(n29), .D(n108), .Y(n500) );
  oa21d1_hd U121 ( .A(n573), .B(n108), .C(n110), .Y(n501) );
  scg6d1_hd U122 ( .A(n111), .B(DP_OP_154J1_137_6175_n25), .C(n107), .Y(n110)
         );
  oa22d1_hd U123 ( .A(n112), .B(n107), .C(n816), .D(n108), .Y(n502) );
  oa21d1_hd U134 ( .A(n28), .B(n108), .C(n124), .Y(n505) );
  scg6d1_hd U135 ( .A(n728), .B(n812), .C(n107), .Y(n124) );
  nd4d1_hd U137 ( .A(n111), .B(n127), .C(n103), .D(n18), .Y(n108) );
  nr4d1_hd U138 ( .A(n719), .B(n128), .C(n129), .D(n130), .Y(n127) );
  scg16d1_hd U139 ( .A(n636), .B(N394), .C(N41), .Y(n130) );
  ao211d1_hd U143 ( .A(n721), .B(n132), .C(i_RST), .D(n136), .Y(n506) );
  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J1_137_6175_U10 ( .A(n676), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J1_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J1_137_6175_U9 ( .A(n677), .B(z_e[2]), .CI(
        DP_OP_154J1_137_6175_n9), .CO(DP_OP_154J1_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J1_137_6175_U8 ( .A(n675), .B(z_e[3]), .CI(
        DP_OP_154J1_137_6175_n8), .CO(DP_OP_154J1_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J1_137_6175_U7 ( .A(n677), .B(z_e[4]), .CI(
        DP_OP_154J1_137_6175_n7), .CO(DP_OP_154J1_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J1_137_6175_U6 ( .A(n675), .B(z_e[5]), .CI(
        DP_OP_154J1_137_6175_n6), .CO(DP_OP_154J1_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J1_137_6175_U5 ( .A(n676), .B(z_e[6]), .CI(
        DP_OP_154J1_137_6175_n5), .CO(DP_OP_154J1_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J1_137_6175_U4 ( .A(n675), .B(z_e[7]), .CI(
        DP_OP_154J1_137_6175_n4), .CO(DP_OP_154J1_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J1_137_6175_U3 ( .A(n677), .B(z_e[8]), .CI(
        DP_OP_154J1_137_6175_n3), .CO(DP_OP_154J1_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n718), .CK(i_CLK), .Q(sum[26]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n718), .CK(i_CLK), .Q(sum[27]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J1_124_6938_U28 ( .A(C2_Z_0), .B(n680), .CI(
        DP_OP_43J1_124_6938_n58), .CO(DP_OP_43J1_124_6938_n27), .S(N310) );
  fad1_hd DP_OP_43J1_124_6938_U27 ( .A(DP_OP_43J1_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J1_124_6938_n27), .CO(DP_OP_43J1_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J1_124_6938_U26 ( .A(DP_OP_43J1_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J1_124_6938_n26), .CO(DP_OP_43J1_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J1_124_6938_U25 ( .A(DP_OP_43J1_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J1_124_6938_n25), .CO(DP_OP_43J1_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J1_124_6938_U24 ( .A(DP_OP_43J1_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J1_124_6938_n24), .CO(DP_OP_43J1_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J1_124_6938_U23 ( .A(DP_OP_43J1_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J1_124_6938_n23), .CO(DP_OP_43J1_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J1_124_6938_U22 ( .A(DP_OP_43J1_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J1_124_6938_n22), .CO(DP_OP_43J1_124_6938_n21), .S(N316)
         );
  fad1_hd DP_OP_43J1_124_6938_U2 ( .A(DP_OP_43J1_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J1_124_6938_n2), .CO(DP_OP_43J1_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J1_124_6938_U3 ( .A(DP_OP_43J1_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J1_124_6938_n3), .CO(DP_OP_43J1_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J1_124_6938_U21 ( .A(DP_OP_43J1_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J1_124_6938_n21), .CO(DP_OP_43J1_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J1_124_6938_U15 ( .A(DP_OP_43J1_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J1_124_6938_n15), .CO(DP_OP_43J1_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J1_124_6938_U16 ( .A(DP_OP_43J1_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J1_124_6938_n16), .CO(DP_OP_43J1_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J1_124_6938_U17 ( .A(DP_OP_43J1_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J1_124_6938_n17), .CO(DP_OP_43J1_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J1_124_6938_U18 ( .A(DP_OP_43J1_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J1_124_6938_n18), .CO(DP_OP_43J1_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J1_124_6938_U19 ( .A(DP_OP_43J1_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J1_124_6938_n19), .CO(DP_OP_43J1_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J1_124_6938_U20 ( .A(DP_OP_43J1_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J1_124_6938_n20), .CO(DP_OP_43J1_124_6938_n19), .S(N318)
         );
  xo2d1_hd DP_OP_154J1_137_6175_U2 ( .A(n675), .B(z_e[9]), .Y(
        DP_OP_154J1_137_6175_n1) );
  xo2d1_hd DP_OP_154J1_137_6175_U1 ( .A(DP_OP_154J1_137_6175_n2), .B(
        DP_OP_154J1_137_6175_n1), .Y(C91_DATA2_9) );
  xo2d1_hd DP_OP_43J1_124_6938_U40 ( .A(n684), .B(C3_Z_17), .Y(
        DP_OP_43J1_124_6938_n41) );
  xo2d1_hd DP_OP_43J1_124_6938_U41 ( .A(n684), .B(C3_Z_16), .Y(
        DP_OP_43J1_124_6938_n42) );
  xo2d1_hd DP_OP_43J1_124_6938_U38 ( .A(C1_Z_0), .B(C3_Z_19), .Y(
        DP_OP_43J1_124_6938_n39) );
  xo2d1_hd DP_OP_43J1_124_6938_U35 ( .A(n681), .B(C3_Z_22), .Y(
        DP_OP_43J1_124_6938_n36) );
  xo2d1_hd DP_OP_43J1_124_6938_U57 ( .A(n682), .B(C3_Z_0), .Y(
        DP_OP_43J1_124_6938_n58) );
  xo2d1_hd DP_OP_43J1_124_6938_U31 ( .A(n682), .B(C3_Z_26), .Y(
        DP_OP_43J1_124_6938_n32) );
  xo2d1_hd DP_OP_43J1_124_6938_U50 ( .A(n683), .B(C3_Z_7), .Y(
        DP_OP_43J1_124_6938_n51) );
  xo2d1_hd DP_OP_43J1_124_6938_U32 ( .A(n682), .B(C3_Z_25), .Y(
        DP_OP_43J1_124_6938_n33) );
  xo2d1_hd DP_OP_43J1_124_6938_U55 ( .A(n680), .B(C3_Z_2), .Y(
        DP_OP_43J1_124_6938_n56) );
  xo2d1_hd DP_OP_43J1_124_6938_U33 ( .A(n682), .B(C3_Z_24), .Y(
        DP_OP_43J1_124_6938_n34) );
  xo2d1_hd DP_OP_43J1_124_6938_U56 ( .A(n680), .B(C3_Z_1), .Y(
        DP_OP_43J1_124_6938_n57) );
  xo2d1_hd DP_OP_43J1_124_6938_U51 ( .A(n683), .B(C3_Z_6), .Y(
        DP_OP_43J1_124_6938_n52) );
  xo2d1_hd DP_OP_43J1_124_6938_U54 ( .A(n680), .B(C3_Z_3), .Y(
        DP_OP_43J1_124_6938_n55) );
  xo2d1_hd DP_OP_43J1_124_6938_U36 ( .A(C1_Z_0), .B(C3_Z_21), .Y(
        DP_OP_43J1_124_6938_n37) );
  xo2d1_hd DP_OP_43J1_124_6938_U39 ( .A(C1_Z_0), .B(C3_Z_18), .Y(
        DP_OP_43J1_124_6938_n40) );
  xo2d1_hd DP_OP_43J1_124_6938_U37 ( .A(C1_Z_0), .B(C3_Z_20), .Y(
        DP_OP_43J1_124_6938_n38) );
  fad1_hd DP_OP_43J1_124_6938_U4 ( .A(DP_OP_43J1_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J1_124_6938_n4), .CO(DP_OP_43J1_124_6938_n3), .S(N334) );
  xo2d1_hd DP_OP_43J1_124_6938_U1 ( .A(DP_OP_43J1_124_6938_n1), .B(n682), .Y(
        N337) );
  xo2d1_hd DP_OP_43J1_124_6938_U34 ( .A(n682), .B(C3_Z_23), .Y(
        DP_OP_43J1_124_6938_n35) );
  xo2d1_hd DP_OP_43J1_124_6938_U52 ( .A(n680), .B(C3_Z_5), .Y(
        DP_OP_43J1_124_6938_n53) );
  xo2d1_hd DP_OP_43J1_124_6938_U49 ( .A(n683), .B(C3_Z_8), .Y(
        DP_OP_43J1_124_6938_n50) );
  xo2d1_hd DP_OP_43J1_124_6938_U44 ( .A(n681), .B(C3_Z_13), .Y(
        DP_OP_43J1_124_6938_n45) );
  xo2d1_hd DP_OP_43J1_124_6938_U42 ( .A(n681), .B(C3_Z_15), .Y(
        DP_OP_43J1_124_6938_n43) );
  xo2d1_hd DP_OP_43J1_124_6938_U43 ( .A(n681), .B(C3_Z_14), .Y(
        DP_OP_43J1_124_6938_n44) );
  xo2d1_hd DP_OP_43J1_124_6938_U53 ( .A(n680), .B(C3_Z_4), .Y(
        DP_OP_43J1_124_6938_n54) );
  xo2d1_hd DP_OP_43J1_124_6938_U48 ( .A(n683), .B(C3_Z_9), .Y(
        DP_OP_43J1_124_6938_n49) );
  xo2d1_hd DP_OP_43J1_124_6938_U45 ( .A(n681), .B(C3_Z_12), .Y(
        DP_OP_43J1_124_6938_n46) );
  xo2d1_hd DP_OP_43J1_124_6938_U47 ( .A(n683), .B(C3_Z_10), .Y(
        DP_OP_43J1_124_6938_n48) );
  xo2d1_hd DP_OP_43J1_124_6938_U46 ( .A(n681), .B(C3_Z_11), .Y(
        DP_OP_43J1_124_6938_n47) );
  fad1_hd DP_OP_43J1_124_6938_U5 ( .A(DP_OP_43J1_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J1_124_6938_n5), .CO(DP_OP_43J1_124_6938_n4), .S(N333) );
  fad1_hd DP_OP_43J1_124_6938_U14 ( .A(DP_OP_43J1_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J1_124_6938_n14), .CO(DP_OP_43J1_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J1_124_6938_U6 ( .A(DP_OP_43J1_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J1_124_6938_n6), .CO(DP_OP_43J1_124_6938_n5), .S(N332) );
  fad1_hd DP_OP_43J1_124_6938_U13 ( .A(DP_OP_43J1_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J1_124_6938_n13), .CO(DP_OP_43J1_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J1_124_6938_U12 ( .A(DP_OP_43J1_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J1_124_6938_n12), .CO(DP_OP_43J1_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J1_124_6938_U11 ( .A(DP_OP_43J1_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J1_124_6938_n11), .CO(DP_OP_43J1_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J1_124_6938_U10 ( .A(DP_OP_43J1_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J1_124_6938_n10), .CO(DP_OP_43J1_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J1_124_6938_U9 ( .A(DP_OP_43J1_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J1_124_6938_n9), .CO(DP_OP_43J1_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J1_124_6938_U8 ( .A(DP_OP_43J1_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J1_124_6938_n8), .CO(DP_OP_43J1_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J1_124_6938_U7 ( .A(DP_OP_43J1_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J1_124_6938_n7), .CO(DP_OP_43J1_124_6938_n6), .S(N331) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n527), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n527), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n526), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n721), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n528), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n528), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n509), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n527), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n522), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n531), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n530), .CK(i_CLK), .Q(b[23]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n517), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n518), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n526), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n526), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n722), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n528), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n517), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n730), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n730), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n720), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n720), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n526), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n509), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n721), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n522), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n518), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n730), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n529), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n516), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n517), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n527), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n720), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n530), .CK(i_CLK), .Q(b[26]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n520), .CK(i_CLK), .Q(b[22]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n531), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n529), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n517), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n516), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n531), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n521), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n516), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n531), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n530), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n516), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n519), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n520), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n519), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n529), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n522), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n518), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n516), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n530), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n520), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n521), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n722), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n722), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n528), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n720), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n527), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n527), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n519), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n520), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n520), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n518), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n521), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n521), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n522), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n520), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n522), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n517), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n519), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n730), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n518), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n529), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n529), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n530), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n516), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n730), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n265), .CK(i_CLK), .Q(guard) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1376), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1376), .CK(i_CLK), .Q(a_s) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n531), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n522), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n521), .CK(i_CLK), .Q(b[28]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n519), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n526), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n722), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n528), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n528), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n720), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n722), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n529), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n518), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n519), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n531), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n530), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n521), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n93), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n525), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n93), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n523), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n715), .CK(i_CLK), .Q(sum[1]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n524), .CK(i_CLK), .Q(sum[2]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n524), .CK(i_CLK), .Q(sum[3]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n525), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n719), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n715), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n715), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n524), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n523), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n719), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n718), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n715), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n525), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n523), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n523), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n719), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n524), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n525), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n525), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n523), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n715), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n524), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n524), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n525), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n719), .CK(i_CLK), .Q(sum[25]) );
  clknd2d1_hd U523 ( .A(n557), .B(n946), .Y(n837) );
  clknd2d1_hd U524 ( .A(n559), .B(n548), .Y(n838) );
  clknd2d1_hd U525 ( .A(n549), .B(n558), .Y(n868) );
  clknd2d1_hd U526 ( .A(n1335), .B(b_e[2]), .Y(n905) );
  clknd2d1_hd U527 ( .A(n1251), .B(a_e[9]), .Y(n922) );
  clknd2d1_hd U528 ( .A(b_e[3]), .B(n1343), .Y(n906) );
  clknd2d1_hd U529 ( .A(b_e[7]), .B(n1385), .Y(n917) );
  clknd2d1_hd U530 ( .A(b_e[0]), .B(n1328), .Y(n901) );
  clknd2d1_hd U531 ( .A(z_e[7]), .B(z_e[8]), .Y(n1001) );
  clknd2d1_hd U532 ( .A(n822), .B(n821), .Y(n896) );
  clknd2d1_hd U533 ( .A(n884), .B(n885), .Y(n808) );
  clknd2d1_hd U534 ( .A(n883), .B(n882), .Y(n884) );
  clknd2d1_hd U535 ( .A(n922), .B(n921), .Y(n957) );
  clknd2d1_hd U536 ( .A(n1358), .B(n957), .Y(n1247) );
  clknd2d1_hd U537 ( .A(n1012), .B(n1040), .Y(n1050) );
  clknd2d1_hd U538 ( .A(z_m[0]), .B(n563), .Y(n1011) );
  clknd2d1_hd U539 ( .A(n28), .B(state[2]), .Y(n995) );
  clknd2d1_hd U540 ( .A(n1020), .B(n1123), .Y(n1021) );
  clknd2d1_hd U541 ( .A(n1014), .B(n1060), .Y(n1070) );
  clknd2d1_hd U542 ( .A(n1016), .B(n1080), .Y(n1090) );
  clknd2d1_hd U543 ( .A(n1018), .B(n1100), .Y(n1111) );
  clknd2d1_hd U544 ( .A(n1184), .B(n1183), .Y(n1185) );
  clknd2d1_hd U545 ( .A(n1190), .B(n1189), .Y(n1191) );
  clknd2d1_hd U546 ( .A(n814), .B(n1210), .Y(n1158) );
  clknd2d1_hd U547 ( .A(n1205), .B(n1210), .Y(n1176) );
  clknd2d1_hd U548 ( .A(n813), .B(n1207), .Y(n1157) );
  clknd2d1_hd U549 ( .A(n808), .B(n809), .Y(n811) );
  clknd2d1_hd U550 ( .A(n813), .B(n741), .Y(n1204) );
  clknd2d1_hd U551 ( .A(n1388), .B(n1160), .Y(n1207) );
  clknd2d1_hd U552 ( .A(n573), .B(state[0]), .Y(n1156) );
  clknd2d1_hd U553 ( .A(n818), .B(n1189), .Y(n1173) );
  clknd2d1_hd U554 ( .A(n567), .B(z_m[10]), .Y(n1015) );
  clknd2d1_hd U555 ( .A(n571), .B(z_m[18]), .Y(n1019) );
  clknd2d1_hd U556 ( .A(n614), .B(z_m[6]), .Y(n1013) );
  clknd2d1_hd U557 ( .A(n569), .B(z_m[14]), .Y(n1017) );
  nid1_hd U558 ( .A(n810), .Y(n693) );
  nid1_hd U559 ( .A(n810), .Y(n694) );
  clknd2d1_hd U560 ( .A(n678), .B(n811), .Y(C1_Z_0) );
  nid1_hd U561 ( .A(n694), .Y(n685) );
  nid1_hd U562 ( .A(n693), .Y(n690) );
  nid1_hd U563 ( .A(n684), .Y(n681) );
  ivd1_hd U564 ( .A(n705), .Y(n701) );
  nid1_hd U565 ( .A(n694), .Y(n686) );
  nid1_hd U566 ( .A(n693), .Y(n691) );
  nid1_hd U567 ( .A(C1_Z_0), .Y(n683) );
  nid1_hd U568 ( .A(n694), .Y(n687) );
  nid1_hd U569 ( .A(n683), .Y(n680) );
  or2d2_hd U570 ( .A(n808), .B(n815), .Y(n678) );
  nid1_hd U571 ( .A(n678), .Y(n705) );
  nid1_hd U572 ( .A(n103), .Y(n105) );
  clknd2d1_hd U573 ( .A(n1369), .B(n1368), .Y(n1370) );
  clknd2d1_hd U574 ( .A(n93), .B(n1323), .Y(n1373) );
  clknd2d1_hd U575 ( .A(n573), .B(n1243), .Y(n1258) );
  clknd2d1_hd U576 ( .A(n817), .B(n816), .Y(n1257) );
  clknd2d1_hd U577 ( .A(n577), .B(n1264), .Y(n1271) );
  clknd2d1_hd U578 ( .A(b[24]), .B(b[23]), .Y(n1269) );
  clknd2d1_hd U579 ( .A(n1365), .B(n1329), .Y(n1336) );
  clknd2d1_hd U580 ( .A(a[24]), .B(a[23]), .Y(n1334) );
  clknd2d1_hd U581 ( .A(b_e[4]), .B(n1282), .Y(n1293) );
  clknd2d1_hd U582 ( .A(n578), .B(n1294), .Y(n1300) );
  clknd2d1_hd U583 ( .A(n817), .B(n573), .Y(n1259) );
  clknd2d1_hd U584 ( .A(N41), .B(n108), .Y(n107) );
  clknd2d1_hd U585 ( .A(a_e[4]), .B(n1347), .Y(n1359) );
  clknd2d1_hd U586 ( .A(n1365), .B(n1360), .Y(n1368) );
  clknd2d1_hd U587 ( .A(n1361), .B(a[28]), .Y(n1367) );
  clknd2d1_hd U588 ( .A(n1295), .B(b[28]), .Y(n1303) );
  clknd2d1_hd U589 ( .A(n1301), .B(n1300), .Y(n1306) );
  clknd2d1_hd U590 ( .A(n1323), .B(n1358), .Y(n1379) );
  clknd2d1_hd U591 ( .A(a_e[6]), .B(n1364), .Y(n1378) );
  clknd2d1_hd U592 ( .A(n1372), .B(n1377), .Y(n1383) );
  clknd2d1_hd U593 ( .A(n648), .B(n1298), .Y(n1316) );
  clknd2d1_hd U594 ( .A(n1305), .B(n1310), .Y(n1318) );
  clknd2d1_hd U595 ( .A(n615), .B(n1029), .Y(n1033) );
  clknd2d1_hd U596 ( .A(n659), .B(n1040), .Y(n1045) );
  clknd2d1_hd U597 ( .A(n1152), .B(sum[27]), .Y(n1025) );
  clknd2d1_hd U598 ( .A(n657), .B(n1060), .Y(n1065) );
  clknd2d1_hd U599 ( .A(n658), .B(n1217), .Y(n1029) );
  clknd2d1_hd U600 ( .A(z_m[21]), .B(n1136), .Y(n1139) );
  clknd2d1_hd U601 ( .A(n658), .B(n1080), .Y(n1085) );
  clknd2d1_hd U602 ( .A(n659), .B(n1100), .Y(n1105) );
  clknd2d1_hd U603 ( .A(n657), .B(n1123), .Y(n1129) );
  clknd2d1_hd U604 ( .A(n753), .B(n752), .Y(n758) );
  clknd2d1_hd U605 ( .A(n763), .B(n762), .Y(n768) );
  clknd2d1_hd U606 ( .A(n773), .B(n772), .Y(n779) );
  clknd2d1_hd U607 ( .A(n1244), .B(n1238), .Y(n1201) );
  clknd2d1_hd U608 ( .A(n811), .B(n809), .Y(n810) );
  nid1_hd U609 ( .A(n684), .Y(n682) );
  clknd2d1_hd U610 ( .A(n814), .B(b_s), .Y(n1203) );
  clknd2d1_hd U611 ( .A(n814), .B(n1207), .Y(n1209) );
  nr3d1_hd U612 ( .A(state[2]), .B(n28), .C(n1156), .Y(n1244) );
  clknd2d1_hd U613 ( .A(n1175), .B(n1174), .Y(n1238) );
  clknd2d1_hd U614 ( .A(n1237), .B(n1236), .Y(n1239) );
  clknd2d1_hd U615 ( .A(n649), .B(n1267), .Y(n1277) );
  clknd2d1_hd U616 ( .A(n578), .B(n1278), .Y(n1286) );
  clknd2d1_hd U617 ( .A(n1279), .B(b[26]), .Y(n1284) );
  clknd2d1_hd U618 ( .A(a_e[2]), .B(n1332), .Y(n1342) );
  clknd2d1_hd U619 ( .A(n1365), .B(n1343), .Y(n1351) );
  clknd2d1_hd U620 ( .A(n1344), .B(a[26]), .Y(n1349) );
  nid1_hd U621 ( .A(n523), .Y(n715) );
  clknd2d1_hd U622 ( .A(n1150), .B(n1006), .Y(n265) );
  ivd1_hd U623 ( .A(n103), .Y(n530) );
  clknd2d1_hd U624 ( .A(n577), .B(n1267), .Y(n1276) );
  clknd2d1_hd U625 ( .A(n647), .B(n1364), .Y(n1375) );
  clknd2d1_hd U626 ( .A(n1367), .B(n1366), .Y(n1371) );
  clknd2d1_hd U627 ( .A(n647), .B(n1347), .Y(n1356) );
  clknd2d1_hd U628 ( .A(n578), .B(n1282), .Y(n1291) );
  clknd2d1_hd U629 ( .A(n647), .B(n1332), .Y(n1341) );
  clknd2d1_hd U630 ( .A(n578), .B(n1298), .Y(n1309) );
  clknd2d1_hd U631 ( .A(n1303), .B(n1302), .Y(n1304) );
  clknd2d1_hd U632 ( .A(n653), .B(z_e[5]), .Y(n790) );
  clknd2d1_hd U633 ( .A(C91_DATA2_5), .B(n618), .Y(n791) );
  clknd2d1_hd U634 ( .A(n805), .B(z_e[1]), .Y(n798) );
  clknd2d1_hd U635 ( .A(n617), .B(C91_DATA2_1), .Y(n799) );
  clknd2d1_hd U636 ( .A(n653), .B(z_e[6]), .Y(n788) );
  clknd2d1_hd U637 ( .A(C91_DATA2_6), .B(n617), .Y(n789) );
  clknd2d1_hd U638 ( .A(n653), .B(z_e[7]), .Y(n786) );
  clknd2d1_hd U639 ( .A(C91_DATA2_7), .B(n617), .Y(n787) );
  clknd2d1_hd U640 ( .A(n805), .B(z_e[3]), .Y(n794) );
  clknd2d1_hd U641 ( .A(C91_DATA2_3), .B(n618), .Y(n795) );
  clknd2d1_hd U642 ( .A(n805), .B(z_e[2]), .Y(n796) );
  clknd2d1_hd U643 ( .A(C91_DATA2_2), .B(n617), .Y(n797) );
  clknd2d1_hd U644 ( .A(n805), .B(z_e[4]), .Y(n792) );
  clknd2d1_hd U645 ( .A(C91_DATA2_4), .B(n618), .Y(n793) );
  clknd2d1_hd U646 ( .A(n653), .B(z_e[8]), .Y(n806) );
  clknd2d1_hd U647 ( .A(C91_DATA2_8), .B(n618), .Y(n807) );
  clknd2d1_hd U648 ( .A(n718), .B(a_e[9]), .Y(n802) );
  clknd2d1_hd U649 ( .A(C91_DATA2_9), .B(n617), .Y(n803) );
  clknd2d1_hd U650 ( .A(n1146), .B(sum[3]), .Y(n1026) );
  clknd2d1_hd U651 ( .A(n724), .B(z[31]), .Y(n1241) );
  ivd1_hd U652 ( .A(n105), .Y(n531) );
  ivd1_hd U653 ( .A(n105), .Y(n516) );
  ivd1_hd U654 ( .A(n105), .Y(n517) );
  ivd1_hd U655 ( .A(n103), .Y(n518) );
  ivd1_hd U656 ( .A(n103), .Y(n519) );
  ivd1_hd U657 ( .A(n105), .Y(n520) );
  ivd1_hd U658 ( .A(n103), .Y(n521) );
  ivd1_hd U659 ( .A(n105), .Y(n522) );
  or2d1_hd U660 ( .A(state[0]), .B(n1259), .Y(n511) );
  ivd1_hd U661 ( .A(n511), .Y(n523) );
  ivd1_hd U662 ( .A(n511), .Y(n524) );
  ivd1_hd U663 ( .A(n511), .Y(n525) );
  nid1_hd U664 ( .A(n509), .Y(n526) );
  nid1_hd U665 ( .A(n509), .Y(n527) );
  nid1_hd U666 ( .A(n509), .Y(n528) );
  ivd1_hd U667 ( .A(n105), .Y(n529) );
  nid1_hd U668 ( .A(n678), .Y(n706) );
  nid1_hd U669 ( .A(C1_Z_0), .Y(n684) );
  xn2d1_hd U670 ( .A(a_s), .B(b_s), .Y(n815) );
  ivd1_hd U671 ( .A(n815), .Y(n809) );
  nid1_hd U672 ( .A(n694), .Y(n689) );
  ivd1_hd U673 ( .A(n705), .Y(n702) );
  xo2d1_hd U674 ( .A(n780), .B(n779), .Y(n784) );
  scg6d1_hd U675 ( .A(n812), .B(n785), .C(n805), .Y(n804) );
  scg2d1_hd U676 ( .A(n686), .B(a_m[12]), .C(b_m[12]), .D(n701), .Y(C2_Z_12)
         );
  scg2d1_hd U677 ( .A(n689), .B(b_m[20]), .C(n604), .D(n698), .Y(C3_Z_20) );
  scg2d1_hd U678 ( .A(n691), .B(b_m[9]), .C(n553), .D(n696), .Y(C3_Z_9) );
  scg2d1_hd U679 ( .A(n686), .B(a_m[9]), .C(b_m[9]), .D(n701), .Y(C2_Z_9) );
  scg2d1_hd U680 ( .A(n686), .B(a_m[13]), .C(b_m[13]), .D(n701), .Y(C2_Z_13)
         );
  scg2d1_hd U681 ( .A(n688), .B(b_m[26]), .C(a_m[26]), .D(n699), .Y(C3_Z_26)
         );
  scg2d1_hd U682 ( .A(n692), .B(b_m[0]), .C(a_m[0]), .D(n695), .Y(C3_Z_0) );
  scg2d1_hd U683 ( .A(n689), .B(b_m[18]), .C(n594), .D(n697), .Y(C3_Z_18) );
  scg2d1_hd U684 ( .A(n691), .B(b_m[10]), .C(n596), .D(n696), .Y(C3_Z_10) );
  scg2d1_hd U685 ( .A(n690), .B(n608), .C(n600), .D(n696), .Y(C3_Z_12) );
  scg2d1_hd U686 ( .A(n689), .B(b_m[22]), .C(n541), .D(n698), .Y(C3_Z_22) );
  scg2d1_hd U687 ( .A(n690), .B(b_m[15]), .C(a_m[15]), .D(n697), .Y(C3_Z_15)
         );
  scg2d1_hd U688 ( .A(n690), .B(n557), .C(a_m[17]), .D(n697), .Y(C3_Z_17) );
  scg2d1_hd U689 ( .A(n686), .B(a_m[10]), .C(b_m[10]), .D(n701), .Y(C2_Z_10)
         );
  scg2d1_hd U690 ( .A(n690), .B(b_m[16]), .C(n590), .D(n697), .Y(C3_Z_16) );
  scg2d1_hd U691 ( .A(n690), .B(b_m[13]), .C(n547), .D(n697), .Y(C3_Z_13) );
  scg2d1_hd U692 ( .A(n691), .B(n543), .C(n539), .D(n699), .Y(C3_Z_11) );
  scg2d1_hd U693 ( .A(n686), .B(a_m[14]), .C(n551), .D(n701), .Y(C2_Z_14) );
  scg2d1_hd U694 ( .A(n685), .B(n606), .C(b_m[15]), .D(n702), .Y(C2_Z_15) );
  scg2d1_hd U695 ( .A(n690), .B(n551), .C(n592), .D(n697), .Y(C3_Z_14) );
  scg2d1_hd U696 ( .A(n685), .B(n549), .C(b_m[19]), .D(n702), .Y(C2_Z_19) );
  scg2d1_hd U697 ( .A(n688), .B(b_m[24]), .C(n561), .D(n698), .Y(C3_Z_24) );
  scg2d1_hd U698 ( .A(n686), .B(n539), .C(b_m[11]), .D(n701), .Y(C2_Z_11) );
  scg2d1_hd U699 ( .A(n685), .B(n594), .C(b_m[18]), .D(n702), .Y(C2_Z_18) );
  scg2d1_hd U700 ( .A(n689), .B(n610), .C(a_m[23]), .D(n698), .Y(C3_Z_23) );
  scg2d1_hd U701 ( .A(n685), .B(a_m[20]), .C(n586), .D(n702), .Y(C2_Z_20) );
  scg2d1_hd U702 ( .A(n689), .B(b_m[21]), .C(a_m[21]), .D(n698), .Y(C3_Z_21)
         );
  scg2d1_hd U703 ( .A(n685), .B(a_m[16]), .C(b_m[16]), .D(n702), .Y(C2_Z_16)
         );
  scg2d1_hd U704 ( .A(n685), .B(a_m[17]), .C(b_m[17]), .D(n702), .Y(C2_Z_17)
         );
  scg2d1_hd U705 ( .A(n689), .B(b_m[19]), .C(a_m[19]), .D(n698), .Y(C3_Z_19)
         );
  scg2d1_hd U706 ( .A(n692), .B(b_m[1]), .C(a_m[1]), .D(n695), .Y(C3_Z_1) );
  scg2d1_hd U707 ( .A(n688), .B(a_m[2]), .C(b_m[2]), .D(n699), .Y(C2_Z_2) );
  scg2d1_hd U708 ( .A(n688), .B(a_m[1]), .C(b_m[1]), .D(n699), .Y(C2_Z_1) );
  scg2d1_hd U709 ( .A(n692), .B(b_m[2]), .C(a_m[2]), .D(n695), .Y(C3_Z_2) );
  scg2d1_hd U710 ( .A(n687), .B(a_m[3]), .C(b_m[3]), .D(n700), .Y(C2_Z_3) );
  scg2d1_hd U711 ( .A(n692), .B(b_m[3]), .C(a_m[3]), .D(n695), .Y(C3_Z_3) );
  scg2d1_hd U712 ( .A(n687), .B(a_m[4]), .C(b_m[4]), .D(n700), .Y(C2_Z_4) );
  scg2d1_hd U713 ( .A(n692), .B(b_m[4]), .C(n584), .D(n695), .Y(C3_Z_4) );
  scg2d1_hd U714 ( .A(n687), .B(a_m[5]), .C(b_m[5]), .D(n700), .Y(C2_Z_5) );
  scg2d1_hd U715 ( .A(n692), .B(n537), .C(a_m[5]), .D(n695), .Y(C3_Z_5) );
  scg2d1_hd U716 ( .A(n687), .B(a_m[6]), .C(b_m[6]), .D(n700), .Y(C2_Z_6) );
  scg2d1_hd U717 ( .A(n691), .B(b_m[6]), .C(n582), .D(n696), .Y(C3_Z_6) );
  scg2d1_hd U718 ( .A(n688), .B(a_m[0]), .C(b_m[0]), .D(n699), .Y(C2_Z_0) );
  scg2d1_hd U719 ( .A(n691), .B(n545), .C(n588), .D(n696), .Y(C3_Z_8) );
  scg2d1_hd U720 ( .A(n687), .B(a_m[8]), .C(b_m[8]), .D(n700), .Y(C2_Z_8) );
  scg2d1_hd U721 ( .A(n688), .B(b_m[25]), .C(a_m[25]), .D(n699), .Y(C3_Z_25)
         );
  scg2d1_hd U722 ( .A(n687), .B(a_m[7]), .C(b_m[7]), .D(n700), .Y(C2_Z_7) );
  scg2d1_hd U723 ( .A(n691), .B(n602), .C(a_m[7]), .D(n696), .Y(C3_Z_7) );
  nid1_hd U724 ( .A(n694), .Y(n688) );
  nid1_hd U725 ( .A(n693), .Y(n692) );
  or2d1_hd U726 ( .A(n1050), .B(n619), .Y(n1054) );
  or2d1_hd U727 ( .A(n1090), .B(n619), .Y(n1094) );
  or2d1_hd U728 ( .A(n1070), .B(n620), .Y(n1074) );
  or2d1_hd U729 ( .A(n1111), .B(n620), .Y(n1116) );
  scg2d1_hd U730 ( .A(n693), .B(a_m[23]), .C(b_m[23]), .D(n703), .Y(C2_Z_23)
         );
  scg2d1_hd U731 ( .A(n693), .B(a_m[22]), .C(n598), .D(n703), .Y(C2_Z_22) );
  scg2d1_hd U732 ( .A(n694), .B(n555), .C(b_m[21]), .D(n703), .Y(C2_Z_21) );
  scg2d1_hd U733 ( .A(n693), .B(a_m[24]), .C(n612), .D(n703), .Y(C2_Z_24) );
  scg2d1_hd U734 ( .A(n810), .B(a_m[25]), .C(b_m[25]), .D(n703), .Y(C2_Z_25)
         );
  scg2d1_hd U735 ( .A(n810), .B(a_m[26]), .C(n703), .D(b_m[26]), .Y(C2_Z_26)
         );
  nr2d1_hd U736 ( .A(n532), .B(n1250), .Y(n1307) );
  ad2d1_hd U737 ( .A(n615), .B(n1010), .Y(n1118) );
  or2d1_hd U738 ( .A(n532), .B(n1260), .Y(n1299) );
  or2d1_hd U739 ( .A(n1260), .B(n572), .Y(n1253) );
  scg6d1_hd U740 ( .A(n1388), .B(n1390), .C(n660), .Y(n1292) );
  or2d1_hd U741 ( .A(DP_OP_154J1_137_6175_n25), .B(n576), .Y(n1113) );
  ad2d1_hd U742 ( .A(n654), .B(n1358), .Y(n955) );
  nid1_hd U743 ( .A(n739), .Y(n738) );
  nid1_hd U744 ( .A(n125), .Y(n729) );
  nid1_hd U745 ( .A(n739), .Y(n737) );
  nid1_hd U746 ( .A(n731), .Y(n732) );
  nid1_hd U747 ( .A(n731), .Y(n739) );
  nid1_hd U748 ( .A(n1151), .Y(n714) );
  nid1_hd U749 ( .A(RSOP_150_C1_CONTROL1), .Y(n734) );
  nid1_hd U750 ( .A(RSOP_150_C1_CONTROL1), .Y(n735) );
  nid1_hd U751 ( .A(n1151), .Y(n713) );
  scg2d1_hd U752 ( .A(n778), .B(a_e[5]), .C(n777), .D(b_e[5]), .Y(n767) );
  or2d1_hd U753 ( .A(n1009), .B(n265), .Y(n1110) );
  scg9d1_hd U754 ( .A(n957), .B(n1260), .C(n625), .Y(n1255) );
  nid1_hd U755 ( .A(RSOP_150_C1_CONTROL1), .Y(n733) );
  nid1_hd U756 ( .A(n1151), .Y(n712) );
  nid1_hd U757 ( .A(RSOP_150_C1_CONTROL1), .Y(n736) );
  nid1_hd U758 ( .A(n1151), .Y(n711) );
  nid1_hd U759 ( .A(RSOP_150_C1_CONTROL1), .Y(n731) );
  scg6d1_hd U760 ( .A(n93), .B(n1157), .C(n1244), .Y(n125) );
  nid1_hd U761 ( .A(n707), .Y(n709) );
  nid1_hd U762 ( .A(n707), .Y(n708) );
  or2d1_hd U763 ( .A(n1250), .B(n1204), .Y(n1164) );
  nid1_hd U764 ( .A(n1146), .Y(n707) );
  nid1_hd U765 ( .A(n517), .Y(n730) );
  nid1_hd U766 ( .A(n1146), .Y(n710) );
  nid1_hd U767 ( .A(n719), .Y(n718) );
  scg2d1_hd U768 ( .A(n677), .B(z_m[23]), .C(n721), .D(n132), .Y(n129) );
  nid1_hd U769 ( .A(n722), .Y(n721) );
  nid1_hd U770 ( .A(n715), .Y(n719) );
  nid1_hd U771 ( .A(n720), .Y(n722) );
  ad2d1_hd U772 ( .A(n29), .B(n1245), .Y(n1376) );
  nr2bd1_hd U773 ( .AN(n1244), .B(n1177), .Y(n1163) );
  nid1_hd U774 ( .A(n526), .Y(n720) );
  ad4d1_hd U775 ( .A(n906), .B(n901), .C(n900), .D(n917), .Y(n902) );
  scg2d1_hd U776 ( .A(n540), .B(n598), .C(n953), .D(n610), .Y(n873) );
  or3d1_hd U777 ( .A(n816), .B(n574), .C(n995), .Y(n131) );
  ad4d1_hd U778 ( .A(n828), .B(n827), .C(n826), .D(n825), .Y(n829) );
  or4d1_hd U779 ( .A(a_e[3]), .B(a_e[2]), .C(a_e[1]), .D(n823), .Y(n824) );
  ad4d1_hd U780 ( .A(n1263), .B(n1251), .C(n1264), .D(n1249), .Y(n679) );
  ad2d1_hd U781 ( .A(i_Z_ACK), .B(o_Z_STB), .Y(n132) );
  or2d1_hd U782 ( .A(z_e[3]), .B(z_e[2]), .Y(n1172) );
  ivd1_hd U783 ( .A(n1292), .Y(n532) );
  ivd1_hd U784 ( .A(n1292), .Y(n533) );
  ivd1_hd U785 ( .A(n1307), .Y(n534) );
  ivd1_hd U786 ( .A(n1307), .Y(n535) );
  ivd1_hd U787 ( .A(b_m[5]), .Y(n536) );
  ivd1_hd U788 ( .A(n536), .Y(n537) );
  ivd1_hd U789 ( .A(a_m[11]), .Y(n538) );
  ivd1_hd U790 ( .A(n538), .Y(n539) );
  ivd1_hd U791 ( .A(a_m[22]), .Y(n540) );
  ivd1_hd U792 ( .A(n540), .Y(n541) );
  ivd1_hd U793 ( .A(b_m[11]), .Y(n542) );
  ivd1_hd U794 ( .A(n542), .Y(n543) );
  ivd1_hd U795 ( .A(b_m[8]), .Y(n544) );
  ivd1_hd U796 ( .A(n544), .Y(n545) );
  ivd1_hd U797 ( .A(a_m[13]), .Y(n546) );
  ivd1_hd U798 ( .A(n546), .Y(n547) );
  ivd1_hd U799 ( .A(a_m[19]), .Y(n548) );
  ivd1_hd U800 ( .A(n548), .Y(n549) );
  ivd1_hd U801 ( .A(b_m[14]), .Y(n550) );
  ivd1_hd U802 ( .A(n550), .Y(n551) );
  ivd1_hd U803 ( .A(a_m[9]), .Y(n552) );
  ivd1_hd U804 ( .A(n552), .Y(n553) );
  ivd1_hd U805 ( .A(a_m[21]), .Y(n554) );
  ivd1_hd U806 ( .A(n554), .Y(n555) );
  ivd1_hd U807 ( .A(b_m[17]), .Y(n556) );
  ivd1_hd U808 ( .A(n556), .Y(n557) );
  ivd1_hd U809 ( .A(b_m[19]), .Y(n558) );
  ivd1_hd U810 ( .A(n558), .Y(n559) );
  ivd1_hd U811 ( .A(a_m[24]), .Y(n560) );
  ivd1_hd U812 ( .A(n560), .Y(n561) );
  ivd1_hd U813 ( .A(z_m[1]), .Y(n562) );
  ivd1_hd U814 ( .A(n562), .Y(n563) );
  ivd1_hd U815 ( .A(z_m[22]), .Y(n564) );
  ivd1_hd U816 ( .A(n564), .Y(n565) );
  ivd1_hd U817 ( .A(z_m[9]), .Y(n566) );
  ivd1_hd U818 ( .A(n566), .Y(n567) );
  ivd1_hd U819 ( .A(z_m[13]), .Y(n568) );
  ivd1_hd U820 ( .A(n568), .Y(n569) );
  ivd1_hd U821 ( .A(z_m[17]), .Y(n570) );
  ivd1_hd U822 ( .A(n570), .Y(n571) );
  ivd1_hd U823 ( .A(n662), .Y(n572) );
  ivd1_hd U824 ( .A(state[1]), .Y(n573) );
  ivd1_hd U825 ( .A(state[1]), .Y(n574) );
  ivd1_hd U826 ( .A(n1110), .Y(n575) );
  ivd1_hd U827 ( .A(n1110), .Y(n576) );
  ivd1_hd U828 ( .A(n1299), .Y(n577) );
  ivd1_hd U829 ( .A(n1299), .Y(n578) );
  ivd1_hd U830 ( .A(n1113), .Y(n579) );
  ivd1_hd U831 ( .A(n1113), .Y(n580) );
  ivd1_hd U832 ( .A(a_m[6]), .Y(n581) );
  ivd1_hd U833 ( .A(n581), .Y(n582) );
  ivd1_hd U834 ( .A(a_m[4]), .Y(n583) );
  ivd1_hd U835 ( .A(n583), .Y(n584) );
  ivd1_hd U836 ( .A(b_m[20]), .Y(n585) );
  ivd1_hd U837 ( .A(n585), .Y(n586) );
  ivd1_hd U838 ( .A(a_m[8]), .Y(n587) );
  ivd1_hd U839 ( .A(n587), .Y(n588) );
  ivd1_hd U840 ( .A(a_m[16]), .Y(n589) );
  ivd1_hd U841 ( .A(n589), .Y(n590) );
  ivd1_hd U842 ( .A(a_m[14]), .Y(n591) );
  ivd1_hd U843 ( .A(n591), .Y(n592) );
  ivd1_hd U844 ( .A(a_m[18]), .Y(n593) );
  ivd1_hd U845 ( .A(n593), .Y(n594) );
  ivd1_hd U846 ( .A(a_m[10]), .Y(n595) );
  ivd1_hd U847 ( .A(n595), .Y(n596) );
  ivd1_hd U848 ( .A(b_m[22]), .Y(n597) );
  ivd1_hd U849 ( .A(n597), .Y(n598) );
  ivd1_hd U850 ( .A(a_m[12]), .Y(n599) );
  ivd1_hd U851 ( .A(n599), .Y(n600) );
  ivd1_hd U852 ( .A(b_m[7]), .Y(n601) );
  ivd1_hd U853 ( .A(n601), .Y(n602) );
  ivd1_hd U854 ( .A(a_m[20]), .Y(n603) );
  ivd1_hd U855 ( .A(n603), .Y(n604) );
  ivd1_hd U856 ( .A(a_m[15]), .Y(n605) );
  ivd1_hd U857 ( .A(n605), .Y(n606) );
  ivd1_hd U858 ( .A(b_m[12]), .Y(n607) );
  ivd1_hd U859 ( .A(n607), .Y(n608) );
  ivd1_hd U860 ( .A(b_m[23]), .Y(n609) );
  ivd1_hd U861 ( .A(n609), .Y(n610) );
  ivd1_hd U862 ( .A(b_m[24]), .Y(n611) );
  ivd1_hd U863 ( .A(n611), .Y(n612) );
  ivd1_hd U864 ( .A(z_m[5]), .Y(n613) );
  ivd1_hd U865 ( .A(n613), .Y(n614) );
  ivd1_hd U866 ( .A(n575), .Y(n615) );
  ivd1_hd U867 ( .A(n672), .Y(n616) );
  ivd1_hd U868 ( .A(n804), .Y(n617) );
  ivd1_hd U869 ( .A(n804), .Y(n618) );
  ivd1_hd U870 ( .A(n1118), .Y(n619) );
  ivd1_hd U871 ( .A(n1118), .Y(n620) );
  ivd1_hd U872 ( .A(n628), .Y(n621) );
  ivd1_hd U873 ( .A(n628), .Y(n622) );
  ivd1_hd U874 ( .A(n654), .Y(n623) );
  ivd1_hd U875 ( .A(n654), .Y(n624) );
  ivd1_hd U876 ( .A(n1376), .Y(n625) );
  ivd1_hd U877 ( .A(n1376), .Y(n626) );
  ivd1_hd U878 ( .A(n1376), .Y(n627) );
  ivd1_hd U879 ( .A(n955), .Y(n628) );
  ivd1_hd U880 ( .A(n955), .Y(n629) );
  ivd1_hd U881 ( .A(n955), .Y(n630) );
  ivd1_hd U882 ( .A(n1163), .Y(n631) );
  ivd1_hd U883 ( .A(n631), .Y(n632) );
  ivd1_hd U884 ( .A(n631), .Y(n633) );
  ivd1_hd U885 ( .A(n631), .Y(n634) );
  ivd1_hd U886 ( .A(n131), .Y(n635) );
  ivd1_hd U887 ( .A(n131), .Y(n636) );
  ivd1_hd U888 ( .A(n1164), .Y(n637) );
  ivd1_hd U889 ( .A(n1164), .Y(n638) );
  ivd1_hd U890 ( .A(n1164), .Y(n639) );
  ivd1_hd U891 ( .A(n1164), .Y(n640) );
  ivd1_hd U892 ( .A(n1253), .Y(n641) );
  ivd1_hd U893 ( .A(n1253), .Y(n642) );
  ivd1_hd U894 ( .A(n1253), .Y(n643) );
  ivd1_hd U895 ( .A(n1253), .Y(n644) );
  nid1_hd U896 ( .A(n1373), .Y(n645) );
  ivd1_hd U897 ( .A(a_e[7]), .Y(n646) );
  nid1_hd U898 ( .A(n1365), .Y(n647) );
  nid1_hd U899 ( .A(b_e[6]), .Y(n648) );
  ivd1_hd U900 ( .A(n1270), .Y(n649) );
  nid1_hd U901 ( .A(n1200), .Y(n650) );
  ivd1_hd U902 ( .A(n743), .Y(n651) );
  ivd1_hd U903 ( .A(n1010), .Y(n652) );
  ivd1_hd U904 ( .A(n1004), .Y(n653) );
  nid1_hd U905 ( .A(n1389), .Y(n654) );
  nid1_hd U906 ( .A(n1389), .Y(n655) );
  nid1_hd U907 ( .A(n1389), .Y(n656) );
  scg16d1_hd U908 ( .A(n1248), .B(n1247), .C(n626), .Y(n1389) );
  nid1_hd U909 ( .A(n619), .Y(n1128) );
  ivd1_hd U910 ( .A(n1128), .Y(n657) );
  ivd1_hd U911 ( .A(n1128), .Y(n658) );
  ivd1_hd U912 ( .A(n1128), .Y(n659) );
  ivd1_hd U913 ( .A(n1255), .Y(n660) );
  ivd1_hd U914 ( .A(n1255), .Y(n661) );
  ivd1_hd U915 ( .A(n1255), .Y(n662) );
  ivd1_hd U916 ( .A(n1255), .Y(n663) );
  or2d1_hd U917 ( .A(n1168), .B(n1158), .Y(n1165) );
  ivd1_hd U918 ( .A(n1165), .Y(n664) );
  ivd1_hd U919 ( .A(n1165), .Y(n665) );
  ivd1_hd U920 ( .A(n1165), .Y(n666) );
  ivd1_hd U921 ( .A(n1165), .Y(n667) );
  ivd1_hd U922 ( .A(n579), .Y(n668) );
  ivd1_hd U923 ( .A(n579), .Y(n669) );
  ivd1_hd U924 ( .A(n579), .Y(n670) );
  ivd1_hd U925 ( .A(n1260), .Y(n671) );
  ad2d1_hd U926 ( .A(n615), .B(n636), .Y(n1144) );
  ivd1_hd U927 ( .A(n1144), .Y(n672) );
  ivd1_hd U928 ( .A(n1144), .Y(n673) );
  ivd1_hd U929 ( .A(n1144), .Y(n674) );
  or2d1_hd U930 ( .A(n1257), .B(n574), .Y(DP_OP_154J1_137_6175_n25) );
  ivd1_hd U931 ( .A(DP_OP_154J1_137_6175_n25), .Y(n675) );
  ivd1_hd U932 ( .A(DP_OP_154J1_137_6175_n25), .Y(n676) );
  ivd1_hd U933 ( .A(DP_OP_154J1_137_6175_n25), .Y(n677) );
  ivd1_hd U934 ( .A(n705), .Y(n700) );
  ivd1_hd U935 ( .A(n706), .Y(n696) );
  ivd1_hd U936 ( .A(n706), .Y(n697) );
  ivd1_hd U937 ( .A(n1004), .Y(n805) );
  nr2d1_hd U938 ( .A(n816), .B(n904), .Y(n1358) );
  ivd1_hd U939 ( .A(n125), .Y(n724) );
  ivd1_hd U940 ( .A(n678), .Y(n698) );
  ivd1_hd U941 ( .A(n678), .Y(n703) );
  ivd1_hd U942 ( .A(n627), .Y(RSOP_150_C1_CONTROL1) );
  ivd1_hd U943 ( .A(n1358), .Y(n1260) );
  ivd1_hd U944 ( .A(n1010), .Y(n18) );
  ivd1_hd U945 ( .A(n1155), .Y(n1152) );
  nr2d1_hd U946 ( .A(n1250), .B(n724), .Y(n1199) );
  ivd1_hd U947 ( .A(n93), .Y(n1250) );
  ivd1_hd U948 ( .A(n705), .Y(n699) );
  ivd1_hd U949 ( .A(n641), .Y(n994) );
  ivd1_hd U950 ( .A(n718), .Y(n716) );
  ivd1_hd U951 ( .A(n718), .Y(n717) );
  ivd1_hd U952 ( .A(n1379), .Y(n1365) );
  ivd1_hd U953 ( .A(n995), .Y(n817) );
  ivd1_hd U954 ( .A(n1025), .Y(n1151) );
  ivd1_hd U955 ( .A(n125), .Y(n723) );
  ivd1_hd U956 ( .A(n1199), .Y(n783) );
  nd2bd1_hd U957 ( .AN(n896), .B(n679), .Y(n1210) );
  nr2d1_hd U958 ( .A(n1391), .B(n1159), .Y(n814) );
  ivd1_hd U959 ( .A(n706), .Y(n695) );
  nd3d1_hd U960 ( .A(n104), .B(i_AB_STB), .C(o_AB_ACK), .Y(n103) );
  scg12d1_hd U961 ( .A(state[3]), .B(n1243), .C(n574), .Y(n509) );
  ivd1_hd U962 ( .A(n1390), .Y(n1387) );
  ivd1_hd U963 ( .A(a_e[1]), .Y(n1329) );
  nr2d1_hd U964 ( .A(n1250), .B(n1157), .Y(n1390) );
  ivd1_hd U965 ( .A(n125), .Y(n725) );
  ivd1_hd U966 ( .A(n729), .Y(n726) );
  ivd1_hd U967 ( .A(n729), .Y(n727) );
  ivd1_hd U968 ( .A(n1199), .Y(n1168) );
  ivd1_hd U969 ( .A(z_m[23]), .Y(n1145) );
  ivd1_hd U970 ( .A(z_m[0]), .Y(n1217) );
  nd2bd1_hd U971 ( .AN(n995), .B(n740), .Y(n1155) );
  ao22d1_hd U972 ( .A(n1177), .B(n1244), .C(n1199), .D(n1176), .Y(n1200) );
  ivd1_hd U973 ( .A(a_e[3]), .Y(n1343) );
  ivd1_hd U974 ( .A(n1158), .Y(n777) );
  nr2d1_hd U975 ( .A(n897), .B(n896), .Y(n1388) );
  ivd1_hd U976 ( .A(b_e[8]), .Y(n1249) );
  ivd1_hd U977 ( .A(b_e[1]), .Y(n1264) );
  ivd1_hd U978 ( .A(b_e[9]), .Y(n1251) );
  ivd1_hd U979 ( .A(b_e[7]), .Y(n1317) );
  ivd1_hd U980 ( .A(a_e[0]), .Y(n1328) );
  ivd1_hd U981 ( .A(a_e[5]), .Y(n1360) );
  ivd1_hd U982 ( .A(a_e[7]), .Y(n1385) );
  ivd1_hd U983 ( .A(state[3]), .Y(n28) );
  ivd1_hd U984 ( .A(state[2]), .Y(n29) );
  ivd1_hd U985 ( .A(a_m[23]), .Y(n953) );
  ivd1_hd U986 ( .A(b_m[21]), .Y(n990) );
  ivd1_hd U987 ( .A(b_m[16]), .Y(n983) );
  ivd1_hd U988 ( .A(b_m[25]), .Y(n1256) );
  ivd1_hd U989 ( .A(b_m[26]), .Y(n833) );
  scg17d1_hd U990 ( .A(sticky), .B(n1155), .C(n1154), .D(n1153), .Y(n393) );
  scg6d1_hd U991 ( .A(n618), .B(n800), .C(n801), .Y(n427) );
  ivd1_hd U992 ( .A(a[30]), .Y(n1377) );
  nd4d1_hd U993 ( .A(n1003), .B(n1025), .C(n1006), .D(n717), .Y(n1004) );
  ivd1_hd U994 ( .A(n1323), .Y(n1357) );
  oa21d1_hd U995 ( .A(n1391), .B(n1387), .C(n623), .Y(n1323) );
  scg17d1_hd U996 ( .A(b_e[8]), .B(n1320), .C(n1319), .D(n1318), .Y(n490) );
  ivd1_hd U997 ( .A(z_m[6]), .Y(n1221) );
  ivd1_hd U998 ( .A(z_m[14]), .Y(n1229) );
  ivd1_hd U999 ( .A(z_m[18]), .Y(n1225) );
  ivd1_hd U1000 ( .A(z_m[10]), .Y(n1219) );
  ivd1_hd U1001 ( .A(b[30]), .Y(n1310) );
  ivd1_hd U1002 ( .A(b_e[5]), .Y(n1294) );
  ivd1_hd U1003 ( .A(a_e[2]), .Y(n1335) );
  nr2bd1_hd U1004 ( .AN(b_e[6]), .B(a_e[6]), .Y(n916) );
  ivd1_hd U1005 ( .A(z_m[20]), .Y(n1226) );
  ivd1_hd U1006 ( .A(z_m[16]), .Y(n1230) );
  ivd1_hd U1007 ( .A(z_m[15]), .Y(n1231) );
  ivd1_hd U1008 ( .A(z_m[19]), .Y(n1227) );
  ivd1_hd U1009 ( .A(z_m[12]), .Y(n1220) );
  ivd1_hd U1010 ( .A(z_m[8]), .Y(n1222) );
  ivd1_hd U1011 ( .A(z_m[7]), .Y(n1223) );
  ivd1_hd U1012 ( .A(z_m[11]), .Y(n1224) );
  ivd1_hd U1013 ( .A(z_m[4]), .Y(n1215) );
  ivd1_hd U1014 ( .A(z_m[2]), .Y(n1214) );
  nd3d1_hd U1015 ( .A(n675), .B(n1145), .C(n1246), .Y(n1006) );
  nr2d1_hd U1016 ( .A(n28), .B(n1258), .Y(n1010) );
  ivd1_hd U1017 ( .A(state[0]), .Y(n816) );
  nr2d1_hd U1018 ( .A(sum[27]), .B(n1155), .Y(n1146) );
  ivd1_hd U1019 ( .A(z_e[0]), .Y(n800) );
  ivd1_hd U1020 ( .A(z_e[9]), .Y(n1171) );
  ao21d1_hd U1021 ( .A(n1196), .B(n1170), .C(z_e[9]), .Y(n1177) );
  ivd1_hd U1022 ( .A(z_e[8]), .Y(n1170) );
  ivd1_hd U1023 ( .A(z_e[7]), .Y(n1196) );
  ivd1_hd U1024 ( .A(b_e[3]), .Y(n1278) );
  ivd1_hd U1025 ( .A(n1204), .Y(n778) );
  ivd1_hd U1026 ( .A(n1207), .Y(n741) );
  nr2d1_hd U1027 ( .A(n895), .B(n894), .Y(n1160) );
  ivd1_hd U1028 ( .A(b_e[0]), .Y(n1263) );
  ivd1_hd U1029 ( .A(a_e[8]), .Y(n1322) );
  ivd1_hd U1030 ( .A(a_e[6]), .Y(n1005) );
  ivd1_hd U1031 ( .A(a_e[4]), .Y(n1350) );
  nr2d1_hd U1032 ( .A(state[0]), .B(n904), .Y(n93) );
  nd3d1_hd U1033 ( .A(state[1]), .B(n29), .C(n28), .Y(n904) );
  ivd1_hd U1034 ( .A(a_m[25]), .Y(n956) );
  ivd1_hd U1035 ( .A(n836), .Y(n835) );
  ivd1_hd U1036 ( .A(b_m[9]), .Y(n972) );
  ivd1_hd U1037 ( .A(a_m[5]), .Y(n932) );
  ivd1_hd U1038 ( .A(b_m[3]), .Y(n963) );
  ivd1_hd U1039 ( .A(a_m[3]), .Y(n929) );
  ivd1_hd U1040 ( .A(a_m[2]), .Y(n927) );
  ivd1_hd U1041 ( .A(a_m[1]), .Y(n926) );
  ivd1_hd U1042 ( .A(b_m[4]), .Y(n965) );
  ivd1_hd U1043 ( .A(b_m[6]), .Y(n968) );
  ivd1_hd U1044 ( .A(a_m[7]), .Y(n935) );
  ivd1_hd U1045 ( .A(b_m[10]), .Y(n974) );
  ivd1_hd U1046 ( .A(b_m[15]), .Y(n981) );
  ivd1_hd U1047 ( .A(b_m[13]), .Y(n978) );
  ivd1_hd U1048 ( .A(a_m[17]), .Y(n946) );
  ivd1_hd U1049 ( .A(b_m[18]), .Y(n986) );
  ivd1_hd U1050 ( .A(b_m[1]), .Y(n960) );
  ivd1_hd U1051 ( .A(b_m[2]), .Y(n961) );
  nr2d1_hd U1052 ( .A(state[3]), .B(n1258), .Y(n104) );
  nr2d1_hd U1053 ( .A(n676), .B(n1152), .Y(n785) );
  nr2d1_hd U1054 ( .A(n1010), .B(n635), .Y(n812) );
  nr2d1_hd U1055 ( .A(n1156), .B(state[3]), .Y(n1245) );
  nr2d1_hd U1056 ( .A(n1249), .B(a_e[8]), .Y(n920) );
  nr2d1_hd U1057 ( .A(state[2]), .B(state[0]), .Y(n1243) );
  nr2d1_hd U1058 ( .A(n1317), .B(b_e[6]), .Y(n822) );
  ivd1_hd U1059 ( .A(a_e[9]), .Y(n1324) );
  ao22d1_hd U1060 ( .A(n835), .B(n834), .C(a_m[26]), .D(n833), .Y(n885) );
  oa22d1_hd U1061 ( .A(n833), .B(a_m[26]), .C(n1256), .D(a_m[25]), .Y(n836) );
  oa211d1_hd U1062 ( .A(n717), .B(n1005), .C(n789), .D(n788), .Y(n421) );
  oa211d1_hd U1063 ( .A(n716), .B(n1350), .C(n793), .D(n792), .Y(n423) );
  oa211d1_hd U1064 ( .A(n717), .B(n1360), .C(n791), .D(n790), .Y(n422) );
  oa211d1_hd U1065 ( .A(n716), .B(n1335), .C(n797), .D(n796), .Y(n425) );
  oa211d1_hd U1066 ( .A(n716), .B(n1343), .C(n795), .D(n794), .Y(n424) );
  oa211d1_hd U1067 ( .A(n716), .B(n1329), .C(n799), .D(n798), .Y(n426) );
  oa211d1_hd U1068 ( .A(n716), .B(n646), .C(n787), .D(n786), .Y(n420) );
  oa211d1_hd U1069 ( .A(n1322), .B(n716), .C(n807), .D(n806), .Y(n419) );
  oa211d1_hd U1070 ( .A(n1004), .B(n1171), .C(n803), .D(n802), .Y(n428) );
  nr2d1_hd U1071 ( .A(n1171), .B(n820), .Y(N394) );
  ivd1_hd U1072 ( .A(n1156), .Y(n740) );
  oa211d1_hd U1073 ( .A(n783), .B(n748), .C(n1200), .D(n744), .Y(n369) );
  oa211d1_hd U1074 ( .A(n783), .B(n761), .C(n1200), .D(n760), .Y(n366) );
  oa211d1_hd U1075 ( .A(n784), .B(n783), .C(n1200), .D(n782), .Y(n362) );
  oa211d1_hd U1076 ( .A(n783), .B(n751), .C(n1200), .D(n750), .Y(n368) );
  oa211d1_hd U1077 ( .A(n783), .B(n771), .C(n650), .D(n770), .Y(n364) );
  ivd1_hd U1078 ( .A(a_e[0]), .Y(n742) );
  nr2d1_hd U1079 ( .A(n814), .B(n1176), .Y(n813) );
  ivd1_hd U1080 ( .A(n1210), .Y(n1206) );
  oa22d1_hd U1081 ( .A(n1004), .B(n800), .C(n717), .D(n1328), .Y(n801) );
  ivd1_hd U1082 ( .A(n729), .Y(n728) );
  ivd1_hd U1083 ( .A(a_s), .Y(n886) );
  ivd1_hd U1084 ( .A(b_s), .Y(n1208) );
  ivd1_hd U1085 ( .A(n678), .Y(n704) );
  scg17d1_hd U1086 ( .A(n1199), .B(n766), .C(n765), .D(n650), .Y(n365) );
  oa22d1_hd U1087 ( .A(n125), .B(n764), .C(n1201), .D(n1188), .Y(n765) );
  ivd1_hd U1088 ( .A(z[27]), .Y(n764) );
  oa21d1_hd U1089 ( .A(n763), .B(n762), .C(n768), .Y(n766) );
  scg17d1_hd U1090 ( .A(n1199), .B(n756), .C(n755), .D(n650), .Y(n367) );
  oa22d1_hd U1091 ( .A(n729), .B(n754), .C(n1201), .D(n1182), .Y(n755) );
  ivd1_hd U1092 ( .A(z[25]), .Y(n754) );
  oa21d1_hd U1093 ( .A(n753), .B(n752), .C(n758), .Y(n756) );
  scg17d1_hd U1094 ( .A(n1199), .B(n776), .C(n775), .D(n650), .Y(n363) );
  oa22d1_hd U1095 ( .A(n125), .B(n774), .C(n1201), .D(n1195), .Y(n775) );
  ivd1_hd U1096 ( .A(z[29]), .Y(n774) );
  oa21d1_hd U1097 ( .A(n773), .B(n772), .C(n779), .Y(n776) );
  ao22d1_hd U1098 ( .A(n723), .B(z[23]), .C(n743), .D(n800), .Y(n744) );
  ivd1_hd U1099 ( .A(n1201), .Y(n743) );
  ao21d1_hd U1100 ( .A(n723), .B(z[26]), .C(n759), .Y(n760) );
  nr2d1_hd U1101 ( .A(n651), .B(n1186), .Y(n759) );
  ao21d1_hd U1102 ( .A(n758), .B(n757), .C(n763), .Y(n761) );
  ao21d1_hd U1103 ( .A(n723), .B(z[30]), .C(n781), .Y(n782) );
  nr2d1_hd U1104 ( .A(n1202), .B(n651), .Y(n781) );
  ao22d1_hd U1105 ( .A(n778), .B(a_e[6]), .C(n777), .D(n648), .Y(n772) );
  ao22d1_hd U1106 ( .A(n778), .B(a_e[7]), .C(n777), .D(b_e[7]), .Y(n780) );
  ao21d1_hd U1107 ( .A(n723), .B(z[24]), .C(n749), .Y(n750) );
  nr2d1_hd U1108 ( .A(n651), .B(n1180), .Y(n749) );
  ao21d1_hd U1109 ( .A(n748), .B(n747), .C(n753), .Y(n751) );
  ao21d1_hd U1110 ( .A(n723), .B(z[28]), .C(n769), .Y(n770) );
  nr2d1_hd U1111 ( .A(n1192), .B(n651), .Y(n769) );
  ao21d1_hd U1112 ( .A(n768), .B(n767), .C(n773), .Y(n771) );
  nr2d1_hd U1113 ( .A(n768), .B(n767), .Y(n773) );
  ao22d1_hd U1114 ( .A(n778), .B(a_e[4]), .C(n777), .D(b_e[4]), .Y(n762) );
  nr2d1_hd U1115 ( .A(n758), .B(n757), .Y(n763) );
  oa22d1_hd U1116 ( .A(n1204), .B(n1343), .C(n1158), .D(n1278), .Y(n757) );
  ao22d1_hd U1117 ( .A(n778), .B(a_e[2]), .C(n777), .D(b_e[2]), .Y(n752) );
  nr2d1_hd U1118 ( .A(n748), .B(n747), .Y(n753) );
  oa22d1_hd U1119 ( .A(n1204), .B(n746), .C(n1158), .D(n745), .Y(n747) );
  ivd1_hd U1120 ( .A(b_e[1]), .Y(n745) );
  ivd1_hd U1121 ( .A(a_e[1]), .Y(n746) );
  oa22d1_hd U1122 ( .A(n1204), .B(n742), .C(n1158), .D(n1263), .Y(n748) );
  ivd1_hd U1123 ( .A(z_e[1]), .Y(n1178) );
  nr2d1_hd U1124 ( .A(z_e[6]), .B(z_e[5]), .Y(n818) );
  ivd1_hd U1125 ( .A(z_e[4]), .Y(n1189) );
  nr2d1_hd U1126 ( .A(n1172), .B(n1173), .Y(n819) );
  ao21d1_hd U1127 ( .A(n1178), .B(n819), .C(n1001), .Y(n820) );
  nr4d1_hd U1128 ( .A(b_e[3]), .B(b_e[2]), .C(b_e[4]), .D(b_e[5]), .Y(n821) );
  nd3d1_hd U1129 ( .A(n1350), .B(n1360), .C(n1005), .Y(n823) );
  nr2d1_hd U1130 ( .A(n1385), .B(n824), .Y(n898) );
  nd4d1_hd U1131 ( .A(a_e[0]), .B(a_e[9]), .C(a_e[8]), .D(n898), .Y(n1391) );
  nr4d1_hd U1132 ( .A(n541), .B(n590), .C(a_m[23]), .D(n549), .Y(n832) );
  nr4d1_hd U1133 ( .A(n555), .B(a_m[17]), .C(a_m[7]), .D(a_m[15]), .Y(n831) );
  nr3d1_hd U1134 ( .A(n604), .B(a_m[25]), .C(n561), .Y(n830) );
  nr4d1_hd U1135 ( .A(a_m[0]), .B(n584), .C(a_m[1]), .D(a_m[2]), .Y(n828) );
  nr4d1_hd U1136 ( .A(n596), .B(a_m[5]), .C(a_m[3]), .D(a_m[26]), .Y(n827) );
  nr4d1_hd U1137 ( .A(n553), .B(a_m[11]), .C(n588), .D(a_m[18]), .Y(n826) );
  nr4d1_hd U1138 ( .A(n582), .B(n600), .C(n592), .D(n547), .Y(n825) );
  nd4d1_hd U1139 ( .A(n832), .B(n831), .C(n830), .D(n829), .Y(n1159) );
  oa22d1_hd U1140 ( .A(b_m[25]), .B(n956), .C(n612), .D(n560), .Y(n834) );
  ao21d1_hd U1141 ( .A(n612), .B(n560), .C(n836), .Y(n883) );
  oa211d1_hd U1142 ( .A(n594), .B(n986), .C(n838), .D(n837), .Y(n881) );
  nr2d1_hd U1143 ( .A(n555), .B(n990), .Y(n871) );
  ao211d1_hd U1144 ( .A(n586), .B(n603), .C(n871), .D(n873), .Y(n878) );
  nr2d1_hd U1145 ( .A(n547), .B(n978), .Y(n858) );
  nr2d1_hd U1146 ( .A(n608), .B(n858), .Y(n839) );
  ao22d1_hd U1147 ( .A(n839), .B(n600), .C(n547), .D(n978), .Y(n866) );
  oa22d1_hd U1148 ( .A(n606), .B(n981), .C(n592), .D(n550), .Y(n865) );
  nr2d1_hd U1149 ( .A(a_m[15]), .B(n981), .Y(n840) );
  nr2d1_hd U1150 ( .A(n551), .B(n840), .Y(n841) );
  ao22d1_hd U1151 ( .A(n841), .B(n592), .C(n606), .D(n981), .Y(n864) );
  oa22d1_hd U1152 ( .A(n542), .B(n539), .C(n974), .D(n596), .Y(n856) );
  ivd1_hd U1153 ( .A(n856), .Y(n853) );
  ao22d1_hd U1154 ( .A(b_m[1]), .B(n926), .C(b_m[2]), .D(n927), .Y(n844) );
  ivd1_hd U1155 ( .A(a_m[0]), .Y(n925) );
  oa211d1_hd U1156 ( .A(b_m[1]), .B(n926), .C(b_m[0]), .D(n925), .Y(n843) );
  oa22d1_hd U1157 ( .A(b_m[3]), .B(n929), .C(b_m[2]), .D(n927), .Y(n842) );
  ao21d1_hd U1158 ( .A(n844), .B(n843), .C(n842), .Y(n846) );
  oa22d1_hd U1159 ( .A(a_m[3]), .B(n963), .C(n584), .D(n965), .Y(n845) );
  oa22d1_hd U1160 ( .A(n846), .B(n845), .C(n537), .D(n932), .Y(n847) );
  ao21d1_hd U1161 ( .A(n584), .B(n965), .C(n847), .Y(n849) );
  oa22d1_hd U1162 ( .A(a_m[5]), .B(n536), .C(n582), .D(n968), .Y(n848) );
  oa22d1_hd U1163 ( .A(n849), .B(n848), .C(n602), .D(n935), .Y(n850) );
  ao21d1_hd U1164 ( .A(n582), .B(n968), .C(n850), .Y(n851) );
  nr2d1_hd U1165 ( .A(n553), .B(n972), .Y(n854) );
  ao211d1_hd U1166 ( .A(n602), .B(n935), .C(n851), .D(n854), .Y(n852) );
  oa211d1_hd U1167 ( .A(n588), .B(n544), .C(n853), .D(n852), .Y(n862) );
  oa211d1_hd U1168 ( .A(n539), .B(n542), .C(n596), .D(n974), .Y(n861) );
  nr2d1_hd U1169 ( .A(n545), .B(n854), .Y(n855) );
  ao22d1_hd U1170 ( .A(n855), .B(n588), .C(n553), .D(n972), .Y(n857) );
  oa22d1_hd U1171 ( .A(n543), .B(n538), .C(n857), .D(n856), .Y(n860) );
  ao211d1_hd U1172 ( .A(n608), .B(n599), .C(n858), .D(n865), .Y(n859) );
  scg22d1_hd U1173 ( .A(n862), .B(n861), .C(n860), .D(n859), .Y(n863) );
  oa211d1_hd U1174 ( .A(n866), .B(n865), .C(n864), .D(n863), .Y(n867) );
  oa211d1_hd U1175 ( .A(n590), .B(n983), .C(n878), .D(n867), .Y(n880) );
  ao22d1_hd U1176 ( .A(a_m[17]), .B(n556), .C(n590), .D(n983), .Y(n870) );
  oa211d1_hd U1177 ( .A(n549), .B(n558), .C(n594), .D(n986), .Y(n869) );
  oa211d1_hd U1178 ( .A(n870), .B(n881), .C(n869), .D(n868), .Y(n877) );
  ao211d1_hd U1179 ( .A(n610), .B(n953), .C(n598), .D(n540), .Y(n876) );
  nr2d1_hd U1180 ( .A(n586), .B(n871), .Y(n872) );
  ao22d1_hd U1181 ( .A(n872), .B(n604), .C(n555), .D(n990), .Y(n874) );
  oa22d1_hd U1182 ( .A(n610), .B(n953), .C(n874), .D(n873), .Y(n875) );
  ao211d1_hd U1183 ( .A(n878), .B(n877), .C(n876), .D(n875), .Y(n879) );
  oa21d1_hd U1184 ( .A(n881), .B(n880), .C(n879), .Y(n882) );
  ao22d1_hd U1185 ( .A(n704), .B(n1208), .C(n886), .D(n705), .Y(N338) );
  nr4d1_hd U1186 ( .A(b_m[3]), .B(n608), .C(b_m[5]), .D(n602), .Y(n890) );
  nr4d1_hd U1187 ( .A(b_m[6]), .B(b_m[1]), .C(b_m[0]), .D(b_m[2]), .Y(n889) );
  nr4d1_hd U1188 ( .A(b_m[26]), .B(n612), .C(b_m[25]), .D(b_m[18]), .Y(n888)
         );
  nr4d1_hd U1189 ( .A(n551), .B(b_m[15]), .C(b_m[10]), .D(b_m[8]), .Y(n887) );
  nd4d1_hd U1190 ( .A(n890), .B(n889), .C(n888), .D(n887), .Y(n895) );
  nr4d1_hd U1191 ( .A(b_m[16]), .B(b_m[17]), .C(n598), .D(n586), .Y(n893) );
  nr2d1_hd U1192 ( .A(b_m[23]), .B(b_m[19]), .Y(n892) );
  nr4d1_hd U1193 ( .A(b_m[13]), .B(n543), .C(b_m[4]), .D(b_m[9]), .Y(n891) );
  nd4d1_hd U1194 ( .A(n893), .B(n892), .C(n891), .D(n990), .Y(n894) );
  nd4d1_hd U1195 ( .A(b_e[9]), .B(b_e[0]), .C(b_e[8]), .D(n1264), .Y(n897) );
  nd4d1_hd U1196 ( .A(n898), .B(n1328), .C(n1324), .D(n1322), .Y(n1205) );
  nr2d1_hd U1197 ( .A(n1264), .B(a_e[1]), .Y(n899) );
  nr2d1_hd U1198 ( .A(n1294), .B(a_e[5]), .Y(n909) );
  nr4d1_hd U1199 ( .A(n899), .B(n909), .C(n920), .D(n916), .Y(n903) );
  ivd1_hd U1200 ( .A(b_e[4]), .Y(n1285) );
  nr2d1_hd U1201 ( .A(n1285), .B(a_e[4]), .Y(n910) );
  ivd1_hd U1202 ( .A(n910), .Y(n900) );
  nd4d1_hd U1203 ( .A(n922), .B(n905), .C(n903), .D(n902), .Y(n1248) );
  ao22d1_hd U1204 ( .A(a_e[3]), .B(n1278), .C(a_e[4]), .D(n1285), .Y(n912) );
  ao211d1_hd U1205 ( .A(b_e[1]), .B(n1329), .C(b_e[0]), .D(n1328), .Y(n908) );
  oa22d1_hd U1206 ( .A(b_e[2]), .B(n1335), .C(b_e[1]), .D(n1329), .Y(n907) );
  oa211d1_hd U1207 ( .A(n908), .B(n907), .C(n906), .D(n905), .Y(n911) );
  ao211d1_hd U1208 ( .A(n912), .B(n911), .C(n910), .D(n909), .Y(n914) );
  oa22d1_hd U1209 ( .A(b_e[5]), .B(n1360), .C(b_e[6]), .D(n1005), .Y(n913) );
  nr2d1_hd U1210 ( .A(n914), .B(n913), .Y(n915) );
  oa22d1_hd U1211 ( .A(n916), .B(n915), .C(b_e[7]), .D(n1385), .Y(n918) );
  ao22d1_hd U1212 ( .A(a_e[8]), .B(n1249), .C(n918), .D(n917), .Y(n919) );
  oa22d1_hd U1213 ( .A(n920), .B(n919), .C(a_e[9]), .D(n1251), .Y(n921) );
  nr2d1_hd U1214 ( .A(n1328), .B(n1329), .Y(n1332) );
  nr2d1_hd U1215 ( .A(n1343), .B(n1342), .Y(n1347) );
  nr2d1_hd U1216 ( .A(n1360), .B(n1359), .Y(n1364) );
  ao21d1_hd U1217 ( .A(n1358), .B(n1378), .C(n1357), .Y(n1386) );
  oa21d1_hd U1218 ( .A(a_e[7]), .B(n1379), .C(n1386), .Y(n1321) );
  nr4d1_hd U1219 ( .A(a_e[8]), .B(n1385), .C(n1379), .D(n1378), .Y(n923) );
  ivd1_hd U1220 ( .A(a[25]), .Y(n1333) );
  nr2d1_hd U1221 ( .A(n1334), .B(n1333), .Y(n1344) );
  ivd1_hd U1222 ( .A(a[27]), .Y(n1348) );
  nr2d1_hd U1223 ( .A(n1349), .B(n1348), .Y(n1361) );
  ivd1_hd U1224 ( .A(a[29]), .Y(n1366) );
  nr2d1_hd U1225 ( .A(n1367), .B(n1366), .Y(n1382) );
  nr2d1_hd U1226 ( .A(n1382), .B(n626), .Y(n1372) );
  scg17d1_hd U1227 ( .A(a_e[8]), .B(n1321), .C(n923), .D(n1383), .Y(n480) );
  ao22d1_hd U1228 ( .A(RSOP_150_C1_CONTROL1), .B(a[22]), .C(a_m[26]), .D(n621), 
        .Y(n924) );
  oa21d1_hd U1229 ( .A(n654), .B(n956), .C(n924), .Y(n479) );
  nr2d1_hd U1230 ( .A(n671), .B(n627), .Y(n959) );
  oa22d1_hd U1231 ( .A(n959), .B(n925), .C(n926), .D(n628), .Y(n478) );
  oa22d1_hd U1232 ( .A(n656), .B(n926), .C(n927), .D(n630), .Y(n477) );
  oa22d1_hd U1233 ( .A(n655), .B(n927), .C(n929), .D(n629), .Y(n476) );
  ao22d1_hd U1234 ( .A(n737), .B(a[0]), .C(a_m[4]), .D(n622), .Y(n928) );
  oa21d1_hd U1235 ( .A(n654), .B(n929), .C(n928), .Y(n475) );
  ao22d1_hd U1236 ( .A(n737), .B(a[1]), .C(n624), .D(n584), .Y(n930) );
  oa21d1_hd U1237 ( .A(n932), .B(n630), .C(n930), .Y(n474) );
  ao22d1_hd U1238 ( .A(n737), .B(a[2]), .C(a_m[6]), .D(n621), .Y(n931) );
  oa21d1_hd U1239 ( .A(n656), .B(n932), .C(n931), .Y(n473) );
  ao22d1_hd U1240 ( .A(n737), .B(a[3]), .C(n623), .D(n582), .Y(n933) );
  oa21d1_hd U1241 ( .A(n935), .B(n629), .C(n933), .Y(n472) );
  ao22d1_hd U1242 ( .A(n737), .B(a[4]), .C(a_m[8]), .D(n622), .Y(n934) );
  oa21d1_hd U1243 ( .A(n655), .B(n935), .C(n934), .Y(n471) );
  ao22d1_hd U1244 ( .A(n737), .B(a[5]), .C(n623), .D(n588), .Y(n936) );
  oa21d1_hd U1245 ( .A(n552), .B(n628), .C(n936), .Y(n470) );
  ao22d1_hd U1246 ( .A(n731), .B(a[6]), .C(a_m[10]), .D(n621), .Y(n937) );
  oa21d1_hd U1247 ( .A(n656), .B(n552), .C(n937), .Y(n469) );
  ao22d1_hd U1248 ( .A(n731), .B(a[7]), .C(n624), .D(n596), .Y(n938) );
  oa21d1_hd U1249 ( .A(n538), .B(n630), .C(n938), .Y(n468) );
  ao22d1_hd U1250 ( .A(n739), .B(a[8]), .C(a_m[12]), .D(n622), .Y(n939) );
  oa21d1_hd U1251 ( .A(n655), .B(n538), .C(n939), .Y(n467) );
  ao22d1_hd U1252 ( .A(n731), .B(a[9]), .C(n624), .D(n600), .Y(n940) );
  oa21d1_hd U1253 ( .A(n546), .B(n629), .C(n940), .Y(n466) );
  ao22d1_hd U1254 ( .A(n739), .B(a[10]), .C(a_m[14]), .D(n621), .Y(n941) );
  oa21d1_hd U1255 ( .A(n656), .B(n546), .C(n941), .Y(n465) );
  ao22d1_hd U1256 ( .A(n739), .B(a[11]), .C(n624), .D(n592), .Y(n942) );
  oa21d1_hd U1257 ( .A(n605), .B(n628), .C(n942), .Y(n464) );
  ao22d1_hd U1258 ( .A(n736), .B(a[12]), .C(a_m[16]), .D(n622), .Y(n943) );
  oa21d1_hd U1259 ( .A(n655), .B(n605), .C(n943), .Y(n463) );
  ao22d1_hd U1260 ( .A(n736), .B(a[13]), .C(n623), .D(n590), .Y(n944) );
  oa21d1_hd U1261 ( .A(n946), .B(n630), .C(n944), .Y(n462) );
  ao22d1_hd U1262 ( .A(n736), .B(a[14]), .C(a_m[18]), .D(n621), .Y(n945) );
  oa21d1_hd U1263 ( .A(n656), .B(n946), .C(n945), .Y(n461) );
  ao22d1_hd U1264 ( .A(n736), .B(a[15]), .C(n623), .D(n594), .Y(n947) );
  oa21d1_hd U1265 ( .A(n548), .B(n629), .C(n947), .Y(n460) );
  ao22d1_hd U1266 ( .A(n736), .B(a[16]), .C(n604), .D(n622), .Y(n948) );
  oa21d1_hd U1267 ( .A(n655), .B(n548), .C(n948), .Y(n459) );
  ao22d1_hd U1268 ( .A(n736), .B(a[17]), .C(n624), .D(a_m[20]), .Y(n949) );
  oa21d1_hd U1269 ( .A(n554), .B(n628), .C(n949), .Y(n458) );
  ao22d1_hd U1270 ( .A(n735), .B(a[18]), .C(n541), .D(n621), .Y(n950) );
  oa21d1_hd U1271 ( .A(n656), .B(n554), .C(n950), .Y(n457) );
  ao22d1_hd U1272 ( .A(n735), .B(a[19]), .C(n624), .D(a_m[22]), .Y(n951) );
  oa21d1_hd U1273 ( .A(n953), .B(n630), .C(n951), .Y(n456) );
  ao22d1_hd U1274 ( .A(n735), .B(a[20]), .C(n561), .D(n622), .Y(n952) );
  oa21d1_hd U1275 ( .A(n655), .B(n953), .C(n952), .Y(n455) );
  ao22d1_hd U1276 ( .A(n735), .B(a[21]), .C(n623), .D(a_m[24]), .Y(n954) );
  oa21d1_hd U1277 ( .A(n956), .B(n629), .C(n954), .Y(n454) );
  ivd1_hd U1278 ( .A(b_m[0]), .Y(n958) );
  oa22d1_hd U1279 ( .A(n959), .B(n958), .C(n960), .D(n994), .Y(n453) );
  oa22d1_hd U1280 ( .A(n960), .B(n663), .C(n961), .D(n994), .Y(n452) );
  oa22d1_hd U1281 ( .A(n961), .B(n662), .C(n963), .D(n994), .Y(n451) );
  ao22d1_hd U1282 ( .A(n735), .B(b[0]), .C(b_m[4]), .D(n644), .Y(n962) );
  oa21d1_hd U1283 ( .A(n963), .B(n661), .C(n962), .Y(n450) );
  ao22d1_hd U1284 ( .A(n734), .B(b[1]), .C(b_m[5]), .D(n641), .Y(n964) );
  oa21d1_hd U1285 ( .A(n965), .B(n660), .C(n964), .Y(n449) );
  ao22d1_hd U1286 ( .A(n734), .B(b[2]), .C(b_m[6]), .D(n641), .Y(n966) );
  oa21d1_hd U1287 ( .A(n536), .B(n663), .C(n966), .Y(n448) );
  ao22d1_hd U1288 ( .A(n734), .B(b[3]), .C(b_m[7]), .D(n642), .Y(n967) );
  oa21d1_hd U1289 ( .A(n968), .B(n662), .C(n967), .Y(n447) );
  ao22d1_hd U1290 ( .A(n734), .B(b[4]), .C(b_m[8]), .D(n644), .Y(n969) );
  scg14d1_hd U1291 ( .A(b_m[7]), .B(n1255), .C(n969), .Y(n446) );
  ao22d1_hd U1292 ( .A(n734), .B(b[5]), .C(b_m[9]), .D(n643), .Y(n970) );
  oa21d1_hd U1293 ( .A(n544), .B(n661), .C(n970), .Y(n445) );
  ao22d1_hd U1294 ( .A(n734), .B(b[6]), .C(b_m[10]), .D(n641), .Y(n971) );
  oa21d1_hd U1295 ( .A(n972), .B(n660), .C(n971), .Y(n444) );
  ao22d1_hd U1296 ( .A(n733), .B(b[7]), .C(b_m[11]), .D(n643), .Y(n973) );
  oa21d1_hd U1297 ( .A(n974), .B(n663), .C(n973), .Y(n443) );
  ao22d1_hd U1298 ( .A(n733), .B(b[8]), .C(b_m[12]), .D(n644), .Y(n975) );
  oa21d1_hd U1299 ( .A(n542), .B(n662), .C(n975), .Y(n442) );
  ao22d1_hd U1300 ( .A(n733), .B(b[9]), .C(b_m[13]), .D(n641), .Y(n976) );
  scg14d1_hd U1301 ( .A(b_m[12]), .B(n572), .C(n976), .Y(n441) );
  ao22d1_hd U1302 ( .A(n733), .B(b[10]), .C(n551), .D(n642), .Y(n977) );
  oa21d1_hd U1303 ( .A(n978), .B(n661), .C(n977), .Y(n440) );
  ao22d1_hd U1304 ( .A(n733), .B(b[11]), .C(b_m[15]), .D(n642), .Y(n979) );
  oa21d1_hd U1305 ( .A(n550), .B(n660), .C(n979), .Y(n439) );
  ao22d1_hd U1306 ( .A(n733), .B(b[12]), .C(b_m[16]), .D(n642), .Y(n980) );
  oa21d1_hd U1307 ( .A(n981), .B(n663), .C(n980), .Y(n438) );
  ao22d1_hd U1308 ( .A(n732), .B(b[13]), .C(b_m[17]), .D(n644), .Y(n982) );
  oa21d1_hd U1309 ( .A(n983), .B(n662), .C(n982), .Y(n437) );
  ao22d1_hd U1310 ( .A(n732), .B(b[14]), .C(b_m[18]), .D(n644), .Y(n984) );
  oa21d1_hd U1311 ( .A(n556), .B(n661), .C(n984), .Y(n436) );
  ao22d1_hd U1312 ( .A(n732), .B(b[15]), .C(b_m[19]), .D(n643), .Y(n985) );
  oa21d1_hd U1313 ( .A(n986), .B(n660), .C(n985), .Y(n435) );
  ao22d1_hd U1314 ( .A(n732), .B(b[16]), .C(b_m[20]), .D(n641), .Y(n987) );
  oa21d1_hd U1315 ( .A(n558), .B(n663), .C(n987), .Y(n434) );
  ao22d1_hd U1316 ( .A(n732), .B(b[17]), .C(n586), .D(n572), .Y(n988) );
  oa21d1_hd U1317 ( .A(n990), .B(n994), .C(n988), .Y(n433) );
  ao22d1_hd U1318 ( .A(n735), .B(b[18]), .C(b_m[22]), .D(n643), .Y(n989) );
  oa21d1_hd U1319 ( .A(n990), .B(n662), .C(n989), .Y(n432) );
  ao22d1_hd U1320 ( .A(n732), .B(b[19]), .C(n598), .D(n572), .Y(n991) );
  oa21d1_hd U1321 ( .A(n609), .B(n994), .C(n991), .Y(n431) );
  ao22d1_hd U1322 ( .A(n1376), .B(b[20]), .C(b_m[24]), .D(n642), .Y(n992) );
  oa21d1_hd U1323 ( .A(n609), .B(n661), .C(n992), .Y(n430) );
  ao22d1_hd U1324 ( .A(n739), .B(b[21]), .C(n612), .D(n572), .Y(n993) );
  oa21d1_hd U1325 ( .A(n1256), .B(n994), .C(n993), .Y(n429) );
  nr2d1_hd U1326 ( .A(n1231), .B(n1230), .Y(n1018) );
  nr2d1_hd U1327 ( .A(n1224), .B(n1220), .Y(n1016) );
  nr2d1_hd U1328 ( .A(n1223), .B(n1222), .Y(n1014) );
  nd3d1_hd U1329 ( .A(n1018), .B(n1016), .C(n1014), .Y(n997) );
  ivd1_hd U1330 ( .A(z_m[3]), .Y(n1216) );
  nr2d1_hd U1331 ( .A(n1216), .B(n1215), .Y(n1012) );
  ivd1_hd U1332 ( .A(n1011), .Y(n1035) );
  nd4d1_hd U1333 ( .A(z_m[23]), .B(n1012), .C(z_m[2]), .D(n1035), .Y(n996) );
  nr4d1_hd U1334 ( .A(n1017), .B(n1013), .C(n997), .D(n996), .Y(n1000) );
  nr2d1_hd U1335 ( .A(n1227), .B(n1226), .Y(n1020) );
  nd4d1_hd U1336 ( .A(n565), .B(guard), .C(z_m[21]), .D(n1020), .Y(n998) );
  nr4d1_hd U1337 ( .A(n18), .B(n1015), .C(n1019), .D(n998), .Y(n999) );
  ao22d1_hd U1338 ( .A(n635), .B(N394), .C(n1000), .D(n999), .Y(n1003) );
  ao211d1_hd U1339 ( .A(z_e[1]), .B(z_e[0]), .C(n1172), .D(n1173), .Y(n1002)
         );
  oa21d1_hd U1340 ( .A(n1002), .B(n1001), .C(z_e[9]), .Y(n1246) );
  ao21d1_hd U1341 ( .A(n635), .B(N394), .C(n1152), .Y(n1150) );
  nr2d1_hd U1342 ( .A(round_bit), .B(sticky), .Y(n1008) );
  ivd1_hd U1343 ( .A(guard), .Y(n1007) );
  ao211d1_hd U1344 ( .A(n1008), .B(n1217), .C(n18), .D(n1007), .Y(n1009) );
  nr2d1_hd U1345 ( .A(n1214), .B(n1011), .Y(n1040) );
  nr2d1_hd U1346 ( .A(n1050), .B(n1013), .Y(n1060) );
  nr2d1_hd U1347 ( .A(n1070), .B(n1015), .Y(n1080) );
  nr2d1_hd U1348 ( .A(n1017), .B(n1090), .Y(n1100) );
  nr2d1_hd U1349 ( .A(n1111), .B(n1019), .Y(n1123) );
  ao21d1_hd U1350 ( .A(n657), .B(n1021), .C(n575), .Y(n1134) );
  oa21d1_hd U1351 ( .A(z_m[21]), .B(n619), .C(n1134), .Y(n1141) );
  ao21d1_hd U1352 ( .A(n659), .B(n564), .C(n1141), .Y(n1024) );
  nr2d1_hd U1353 ( .A(n620), .B(n1021), .Y(n1136) );
  oa21d1_hd U1354 ( .A(z_m[23]), .B(n1139), .C(n669), .Y(n1022) );
  ao22d1_hd U1355 ( .A(n1152), .B(sum[26]), .C(n565), .D(n1022), .Y(n1023) );
  oa211d1_hd U1356 ( .A(n1024), .B(n1145), .C(n1023), .D(n1025), .Y(n418) );
  scg4d1_hd U1357 ( .A(n714), .B(sum[3]), .C(n636), .D(z_m[0]), .E(round_bit), 
        .F(n676), .G(n710), .H(sum[2]), .Y(n266) );
  ao22d1_hd U1358 ( .A(n714), .B(sum[4]), .C(z_m[0]), .D(n576), .Y(n1028) );
  ao22d1_hd U1359 ( .A(guard), .B(n580), .C(z_m[1]), .D(n616), .Y(n1027) );
  nd4d1_hd U1360 ( .A(n1028), .B(n1027), .C(n1029), .D(n1026), .Y(n417) );
  nr2d1_hd U1361 ( .A(n563), .B(n620), .Y(n1034) );
  nr2d1_hd U1362 ( .A(n580), .B(n1034), .Y(n1032) );
  ao22d1_hd U1363 ( .A(n713), .B(sum[5]), .C(n710), .D(sum[4]), .Y(n1031) );
  ao22d1_hd U1364 ( .A(z_m[2]), .B(n616), .C(n563), .D(n1033), .Y(n1030) );
  oa211d1_hd U1365 ( .A(n1032), .B(n1217), .C(n1031), .D(n1030), .Y(n416) );
  ao22d1_hd U1366 ( .A(n713), .B(sum[6]), .C(n710), .D(sum[5]), .Y(n1039) );
  ao22d1_hd U1367 ( .A(n579), .B(n563), .C(z_m[3]), .D(n616), .Y(n1038) );
  oa21d1_hd U1368 ( .A(n1034), .B(n1033), .C(z_m[2]), .Y(n1037) );
  nd3d1_hd U1369 ( .A(n659), .B(n1035), .C(n1214), .Y(n1036) );
  nd4d1_hd U1370 ( .A(n1039), .B(n1038), .C(n1037), .D(n1036), .Y(n415) );
  ao22d1_hd U1371 ( .A(n713), .B(sum[7]), .C(n710), .D(sum[6]), .Y(n1043) );
  oa21d1_hd U1372 ( .A(n1040), .B(n18), .C(n1110), .Y(n1044) );
  oa22d1_hd U1373 ( .A(z_m[3]), .B(n1045), .C(n669), .D(n1214), .Y(n1041) );
  ao21d1_hd U1374 ( .A(z_m[3]), .B(n1044), .C(n1041), .Y(n1042) );
  oa211d1_hd U1375 ( .A(n1215), .B(n672), .C(n1043), .D(n1042), .Y(n414) );
  ao21d1_hd U1376 ( .A(n657), .B(n1216), .C(n1044), .Y(n1049) );
  ao22d1_hd U1377 ( .A(n713), .B(sum[8]), .C(n710), .D(sum[7]), .Y(n1048) );
  oa21d1_hd U1378 ( .A(z_m[4]), .B(n1045), .C(n669), .Y(n1046) );
  ao22d1_hd U1379 ( .A(z_m[3]), .B(n1046), .C(z_m[5]), .D(n616), .Y(n1047) );
  oa211d1_hd U1380 ( .A(n1049), .B(n1215), .C(n1048), .D(n1047), .Y(n413) );
  ao22d1_hd U1381 ( .A(n713), .B(sum[9]), .C(n710), .D(sum[8]), .Y(n1053) );
  ao21d1_hd U1382 ( .A(n658), .B(n1050), .C(n575), .Y(n1055) );
  ao22d1_hd U1383 ( .A(n614), .B(n1055), .C(n1054), .D(n613), .Y(n1051) );
  ao21d1_hd U1384 ( .A(n579), .B(z_m[4]), .C(n1051), .Y(n1052) );
  oa211d1_hd U1385 ( .A(n1221), .B(n674), .C(n1053), .D(n1052), .Y(n412) );
  ao22d1_hd U1386 ( .A(n713), .B(sum[10]), .C(n707), .D(sum[9]), .Y(n1059) );
  oa21d1_hd U1387 ( .A(z_m[6]), .B(n1054), .C(n670), .Y(n1057) );
  oa21d1_hd U1388 ( .A(z_m[5]), .B(n619), .C(n1055), .Y(n1056) );
  ao22d1_hd U1389 ( .A(z_m[5]), .B(n1057), .C(z_m[6]), .D(n1056), .Y(n1058) );
  oa211d1_hd U1390 ( .A(n1223), .B(n673), .C(n1059), .D(n1058), .Y(n411) );
  ao22d1_hd U1391 ( .A(n712), .B(sum[11]), .C(n707), .D(sum[10]), .Y(n1063) );
  oa21d1_hd U1392 ( .A(n1060), .B(n652), .C(n615), .Y(n1064) );
  oa22d1_hd U1393 ( .A(z_m[7]), .B(n1065), .C(n670), .D(n1221), .Y(n1061) );
  ao21d1_hd U1394 ( .A(z_m[7]), .B(n1064), .C(n1061), .Y(n1062) );
  oa211d1_hd U1395 ( .A(n1222), .B(n672), .C(n1063), .D(n1062), .Y(n410) );
  ao21d1_hd U1396 ( .A(n658), .B(n1223), .C(n1064), .Y(n1069) );
  ao22d1_hd U1397 ( .A(n712), .B(sum[12]), .C(n1146), .D(sum[11]), .Y(n1068)
         );
  oa21d1_hd U1398 ( .A(z_m[8]), .B(n1065), .C(n668), .Y(n1066) );
  ao22d1_hd U1399 ( .A(n567), .B(n1144), .C(z_m[7]), .D(n1066), .Y(n1067) );
  oa211d1_hd U1400 ( .A(n1069), .B(n1222), .C(n1068), .D(n1067), .Y(n409) );
  ao22d1_hd U1401 ( .A(n712), .B(sum[13]), .C(n707), .D(sum[12]), .Y(n1073) );
  ao21d1_hd U1402 ( .A(n659), .B(n1070), .C(n576), .Y(n1075) );
  ao22d1_hd U1403 ( .A(z_m[9]), .B(n1075), .C(n1074), .D(n566), .Y(n1071) );
  ao21d1_hd U1404 ( .A(n580), .B(z_m[8]), .C(n1071), .Y(n1072) );
  oa211d1_hd U1405 ( .A(n1219), .B(n674), .C(n1073), .D(n1072), .Y(n408) );
  ao22d1_hd U1406 ( .A(n712), .B(sum[14]), .C(n707), .D(sum[13]), .Y(n1079) );
  oa21d1_hd U1407 ( .A(z_m[10]), .B(n1074), .C(n670), .Y(n1077) );
  oa21d1_hd U1408 ( .A(n567), .B(n620), .C(n1075), .Y(n1076) );
  ao22d1_hd U1409 ( .A(z_m[9]), .B(n1077), .C(z_m[10]), .D(n1076), .Y(n1078)
         );
  oa211d1_hd U1410 ( .A(n1224), .B(n673), .C(n1079), .D(n1078), .Y(n407) );
  ao22d1_hd U1411 ( .A(n712), .B(sum[15]), .C(n1146), .D(sum[14]), .Y(n1083)
         );
  oa21d1_hd U1412 ( .A(n1080), .B(n652), .C(n1110), .Y(n1084) );
  oa22d1_hd U1413 ( .A(z_m[11]), .B(n1085), .C(n669), .D(n1219), .Y(n1081) );
  ao21d1_hd U1414 ( .A(z_m[11]), .B(n1084), .C(n1081), .Y(n1082) );
  oa211d1_hd U1415 ( .A(n1220), .B(n672), .C(n1083), .D(n1082), .Y(n406) );
  ao21d1_hd U1416 ( .A(n659), .B(n1224), .C(n1084), .Y(n1089) );
  ao22d1_hd U1417 ( .A(n712), .B(sum[16]), .C(n709), .D(sum[15]), .Y(n1088) );
  oa21d1_hd U1418 ( .A(z_m[12]), .B(n1085), .C(n670), .Y(n1086) );
  ao22d1_hd U1419 ( .A(n569), .B(n616), .C(z_m[11]), .D(n1086), .Y(n1087) );
  oa211d1_hd U1420 ( .A(n1089), .B(n1220), .C(n1088), .D(n1087), .Y(n405) );
  ao22d1_hd U1421 ( .A(n711), .B(sum[17]), .C(n709), .D(sum[16]), .Y(n1093) );
  ao21d1_hd U1422 ( .A(n657), .B(n1090), .C(n576), .Y(n1095) );
  ao22d1_hd U1423 ( .A(n569), .B(n1095), .C(n1094), .D(n568), .Y(n1091) );
  ao21d1_hd U1424 ( .A(n579), .B(z_m[12]), .C(n1091), .Y(n1092) );
  oa211d1_hd U1425 ( .A(n1229), .B(n674), .C(n1093), .D(n1092), .Y(n404) );
  ao22d1_hd U1426 ( .A(n711), .B(sum[18]), .C(n709), .D(sum[17]), .Y(n1099) );
  oa21d1_hd U1427 ( .A(z_m[14]), .B(n1094), .C(n669), .Y(n1097) );
  oa21d1_hd U1428 ( .A(n569), .B(n619), .C(n1095), .Y(n1096) );
  ao22d1_hd U1429 ( .A(z_m[13]), .B(n1097), .C(z_m[14]), .D(n1096), .Y(n1098)
         );
  oa211d1_hd U1430 ( .A(n1231), .B(n673), .C(n1099), .D(n1098), .Y(n403) );
  ao22d1_hd U1431 ( .A(n711), .B(sum[19]), .C(n709), .D(sum[18]), .Y(n1103) );
  oa21d1_hd U1432 ( .A(n1100), .B(n652), .C(n615), .Y(n1104) );
  oa22d1_hd U1433 ( .A(z_m[15]), .B(n1105), .C(n668), .D(n1229), .Y(n1101) );
  ao21d1_hd U1434 ( .A(z_m[15]), .B(n1104), .C(n1101), .Y(n1102) );
  oa211d1_hd U1435 ( .A(n1230), .B(n672), .C(n1103), .D(n1102), .Y(n402) );
  ao21d1_hd U1436 ( .A(n657), .B(n1231), .C(n1104), .Y(n1109) );
  ao22d1_hd U1437 ( .A(n711), .B(sum[20]), .C(n709), .D(sum[19]), .Y(n1108) );
  oa21d1_hd U1438 ( .A(z_m[16]), .B(n1105), .C(n669), .Y(n1106) );
  ao22d1_hd U1439 ( .A(n571), .B(n1144), .C(z_m[15]), .D(n1106), .Y(n1107) );
  oa211d1_hd U1440 ( .A(n1109), .B(n1230), .C(n1108), .D(n1107), .Y(n401) );
  ao22d1_hd U1441 ( .A(n711), .B(sum[21]), .C(n709), .D(sum[20]), .Y(n1115) );
  ao21d1_hd U1442 ( .A(n658), .B(n1111), .C(n575), .Y(n1117) );
  ao22d1_hd U1443 ( .A(n571), .B(n1117), .C(n1116), .D(n570), .Y(n1112) );
  ao21d1_hd U1444 ( .A(n580), .B(z_m[16]), .C(n1112), .Y(n1114) );
  oa211d1_hd U1445 ( .A(n1225), .B(n674), .C(n1115), .D(n1114), .Y(n400) );
  ao22d1_hd U1446 ( .A(n711), .B(sum[22]), .C(n708), .D(sum[21]), .Y(n1122) );
  oa21d1_hd U1447 ( .A(z_m[18]), .B(n1116), .C(n668), .Y(n1120) );
  oa21d1_hd U1448 ( .A(n571), .B(n620), .C(n1117), .Y(n1119) );
  ao22d1_hd U1449 ( .A(z_m[17]), .B(n1120), .C(z_m[18]), .D(n1119), .Y(n1121)
         );
  oa211d1_hd U1450 ( .A(n1227), .B(n673), .C(n1122), .D(n1121), .Y(n399) );
  ao22d1_hd U1451 ( .A(n714), .B(sum[23]), .C(n708), .D(sum[22]), .Y(n1126) );
  oa21d1_hd U1452 ( .A(n1123), .B(n652), .C(n1110), .Y(n1127) );
  oa22d1_hd U1453 ( .A(z_m[19]), .B(n1129), .C(n670), .D(n1225), .Y(n1124) );
  ao21d1_hd U1454 ( .A(z_m[19]), .B(n1127), .C(n1124), .Y(n1125) );
  oa211d1_hd U1455 ( .A(n1226), .B(n672), .C(n1126), .D(n1125), .Y(n398) );
  ao21d1_hd U1456 ( .A(n658), .B(n1227), .C(n1127), .Y(n1133) );
  ao22d1_hd U1457 ( .A(n1151), .B(sum[24]), .C(n708), .D(sum[23]), .Y(n1132)
         );
  oa21d1_hd U1458 ( .A(z_m[20]), .B(n1129), .C(n668), .Y(n1130) );
  ao22d1_hd U1459 ( .A(z_m[21]), .B(n1144), .C(z_m[19]), .D(n1130), .Y(n1131)
         );
  oa211d1_hd U1460 ( .A(n1133), .B(n1226), .C(n1132), .D(n1131), .Y(n397) );
  ao22d1_hd U1461 ( .A(n714), .B(sum[25]), .C(n708), .D(sum[24]), .Y(n1138) );
  ivd1_hd U1462 ( .A(z_m[21]), .Y(n1228) );
  oa22d1_hd U1463 ( .A(n1134), .B(n1228), .C(n668), .D(n1226), .Y(n1135) );
  ao21d1_hd U1464 ( .A(n1136), .B(n1228), .C(n1135), .Y(n1137) );
  oa211d1_hd U1465 ( .A(n564), .B(n674), .C(n1138), .D(n1137), .Y(n396) );
  ao22d1_hd U1466 ( .A(n714), .B(sum[26]), .C(n708), .D(sum[25]), .Y(n1143) );
  oa22d1_hd U1467 ( .A(z_m[22]), .B(n1139), .C(n1228), .D(n668), .Y(n1140) );
  ao21d1_hd U1468 ( .A(n565), .B(n1141), .C(n1140), .Y(n1142) );
  oa211d1_hd U1469 ( .A(n1145), .B(n673), .C(n1143), .D(n1142), .Y(n395) );
  ivd1_hd U1470 ( .A(round_bit), .Y(n1149) );
  ao22d1_hd U1471 ( .A(n714), .B(sum[2]), .C(n708), .D(sum[1]), .Y(n1148) );
  nd3d1_hd U1472 ( .A(n636), .B(guard), .C(n265), .Y(n1147) );
  oa211d1_hd U1473 ( .A(n1149), .B(n265), .C(n1148), .D(n1147), .Y(n394) );
  scg12d1_hd U1474 ( .A(round_bit), .B(n635), .C(n1150), .Y(n1154) );
  ao22d1_hd U1475 ( .A(n1152), .B(sum[0]), .C(n1151), .D(sum[1]), .Y(n1153) );
  scg4d1_hd U1476 ( .A(b_m[3]), .B(n664), .C(z_m[0]), .D(n632), .E(a_m[3]), 
        .F(n638), .G(n724), .H(z[0]), .Y(n392) );
  scg4d1_hd U1477 ( .A(b_m[4]), .B(n665), .C(z_m[1]), .D(n633), .E(a_m[4]), 
        .F(n639), .G(n727), .H(z[1]), .Y(n391) );
  scg4d1_hd U1478 ( .A(b_m[5]), .B(n666), .C(z_m[2]), .D(n634), .E(a_m[5]), 
        .F(n640), .G(n727), .H(z[2]), .Y(n390) );
  scg4d1_hd U1479 ( .A(b_m[6]), .B(n667), .C(z_m[3]), .D(n1163), .E(a_m[6]), 
        .F(n637), .G(n727), .H(z[3]), .Y(n389) );
  scg4d1_hd U1480 ( .A(n602), .B(n664), .C(z_m[4]), .D(n632), .E(a_m[7]), .F(
        n638), .G(n727), .H(z[4]), .Y(n388) );
  scg4d1_hd U1481 ( .A(b_m[8]), .B(n665), .C(n614), .D(n633), .E(a_m[8]), .F(
        n639), .G(n727), .H(z[5]), .Y(n387) );
  scg4d1_hd U1482 ( .A(b_m[9]), .B(n666), .C(z_m[6]), .D(n634), .E(n553), .F(
        n640), .G(n727), .H(z[6]), .Y(n386) );
  scg4d1_hd U1483 ( .A(b_m[10]), .B(n667), .C(z_m[7]), .D(n1163), .E(a_m[10]), 
        .F(n637), .G(n726), .H(z[7]), .Y(n385) );
  scg4d1_hd U1484 ( .A(n543), .B(n664), .C(z_m[8]), .D(n632), .E(n539), .F(
        n638), .G(n726), .H(z[8]), .Y(n384) );
  scg4d1_hd U1485 ( .A(n608), .B(n665), .C(n567), .D(n633), .E(a_m[12]), .F(
        n639), .G(n726), .H(z[9]), .Y(n383) );
  scg4d1_hd U1486 ( .A(b_m[13]), .B(n666), .C(z_m[10]), .D(n634), .E(n547), 
        .F(n640), .G(n726), .H(z[10]), .Y(n382) );
  scg4d1_hd U1487 ( .A(n551), .B(n667), .C(z_m[11]), .D(n1163), .E(a_m[14]), 
        .F(n637), .G(n726), .H(z[11]), .Y(n381) );
  scg4d1_hd U1488 ( .A(b_m[15]), .B(n664), .C(z_m[12]), .D(n632), .E(a_m[15]), 
        .F(n638), .G(n725), .H(z[12]), .Y(n380) );
  scg4d1_hd U1489 ( .A(b_m[16]), .B(n665), .C(n569), .D(n633), .E(a_m[16]), 
        .F(n639), .G(n725), .H(z[13]), .Y(n379) );
  scg4d1_hd U1490 ( .A(b_m[17]), .B(n666), .C(z_m[14]), .D(n634), .E(a_m[17]), 
        .F(n640), .G(n725), .H(z[14]), .Y(n378) );
  scg4d1_hd U1491 ( .A(b_m[18]), .B(n667), .C(z_m[15]), .D(n1163), .E(a_m[18]), 
        .F(n637), .G(n725), .H(z[15]), .Y(n377) );
  scg4d1_hd U1492 ( .A(b_m[19]), .B(n664), .C(z_m[16]), .D(n632), .E(a_m[19]), 
        .F(n638), .G(n725), .H(z[16]), .Y(n376) );
  scg4d1_hd U1493 ( .A(b_m[20]), .B(n665), .C(n571), .D(n633), .E(n604), .F(
        n639), .G(n725), .H(z[17]), .Y(n375) );
  scg4d1_hd U1494 ( .A(b_m[21]), .B(n666), .C(z_m[18]), .D(n634), .E(n555), 
        .F(n640), .G(n726), .H(z[18]), .Y(n374) );
  scg4d1_hd U1495 ( .A(b_m[22]), .B(n667), .C(z_m[19]), .D(n1163), .E(n541), 
        .F(n637), .G(n724), .H(z[19]), .Y(n373) );
  scg4d1_hd U1496 ( .A(b_m[23]), .B(n664), .C(z_m[20]), .D(n632), .E(a_m[23]), 
        .F(n638), .G(n724), .H(z[20]), .Y(n372) );
  scg4d1_hd U1497 ( .A(b_m[24]), .B(n665), .C(z_m[21]), .D(n633), .E(n561), 
        .F(n639), .G(n724), .H(z[21]), .Y(n371) );
  nr3d1_hd U1498 ( .A(n815), .B(n1210), .C(n1205), .Y(n1162) );
  ivd1_hd U1499 ( .A(n1159), .Y(n1161) );
  oa22d1_hd U1500 ( .A(n1161), .B(n1205), .C(n1160), .D(n1210), .Y(n1211) );
  nr2d1_hd U1501 ( .A(n1162), .B(n1211), .Y(n1169) );
  ao22d1_hd U1502 ( .A(a_m[25]), .B(n637), .C(z_m[22]), .D(n634), .Y(n1167) );
  ao22d1_hd U1503 ( .A(b_m[25]), .B(n666), .C(n723), .D(z[22]), .Y(n1166) );
  oa211d1_hd U1504 ( .A(n1169), .B(n1168), .C(n1167), .D(n1166), .Y(n370) );
  nr4d1_hd U1505 ( .A(n1171), .B(n1196), .C(n1170), .D(n1178), .Y(n1175) );
  nr4d1_hd U1506 ( .A(z_m[23]), .B(z_e[0]), .C(n1173), .D(n1172), .Y(n1174) );
  nr2bd1_hd U1507 ( .AN(z_e[0]), .B(n1178), .Y(n1179) );
  nr2d1_hd U1508 ( .A(z_e[1]), .B(z_e[0]), .Y(n1184) );
  nr2d1_hd U1509 ( .A(n1179), .B(n1184), .Y(n1180) );
  ivd1_hd U1510 ( .A(n1184), .Y(n1181) );
  ivd1_hd U1511 ( .A(z_e[2]), .Y(n1183) );
  ao22d1_hd U1512 ( .A(z_e[2]), .B(n1181), .C(n1184), .D(n1183), .Y(n1182) );
  nr2d1_hd U1513 ( .A(z_e[3]), .B(n1185), .Y(n1190) );
  ao21d1_hd U1514 ( .A(z_e[3]), .B(n1185), .C(n1190), .Y(n1186) );
  ivd1_hd U1515 ( .A(n1190), .Y(n1187) );
  ao22d1_hd U1516 ( .A(z_e[4]), .B(n1187), .C(n1190), .D(n1189), .Y(n1188) );
  nr2d1_hd U1517 ( .A(z_e[5]), .B(n1191), .Y(n1193) );
  ao21d1_hd U1518 ( .A(z_e[5]), .B(n1191), .C(n1193), .Y(n1192) );
  ivd1_hd U1519 ( .A(n1193), .Y(n1194) );
  nr2d1_hd U1520 ( .A(z_e[6]), .B(n1194), .Y(n1198) );
  ao21d1_hd U1521 ( .A(z_e[6]), .B(n1194), .C(n1198), .Y(n1195) );
  ivd1_hd U1522 ( .A(n1198), .Y(n1197) );
  ao22d1_hd U1523 ( .A(z_e[7]), .B(n1198), .C(n1197), .D(n1196), .Y(n1202) );
  oa211d1_hd U1524 ( .A(n1206), .B(n1205), .C(n1204), .D(n1203), .Y(n1213) );
  ao21d1_hd U1525 ( .A(n1210), .B(n1209), .C(n1208), .Y(n1212) );
  ao211d1_hd U1526 ( .A(a_s), .B(n1213), .C(n1212), .D(n1211), .Y(n1242) );
  nd4d1_hd U1527 ( .A(n1217), .B(n1216), .C(n1215), .D(n1214), .Y(n1218) );
  nr4d1_hd U1528 ( .A(z_m[22]), .B(n563), .C(z_m[5]), .D(n1218), .Y(n1237) );
  nd4d1_hd U1529 ( .A(n568), .B(n1220), .C(n566), .D(n1219), .Y(n1235) );
  nd4d1_hd U1530 ( .A(n1224), .B(n1223), .C(n1222), .D(n1221), .Y(n1234) );
  nd4d1_hd U1531 ( .A(n1228), .B(n1227), .C(n1226), .D(n1225), .Y(n1233) );
  nd4d1_hd U1532 ( .A(n570), .B(n1231), .C(n1230), .D(n1229), .Y(n1232) );
  nr4d1_hd U1533 ( .A(n1235), .B(n1234), .C(n1233), .D(n1232), .Y(n1236) );
  oa211d1_hd U1534 ( .A(n1239), .B(n1238), .C(n1244), .D(z_s), .Y(n1240) );
  oa211d1_hd U1535 ( .A(n1242), .B(n1250), .C(n1241), .D(n1240), .Y(n361) );
  nr2d1_hd U1536 ( .A(n721), .B(o_Z_STB), .Y(n136) );
  nr3d1_hd U1537 ( .A(n1245), .B(n93), .C(n1244), .Y(n111) );
  oa22d1_hd U1538 ( .A(n1248), .B(n1247), .C(DP_OP_154J1_137_6175_n25), .D(
        n1246), .Y(n128) );
  nr2d1_hd U1539 ( .A(n1263), .B(n1264), .Y(n1267) );
  nr2d1_hd U1540 ( .A(n1278), .B(n1277), .Y(n1282) );
  nr2d1_hd U1541 ( .A(n1294), .B(n1293), .Y(n1298) );
  ao21d1_hd U1542 ( .A(n1358), .B(n1316), .C(n533), .Y(n1315) );
  oa21d1_hd U1543 ( .A(b_e[7]), .B(n1299), .C(n1315), .Y(n1320) );
  ao21d1_hd U1544 ( .A(n577), .B(n1249), .C(n1320), .Y(n1252) );
  ivd1_hd U1545 ( .A(b[25]), .Y(n1268) );
  nr2d1_hd U1546 ( .A(n1269), .B(n1268), .Y(n1279) );
  ivd1_hd U1547 ( .A(b[27]), .Y(n1283) );
  nr2d1_hd U1548 ( .A(n1284), .B(n1283), .Y(n1295) );
  ivd1_hd U1549 ( .A(b[29]), .Y(n1302) );
  nr2d1_hd U1550 ( .A(n1303), .B(n1302), .Y(n1312) );
  nr2d1_hd U1551 ( .A(n1312), .B(n625), .Y(n1305) );
  oa211d1_hd U1552 ( .A(n1252), .B(n1251), .C(n535), .D(n1318), .Y(n504) );
  ao22d1_hd U1553 ( .A(n731), .B(b[22]), .C(b_m[26]), .D(n643), .Y(n1254) );
  oa21d1_hd U1554 ( .A(n1256), .B(n660), .C(n1254), .Y(n503) );
  scg12d1_hd U1555 ( .A(n1258), .B(n1257), .C(n1390), .Y(n112) );
  scg12d1_hd U1556 ( .A(n1260), .B(n1259), .C(n677), .Y(n106) );
  nr2d1_hd U1557 ( .A(b_e[0]), .B(n1299), .Y(n1262) );
  ao21d1_hd U1558 ( .A(n532), .B(b_e[0]), .C(n1262), .Y(n1261) );
  oa21d1_hd U1559 ( .A(b[23]), .B(n625), .C(n1261), .Y(n498) );
  nr2d1_hd U1560 ( .A(n533), .B(n1262), .Y(n1272) );
  oa22d1_hd U1561 ( .A(n1272), .B(n1264), .C(n1263), .D(n1271), .Y(n1266) );
  oa211d1_hd U1562 ( .A(b[24]), .B(b[23]), .C(n738), .D(n1269), .Y(n1265) );
  nd3bd1_hd U1563 ( .AN(n1266), .B(n534), .C(n1265), .Y(n497) );
  ao211d1_hd U1564 ( .A(n1269), .B(n1268), .C(n1279), .D(n625), .Y(n1274) );
  ivd1_hd U1565 ( .A(b_e[2]), .Y(n1270) );
  ao21d1_hd U1566 ( .A(n1272), .B(n1271), .C(n1270), .Y(n1273) );
  nr2d1_hd U1567 ( .A(n1274), .B(n1273), .Y(n1275) );
  oa211d1_hd U1568 ( .A(n649), .B(n1276), .C(n1275), .D(n534), .Y(n496) );
  ao21d1_hd U1569 ( .A(n671), .B(n1277), .C(n533), .Y(n1287) );
  oa22d1_hd U1570 ( .A(n1287), .B(n1278), .C(n1277), .D(n1286), .Y(n1281) );
  oa211d1_hd U1571 ( .A(n1279), .B(b[26]), .C(n738), .D(n1284), .Y(n1280) );
  nd3bd1_hd U1572 ( .AN(n1281), .B(n535), .C(n1280), .Y(n495) );
  ao211d1_hd U1573 ( .A(n1284), .B(n1283), .C(n1295), .D(n627), .Y(n1289) );
  ao21d1_hd U1574 ( .A(n1287), .B(n1286), .C(n1285), .Y(n1288) );
  nr2d1_hd U1575 ( .A(n1289), .B(n1288), .Y(n1290) );
  oa211d1_hd U1576 ( .A(b_e[4]), .B(n1291), .C(n1290), .D(n534), .Y(n494) );
  ao21d1_hd U1577 ( .A(n671), .B(n1293), .C(n532), .Y(n1301) );
  oa22d1_hd U1578 ( .A(n1301), .B(n1294), .C(n1293), .D(n1300), .Y(n1297) );
  oa211d1_hd U1579 ( .A(n1295), .B(b[28]), .C(n738), .D(n1303), .Y(n1296) );
  nd3bd1_hd U1580 ( .AN(n1297), .B(n534), .C(n1296), .Y(n493) );
  ao22d1_hd U1581 ( .A(n648), .B(n1306), .C(n1305), .D(n1304), .Y(n1308) );
  oa211d1_hd U1582 ( .A(n648), .B(n1309), .C(n1308), .D(n535), .Y(n492) );
  nr2d1_hd U1583 ( .A(n626), .B(n1310), .Y(n1313) );
  nr2d1_hd U1584 ( .A(n1299), .B(n1316), .Y(n1311) );
  ao22d1_hd U1585 ( .A(n1313), .B(n1312), .C(n1311), .D(n1317), .Y(n1314) );
  oa211d1_hd U1586 ( .A(n1315), .B(n1317), .C(n1314), .D(n1318), .Y(n491) );
  nr4d1_hd U1587 ( .A(b_e[8]), .B(n1317), .C(n1299), .D(n1316), .Y(n1319) );
  ao21d1_hd U1588 ( .A(n647), .B(n1322), .C(n1321), .Y(n1325) );
  oa211d1_hd U1589 ( .A(n1325), .B(n1324), .C(n1383), .D(n645), .Y(n489) );
  nr2d1_hd U1590 ( .A(a_e[0]), .B(n1379), .Y(n1327) );
  ao21d1_hd U1591 ( .A(n1357), .B(a_e[0]), .C(n1327), .Y(n1326) );
  oa21d1_hd U1592 ( .A(a[23]), .B(n626), .C(n1326), .Y(n488) );
  nr2d1_hd U1593 ( .A(n1357), .B(n1327), .Y(n1337) );
  oa22d1_hd U1594 ( .A(n1337), .B(n1329), .C(n1328), .D(n1336), .Y(n1331) );
  oa211d1_hd U1595 ( .A(a[24]), .B(a[23]), .C(n738), .D(n1334), .Y(n1330) );
  nd3bd1_hd U1596 ( .AN(n1331), .B(n645), .C(n1330), .Y(n487) );
  ao211d1_hd U1597 ( .A(n1334), .B(n1333), .C(n1344), .D(n625), .Y(n1339) );
  ao21d1_hd U1598 ( .A(n1337), .B(n1336), .C(n1335), .Y(n1338) );
  nr2d1_hd U1599 ( .A(n1339), .B(n1338), .Y(n1340) );
  oa211d1_hd U1600 ( .A(a_e[2]), .B(n1341), .C(n1340), .D(n1373), .Y(n486) );
  ao21d1_hd U1601 ( .A(n671), .B(n1342), .C(n1357), .Y(n1352) );
  oa22d1_hd U1602 ( .A(n1352), .B(n1343), .C(n1342), .D(n1351), .Y(n1346) );
  oa211d1_hd U1603 ( .A(n1344), .B(a[26]), .C(n738), .D(n1349), .Y(n1345) );
  nd3bd1_hd U1604 ( .AN(n1346), .B(n645), .C(n1345), .Y(n485) );
  ao211d1_hd U1605 ( .A(n1349), .B(n1348), .C(n1361), .D(n626), .Y(n1354) );
  ao21d1_hd U1606 ( .A(n1352), .B(n1351), .C(n1350), .Y(n1353) );
  nr2d1_hd U1607 ( .A(n1354), .B(n1353), .Y(n1355) );
  oa211d1_hd U1608 ( .A(a_e[4]), .B(n1356), .C(n1355), .D(n1373), .Y(n484) );
  ao21d1_hd U1609 ( .A(n671), .B(n1359), .C(n1357), .Y(n1369) );
  oa22d1_hd U1610 ( .A(n1369), .B(n1360), .C(n1359), .D(n1368), .Y(n1363) );
  oa211d1_hd U1611 ( .A(n1361), .B(a[28]), .C(n738), .D(n1367), .Y(n1362) );
  nd3bd1_hd U1612 ( .AN(n1363), .B(n645), .C(n1362), .Y(n483) );
  ao22d1_hd U1613 ( .A(n1372), .B(n1371), .C(a_e[6]), .D(n1370), .Y(n1374) );
  oa211d1_hd U1614 ( .A(a_e[6]), .B(n1375), .C(n1374), .D(n1373), .Y(n482) );
  nr2d1_hd U1615 ( .A(n1377), .B(n627), .Y(n1381) );
  nr2d1_hd U1616 ( .A(n1379), .B(n1378), .Y(n1380) );
  ao22d1_hd U1617 ( .A(n1382), .B(n1381), .C(n1380), .D(n1385), .Y(n1384) );
  oa211d1_hd U1618 ( .A(n1386), .B(n646), .C(n1384), .D(n1383), .Y(n481) );
  oa21d1_hd U1619 ( .A(n1388), .B(n1387), .C(n572), .Y(n2) );
  scg6d1_hd U1620 ( .A(n1391), .B(n1390), .C(n654), .Y(n1) );
endmodule

