module pad_FIR_FILTER(   //top module
	input RESET,CLK,WR,
	input [15:0] iDATA,
	output [38:0] oDATA);

// wires from the package to the pins of the pads
//wire RESET, CLK, WR;
//wire [15:0] iDATA;
//wire [38:0] oDATA;
//wires from the pins of the pads to the core
wire RESET_c, CLK_c, WR_c;
wire [15:0] iDATA_c;
wire [38:0] oDATA_c;
// the core is instantiated with the name "core_FIR_FILTER"
FIR_FILTER core_FIR_FILTER(RESET_c,CLK_c, WR_c, iDATA_c, oDATA_c);

// Top pad (52) 
// input pads, based upon the module phic (PAD,PI,PO,Y)
  phic pad0( .PAD(RESET), .PI(1'b0), .PO(), .Y(RESET_c) );
  phic pad1( .PAD(CLK), .PI(1'b0), .PO(), .Y(CLK_c) );
  phic pad2( .PAD(WR), .PI(1'b0), .PO(), .Y(WR_c) );
  phic pad3( .PAD(iDATA[0]), .PI(1'b0), .PO(), .Y(iDATA_c[0]) );
  phic pad4( .PAD(iDATA[1]), .PI(1'b0), .PO(), .Y(iDATA_c[1]) );
  phic pad5( .PAD(iDATA[2]), .PI(1'b0), .PO(), .Y(iDATA_c[2]) );
  phic pad6( .PAD(iDATA[3]), .PI(1'b0), .PO(), .Y(iDATA_c[3]) );
  phic pad7( .PAD(iDATA[4]), .PI(1'b0), .PO(), .Y(iDATA_c[4]) );
  phic pad8( .PAD(iDATA[5]), .PI(1'b0), .PO(), .Y(iDATA_c[5]) );
  phic pad9( .PAD(iDATA[6]), .PI(1'b0), .PO(), .Y(iDATA_c[6]) );
  phic pad10( .PAD(iDATA[7]), .PI(1'b0), .PO(), .Y(iDATA_c[7]) );
  phic pad11( .PAD(iDATA[8]), .PI(1'b0), .PO(), .Y(iDATA_c[8]) );
  phic pad12( .PAD(iDATA[9]), .PI(1'b0), .PO(), .Y(iDATA_c[9]) );
  phic pad13( .PAD(iDATA[10]), .PI(1'b0), .PO(), .Y(iDATA_c[10]) );
  phic pad14( .PAD(iDATA[11]), .PI(1'b0), .PO(), .Y(iDATA_c[11]) );
  phic pad15( .PAD(iDATA[12]), .PI(1'b0), .PO(), .Y(iDATA_c[12]) );
  phic pad16( .PAD(iDATA[13]), .PI(1'b0), .PO(), .Y(iDATA_c[13]) );
  phic pad17( .PAD(iDATA[14]), .PI(1'b0), .PO(), .Y(iDATA_c[14]) );
  phic pad18( .PAD(iDATA[15]), .PI(1'b0), .PO(), .Y(iDATA_c[15]) ); 
  phic pad19();
  phic pad20();
  phic pad21();
  phic pad22();
  phic pad23();
  phic pad24();
  phic pad25();
  phic pad26();
  phic pad27();
  phic pad28();
  phic pad29();
  phic pad30();
  phic pad31();
  phic pad32();

  vssoh pad33();
  vssoh pad34();
  vssoh pad35();
  vssoh pad36();
  vssoh pad37();
  vssoh pad38();
  vssoh pad39();
// output pads, based upon the module phob12 (A,PAD)
phob12 pad40(.A(oDATA_c[0]), .PAD(oDATA[0])); 
phob12 pad41(.A(oDATA_c[1]), .PAD(oDATA[1])); 
phob12 pad42(.A(oDATA_c[2]), .PAD(oDATA[2])); 
phob12 pad43(.A(oDATA_c[3]), .PAD(oDATA[3])); 
phob12 pad44(.A(oDATA_c[4]), .PAD(oDATA[4])); 
phob12 pad45(.A(oDATA_c[5]), .PAD(oDATA[5])); 
phob12 pad46(.A(oDATA_c[6]), .PAD(oDATA[6])); 
phob12 pad47(.A(oDATA_c[7]), .PAD(oDATA[7])); 
phob12 pad48(.A(oDATA_c[8]), .PAD(oDATA[8])); 
phob12 pad49(.A(oDATA_c[9]), .PAD(oDATA[9])); 
phob12 pad50(.A(oDATA_c[10]), .PAD(oDATA[10])); 
// Right pad(52)
phob12 pad51(.A(oDATA_c[11]), .PAD(oDATA[11])); 
phob12 pad52(.A(oDATA_c[12]), .PAD(oDATA[12])); 
phob12 pad53(.A(oDATA_c[13]), .PAD(oDATA[13])); 
phob12 pad54(.A(oDATA_c[14]), .PAD(oDATA[14])); 
phob12 pad55(.A(oDATA_c[15]), .PAD(oDATA[15])); 
phob12 pad56(.A(oDATA_c[16]), .PAD(oDATA[16])); 
phob12 pad57(.A(oDATA_c[17]), .PAD(oDATA[17])); 
phob12 pad58(.A(oDATA_c[18]), .PAD(oDATA[18])); 
phob12 pad59(.A(oDATA_c[19]), .PAD(oDATA[19])); 
phob12 pad60(.A(oDATA_c[20]), .PAD(oDATA[20])); 
phob12 pad61(.A(oDATA_c[21]), .PAD(oDATA[21])); 
phob12 pad62(.A(oDATA_c[22]), .PAD(oDATA[22])); 
phob12 pad63(.A(oDATA_c[23]), .PAD(oDATA[23])); 
phob12 pad64(.A(oDATA_c[24]), .PAD(oDATA[24])); 
phob12 pad65(.A(oDATA_c[25]), .PAD(oDATA[25])); 
phob12 pad66(.A(oDATA_c[26]), .PAD(oDATA[26])); 
phob12 pad67(.A(oDATA_c[27]), .PAD(oDATA[27])); 
phob12 pad68(.A(oDATA_c[28]), .PAD(oDATA[28])); 
phob12 pad69(.A(oDATA_c[29]), .PAD(oDATA[29])); 
phob12 pad70(.A(oDATA_c[30]), .PAD(oDATA[30])); 
phob12 pad71(.A(oDATA_c[31]), .PAD(oDATA[31])); 
phob12 pad72(.A(oDATA_c[32]), .PAD(oDATA[32])); 
phob12 pad73(.A(oDATA_c[33]), .PAD(oDATA[33])); 
phob12 pad74(.A(oDATA_c[34]), .PAD(oDATA[34])); 
phob12 pad75(.A(oDATA_c[35]), .PAD(oDATA[35])); 
phob12 pad76(.A(oDATA_c[36]), .PAD(oDATA[36])); 
phob12 pad77(.A(oDATA_c[37]), .PAD(oDATA[37])); 
phob12 pad78(.A(oDATA_c[38]), .PAD(oDATA[38])); 
phob12 pad79(); 
phob12 pad80(); 
phob12 pad81(); 
phob12 pad82(); 
phob12 pad83(); 
  vssoh pad84();
  vssoh pad85();
  vssoh pad86();
  vssoh pad87();
  vssoh pad88();
  vssoh pad89();
  vssoh pad90();
  vssoh pad91();
  vssoh pad92();
  vssoh pad93();
  vdd12ih pad94();
  vdd12ih pad95();
  vdd12ih pad96();
  vdd12ih pad97();
  vdd12ih pad98();
  vdd12ih pad99();
  vdd12ih pad100();
  vdd12ih pad101();
  vdd12ih pad102();
  vdd12ih pad103();

// Left pad -(52)
  phob12 pad104();
  phob12 pad105();
  phob12 pad106();
  phob12 pad109();
  phob12 pad110();
  phob12 pad111();
  phob12 pad112();
  phob12 pad113();
  phob12 pad114();
  phob12 pad115();
  phob12 pad116();
  phob12 pad117();
  phob12 pad118();
  phob12 pad119();
  phob12 pad120();
  phob12 pad121();
  phob12 pad122();
  phob12 pad123();
  phob12 pad124();
  phob12 pad125();
  phob12 pad126();
  phob12 pad127();
  phob12 pad128();
  phob12 pad129();
  phob12 pad130();
  phob12 pad132();
  phob12 pad133();
  phob12 pad134();
  phob12 pad135();
  vssoh pad136();
  vssoh pad137();
  vssoh pad138();
  vssoh pad139();
  vssoh pad140();
  vssoh pad141();
  vssoh pad142();
  vssoh pad143();
  vssoh pad144();
  vssoh pad145();
  vdd12ih pad146();
  vdd12ih pad147();
  vdd12ih pad148();
  vdd12ih pad149();
  vdd12ih pad150();
  vdd12ih pad151();
  vdd12ih pad152();
  vdd12ih pad153();
  vdd12ih pad154();
  vdd12ih pad155();



// Bottom pad (52) 
  vdd33oph pad156();
  vdd33oph pad157();
  vdd33oph pad158();
  vdd33oph pad159();
  vdd33oph pad160();
  vdd33oph pad161();
  vdd33oph pad162();
  vdd33oph pad163();
  vdd33oph pad164();
  vdd33oph pad165();
  phic pad166();
  phic pad167();
  vdd12ih pad168();
  vdd12ih pad169();
  vdd12ih pad170();
  vdd12ih pad171();
  vdd12ih pad172();
  vdd12ih pad173();
  vdd12ih pad174();
  vdd12ih pad175();
  vdd12ih pad176();
  vdd12ih pad177();
  vdd12ih pad178();
  vdd12ih pad179();
  vdd12ih pad180();
  vdd12ih pad181();
  vdd12ih pad182();
  vdd12ih pad183();
  vdd12ih pad184();
  vdd12ih pad185();
  vdd12ih pad186();
  vdd12ih pad187();
  vssoh pad188();
  vssoh pad189();
  vssoh pad190();
  vssoh pad191();
  vssoh pad192();
  vssoh pad193();
  vssoh pad194();
  vssoh pad195();
  vssoh pad196();
  vssoh pad197();
  vssoh pad198();
  vssoh pad199();
  vssoh pad200();
  vssoh pad201();
  vssoh pad202();
  vssoh pad203();
  vssoh pad204();
  vssoh pad205();
  vssoh pad206();
  vssoh pad207();

endmodule
