
module FIR_FILTER_PAD ( RESET, CLK, WR, IDATA, ODATA );
  input [15:0] IDATA;
  output [38:0] ODATA;
  input RESET, CLK, WR;
  wire   w_reset, w_clk, w_wr;
  wire   [15:0] w_idata;
  wire   [38:0] w_odata;

  FIR_FILTER FIR1 ( .RESET(w_reset), .CLK(w_clk), .WR(w_wr), .iDATA(w_idata), .oDATA(
        w_odata) );
  phic pad1 ( .PAD(IDATA[0]), .PI(1'b0), .PO(),  .Y(w_idata[0]) );
  phic pad2 ( .PAD(IDATA[1]), .PI(1'b0), .PO(),  .Y(w_idata[1]) );
  phic pad3 ( .PAD(IDATA[2]), .PI(1'b0), .PO(),  .Y(w_idata[2]) );
  phic pad4 ( .PAD(IDATA[3]), .PI(1'b0), .PO(),  .Y(w_idata[3]) );
  phic pad5 ( .PAD(IDATA[4]), .PI(1'b0), .PO(),  .Y(w_idata[4]) );
  phic pad6 ( .PAD(IDATA[5]), .PI(1'b0), .PO(),  .Y(w_idata[5]) );
  phic pad7 ( .PAD(IDATA[6]), .PI(1'b0), .PO(),  .Y(w_idata[6]) );
  phic pad8 ( .PAD(IDATA[7]), .PI(1'b0), .PO(),  .Y(w_idata[7]) );
  vdd33oph pad9 (  );
  vdd33oph pad10 (  );
  vdd33oph pad11 (  );
  vdd33oph pad12 (  );
  vdd33oph pad13 (  );
  vdd33oph pad14 (  );
  vdd33oph pad15 (  );
  vdd33oph pad16 (  );
  vssoh pad17 (  );
  vssoh pad18 (  );
  vssoh pad19 (  );
  vssoh pad20 (  );
  vssoh pad21 (  );
  vssoh pad22 (  );
  phic pad23 ( .PAD(IDATA[8]), .PI(1'b0), .PO(),  .Y(w_idata[8]) );
  phic pad24 ( .PAD(IDATA[9]), .PI(1'b0), .PO(),  .Y(w_idata[9]) );
  phic pad25 ( .PAD(IDATA[10]), .PI(1'b0), .PO(),  .Y(w_idata[10]) );
  phic pad26 ( .PAD(IDATA[11]), .PI(1'b0), .PO(),  .Y(w_idata[11]) );
  phic pad27 ( .PAD(IDATA[12]), .PI(1'b0), .PO(),  .Y(w_idata[12]) );
  phic pad28 ( .PAD(IDATA[13]), .PI(1'b0), .PO(),  .Y(w_idata[13]) );
  phic pad29 ( .PAD(IDATA[14]), .PI(1'b0), .PO(),  .Y(w_idata[14]) );
  phic pad30 ( .PAD(IDATA[15]), .PI(1'b0), .PO(),  .Y(w_idata[15]) );
  phob12 pad31 (  );
  phob12 pad32 (  );
  phob12 pad33 (  );
  phob12 pad34 (  );
  phob12 pad35 (  );
  phob12 pad36 (  );
  phob12 pad37 ( );
  phob12 pad38 ( .A(w_odata[16]), .PAD(ODATA[16]) );
  vdd33oph pad39 (  );
  vdd33oph pad40 (  );
  vdd33oph pad41 (  );
  vdd33oph pad42 (  );
  vdd33oph pad43 (  );
  vdd33oph pad44 (  );
  vdd33oph pad45 (  );
  vdd33oph pad46 (  );
  vssoh pad47 (  );
  vssoh pad48 (  );
  vssoh pad49 (  );
  vssoh pad50 (  );
  vssoh pad51 (  );
  vssoh pad52 (  );
  phob12 pad53 ( .A(w_odata[0]), .PAD(ODATA[0]) );
  phob12 pad54 ( .A(w_odata[1]), .PAD(ODATA[1]) );
  phob12 pad55 ( .A(w_odata[2]), .PAD(ODATA[2]) );
  phob12 pad56 ( .A(w_odata[3]), .PAD(ODATA[3]) );
  phob12 pad57 ( .A(w_odata[4]), .PAD(ODATA[4]) );
  phob12 pad58 ( .A(w_odata[5]), .PAD(ODATA[5]) );
  phob12 pad59 ( .A(w_odata[6]), .PAD(ODATA[6]) );
  phob12 pad60 ( .A(w_odata[7]), .PAD(ODATA[7]) );
  phob12 pad61 ( .A(w_odata[8]), .PAD(ODATA[8]) );
  phob12 pad62 ( .A(w_odata[9]), .PAD(ODATA[9]) );
  phob12 pad63 ( .A(w_odata[10]), .PAD(ODATA[10]) );
  phob12 pad64 ( .A(w_odata[11]), .PAD(ODATA[11]) );
  phob12 pad65 ( .A(w_odata[12]), .PAD(ODATA[12]) );
  phob12 pad66 ( .A(w_odata[13]), .PAD(ODATA[13]) );
  phob12 pad67 ( .A(w_odata[14]), .PAD(ODATA[14]) );
  phob12 pad68 ( .A(w_odata[15]), .PAD(ODATA[15]) );
  vdd33oph pad69 (  );
  vdd33oph pad70 (  );
  vdd33oph pad71 (  );
  vdd33oph pad72 (  );
  vdd33oph pad73 (  );
  vdd33oph pad74 (  );
  vdd33oph pad75 (  );
  vdd33oph pad76 (  );
  vssoh pad77 (  );
  vssoh pad78 (  );
  vssoh pad79 (  );
  vssoh pad80 (  );
  vssoh pad81 (  );
  vssoh pad82 (  );
  phob12 pad83 ( .A(w_odata[17]), .PAD(ODATA[17]) );
  phob12 pad84 ( .A(w_odata[18]), .PAD(ODATA[18]) );
  phob12 pad85 ( .A(w_odata[19]), .PAD(ODATA[19]) );
  phob12 pad86 ( .A(w_odata[20]), .PAD(ODATA[20]) );
  phob12 pad87 ( .A(w_odata[21]), .PAD(ODATA[21]) );
  phob12 pad88 ( .A(w_odata[22]), .PAD(ODATA[22]) );
  phob12 pad89 ( .A(w_odata[23]), .PAD(ODATA[23]) );
  phob12 pad90 ( .A(w_odata[24]), .PAD(ODATA[24]) );
  phob12 pad91 ( .A(w_odata[25]), .PAD(ODATA[25]) );
  phob12 pad92 ( .A(w_odata[26]), .PAD(ODATA[26]) );
  phob12 pad93 ( .A(w_odata[27]), .PAD(ODATA[27]) );
  phob12 pad94 ( .A(w_odata[28]), .PAD(ODATA[28]) );
  phob12 pad95 ( .A(w_odata[29]), .PAD(ODATA[29]) );
  phob12 pad96 ( .A(w_odata[30]), .PAD(ODATA[30]) );
  phob12 pad97 ( .A(w_odata[31]), .PAD(ODATA[31]) );
  phob12 pad98 ( .A(w_odata[32]), .PAD(ODATA[32]) );
  vdd33oph pad99 (  );
  vdd33oph pad100 (  );
  vdd33oph pad101 (  );
  vdd33oph pad102 (  );
  vdd33oph pad103 (  );
  vdd33oph pad104 (  );
  vdd33oph pad105 (  );
  vdd33oph pad106 (  );
  vssoh pad107 (  );
  vssoh pad108 (  );
  vssoh pad109 (  );
  vssoh pad110 (  );
  vssoh pad111 (  );
  phob12 pad112 ( .A(w_odata[33]), .PAD(ODATA[33]) );
  phob12 pad113 ( .A(w_odata[34]), .PAD(ODATA[34]) );
  phob12 pad114 ( .A(w_odata[35]), .PAD(ODATA[35]) );
  phob12 pad115 ( .A(w_odata[36]), .PAD(ODATA[36]) );
  phob12 pad116 ( .A(w_odata[37]), .PAD(ODATA[37]) );
  phob12 pad117 ( .A(w_odata[38]), .PAD(ODATA[38]) );
  phic pad118 ( .PAD(CLK), .PI(1'b0), .PO(),  .Y(w_clk) );
  phic pad119 ( .PAD(RESET), .PI(1'b0), .PO(),  .Y(w_reset) );
  phic pad120 ( .PAD(WR), .PI(1'b0), .PO(),  .Y(w_wr) );
  
  vdd12ih pad121 (  );
  vdd12ih pad122 (  );
  vdd12ih pad123 (  );
  vdd12ih pad124 (  );
  vdd12ih pad125 (  );
  vdd12ih pad126 (  );
  vssiph pad127 (  );
  vssiph pad128 (  );
  vssiph pad129 (  );
  vssiph pad130 (  );
  vssiph pad131 (  );
  vssiph pad132 (  );
  vssiph pad133 (  );
  vssiph pad134 (  );
  vssiph pad135 (  );
  vssiph pad136 (  );
  vssiph pad137 (  );
  vssiph pad138 (  );
  vssiph pad139 (  );
  vssiph pad140 (  );
  vssiph pad141 (  );
  vssiph pad142 (  );
  vssiph pad143 (  );
  vssiph pad144 (  );
  vssiph pad145 (  );
  vssiph pad146 (  );
  vssiph pad147 (  );
  vssiph pad148 (  );
  vssiph pad149 (  );
  vssiph pad150 (  );
  vssiph pad151 (  );
  vssoh pad152 (  );
  vssoh pad153 (  );
  vssoh pad154 (  );
  vssoh pad155 (  );
  vdd12ih pad156 (  );
  vdd12ih pad157 (  );
  vdd12ih pad158 (  );
  vdd12ih pad159 (  );
  vdd12ih pad160 (  );
  vdd12ih pad161 (  );
  vdd12ih pad162 (  );
  vdd12ih pad163 (  );
  vdd12ih pad164 (  );
  vdd12ih pad165 (  );
  vdd12ih pad166 (  );
  vdd12ih pad167 (  );
  vdd12ih pad168 (  );
  vdd12ih pad169 (  );
  vdd12ih pad170 (  );
  vdd12ih pad171 (  );
  vdd12ih pad172 (  );
  vdd12ih pad173 (  );
  vdd12ih pad174 (  );
  vdd12ih pad175 (  );
  vdd12ih pad176 (  );
  vdd12ih pad177 (  );
  vdd12ih pad178 (  );
  vdd12ih pad179 (  );
  vdd12ih pad180 (  );
  vdd12ih pad181 (  );
  vdd12ih pad182 (  );
  vdd12ih pad183 (  );
  vssoh pad184 (  );
  vssoh pad185 (  );
  vssoh pad186 (  );
  vssoh pad187 (  );
  vssoh pad188 (  );
  vssoh pad189 (  );
  vssoh pad190 (  );
  vssoh pad191 (  );
  vssiph pad192 (  );
  vssiph pad193 (  );
  vssiph pad194 (  );
  vssiph pad195 (  );
  vssiph pad196 (  );
  vssiph pad197 (  );
  vssiph pad198 (  );
  vssiph pad199 (  );
  vssiph pad200 (  );
  vssiph pad201 (  );
  vssiph pad202 (  );
  vssoh pad203 (  );
  vssoh pad204 (  );
  vssoh pad205 (  );
  vssoh pad206 (  );
  vssoh pad207 (  );
  vssoh pad208 (  );
  //vssoh pad209 (  );
  //vssoh pad210 (  );
  //vssoh pad211 (  );
  //vssoh pad212 (  );
  //vssoh pad213 (  );
  //vssoh pad214 (  );
  //vssoh pad215 (  );
  //vssoh pad216 (  );
  //vssoh pad217 (  );
  //vssoh pad218 (  );
  //vssoh pad219 (  );
  //vssoh pad220 (  );
  //vssoh pad221 (  );
  //vssoh pad222 (  );
  //vssoh pad223 (  );
  //vssoh pad224 (  );
  //vssoh pad225 (  );
  //vssoh pad226 (  );
  //vssoh pad227 (  );
  //vssoh pad228 (  );
  //vssoh pad229 (  );
  //vssoh pad230 (  );
  //vssoh pad231 (  );
  //vssoh pad232 (  );
  //vssoh pad233 (  );
  //vssoh pad234 (  );
  //vssoh pad235 (  );
  //vssoh pad236 (  );
  //vssoh pad237 (  );
  //vssoh pad238 (  );
  //vssoh pad239 (  );
  //vssoh pad240 (  );
  //vssoh pad241 (  );
  //vssoh pad242 (  );
  //vssoh pad243 (  );
  //vssoh pad244 (  );
  //vssoh pad245 (  );
  //vssoh pad246 (  );
  //vssoh pad247 (  );
  //vssoh pad248 (  );
  //vssoh pad249 (  );
  //vssoh pad250 (  );
  //vssoh pad251 (  );
  //vssoh pad252 (  );
  //vssoh pad253 (  );
  //vssoh pad254 (  );
  //vssoh pad255 (  );
  //vssoh pad256 (  );
  //vssoh pad257 (  );
  //vssoh pad258 (  );
  //vssoh pad259 (  );
  //vssoh pad260 (  );
  //vssoh pad261 (  );
  //vssoh pad262 (  );
  //vssoh pad263 (  );
  //vssoh pad264 (  );
  //vssoh pad265 (  );
  //vssoh pad266 (  );
  //vssoh pad267 (  );
  //vssoh pad268 (  );
  //vssoh pad269 (  );
  //vssoh pad270 (  );
  //vssoh pad271 (  );
  //vssoh pad272 (  );
  //vssoh pad273 (  );
  //vssoh pad274 (  );
  //vssoh pad275 (  );
  //vssoh pad276 (  );
  //vssoh pad277 (  );
  //vssoh pad278 (  );
  //vssoh pad279 (  );
  //vssoh pad280 (  );
endmodule

