
module float_adder ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n105,
         n109, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n125, n126, n131, n133, n134, n135, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n719, n720, n722,
         n723, n724, n725, n726, n727, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1660;
  wire   [1557:1554] n;

  scg21d1_hd U117 ( .A(o_AB_ACK), .B(n1271), .C(n206), .D(i_RST), .Y(n1117) );
  oa22d1_hd U119 ( .A(n1270), .B(n1269), .C(n1274), .D(n1268), .Y(n1116) );
  oa21d1_hd U121 ( .A(n49), .B(n1268), .C(n1267), .Y(n1115) );
  scg6d1_hd U122 ( .A(n1266), .B(n1028), .C(n1269), .Y(n1267) );
  oa22d1_hd U123 ( .A(n1265), .B(n1269), .C(n67), .D(n1268), .Y(n1114) );
  oa21d1_hd U134 ( .A(n1275), .B(n1268), .C(n1264), .Y(n1111) );
  scg6d1_hd U135 ( .A(n196), .B(n1013), .C(n1269), .Y(n1264) );
  nd4d1_hd U137 ( .A(n1266), .B(n1263), .C(n1272), .D(n896), .Y(n1268) );
  nr4d1_hd U138 ( .A(n204), .B(n1262), .C(n1261), .D(n1260), .Y(n1263) );
  scg16d1_hd U139 ( .A(n20), .B(n1286), .C(n1660), .Y(n1260) );
  ao211d1_hd U143 ( .A(n201), .B(n1259), .C(i_RST), .D(n1258), .Y(n1110) );
  ivd1_hd U485 ( .A(i_RST), .Y(n1660) );
  fad1_hd DP_OP_154J1_137_6175_U10 ( .A(n121), .B(n1377), .CI(n1376), .CO(
        n1027), .S(n1285) );
  fad1_hd DP_OP_154J1_137_6175_U9 ( .A(n122), .B(n1378), .CI(n1027), .CO(n1026), .S(n1284) );
  fad1_hd DP_OP_154J1_137_6175_U8 ( .A(n120), .B(n1379), .CI(n1026), .CO(n1025), .S(n1283) );
  fad1_hd DP_OP_154J1_137_6175_U7 ( .A(n121), .B(n1380), .CI(n1025), .CO(n1024), .S(n1282) );
  fad1_hd DP_OP_154J1_137_6175_U6 ( .A(n122), .B(n1381), .CI(n1024), .CO(n1023), .S(n1281) );
  fad1_hd DP_OP_154J1_137_6175_U5 ( .A(n120), .B(n1382), .CI(n1023), .CO(n1022), .S(n1280) );
  fad1_hd DP_OP_154J1_137_6175_U4 ( .A(n120), .B(n1383), .CI(n1022), .CO(n1021), .S(n1279) );
  fad1_hd DP_OP_154J1_137_6175_U3 ( .A(n121), .B(n1384), .CI(n1021), .CO(n1020), .S(n1278) );
  fd1qd1_hd z_e_reg_0_ ( .D(n1189), .CK(i_CLK), .Q(n1376) );
  fd1qd1_hd a_e_reg_3_ ( .D(n1131), .CK(i_CLK), .Q(n1483) );
  fd1qd1_hd b_e_reg_0_ ( .D(n1118), .CK(i_CLK), .Q(n1443) );
  fd1qd1_hd b_e_reg_3_ ( .D(n1121), .CK(i_CLK), .Q(n1446) );
  fd1qd1_hd z_reg_31_ ( .D(n1255), .CK(i_CLK), .Q(n1347) );
  fd1qd1_hd z_reg_0_ ( .D(n1224), .CK(i_CLK), .Q(n1316) );
  fd1qd1_hd z_reg_1_ ( .D(n1225), .CK(i_CLK), .Q(n1317) );
  fd1qd1_hd z_reg_2_ ( .D(n1226), .CK(i_CLK), .Q(n1318) );
  fd1qd1_hd z_reg_3_ ( .D(n1227), .CK(i_CLK), .Q(n1319) );
  fd1qd1_hd z_reg_4_ ( .D(n1228), .CK(i_CLK), .Q(n1320) );
  fd1qd1_hd z_reg_5_ ( .D(n1229), .CK(i_CLK), .Q(n1321) );
  fd1qd1_hd z_reg_6_ ( .D(n1230), .CK(i_CLK), .Q(n1322) );
  fd1qd1_hd z_reg_7_ ( .D(n1231), .CK(i_CLK), .Q(n1323) );
  fd1qd1_hd z_reg_8_ ( .D(n1232), .CK(i_CLK), .Q(n1324) );
  fd1qd1_hd z_reg_9_ ( .D(n1233), .CK(i_CLK), .Q(n1325) );
  fd1qd1_hd z_reg_10_ ( .D(n1234), .CK(i_CLK), .Q(n1326) );
  fd1qd1_hd z_reg_11_ ( .D(n1235), .CK(i_CLK), .Q(n1327) );
  fd1qd1_hd z_reg_12_ ( .D(n1236), .CK(i_CLK), .Q(n1328) );
  fd1qd1_hd z_reg_13_ ( .D(n1237), .CK(i_CLK), .Q(n1329) );
  fd1qd1_hd z_reg_14_ ( .D(n1238), .CK(i_CLK), .Q(n1330) );
  fd1qd1_hd z_reg_15_ ( .D(n1239), .CK(i_CLK), .Q(n1331) );
  fd1qd1_hd z_reg_16_ ( .D(n1240), .CK(i_CLK), .Q(n1332) );
  fd1qd1_hd z_reg_17_ ( .D(n1241), .CK(i_CLK), .Q(n1333) );
  fd1qd1_hd z_reg_18_ ( .D(n1242), .CK(i_CLK), .Q(n1334) );
  fd1qd1_hd z_reg_19_ ( .D(n1243), .CK(i_CLK), .Q(n1335) );
  fd1qd1_hd z_reg_20_ ( .D(n1244), .CK(i_CLK), .Q(n1336) );
  fd1qd1_hd z_reg_21_ ( .D(n1245), .CK(i_CLK), .Q(n1337) );
  fd1qd1_hd z_reg_22_ ( .D(n1246), .CK(i_CLK), .Q(n1338) );
  fd1qd1_hd z_reg_29_ ( .D(n1253), .CK(i_CLK), .Q(n1345) );
  fd1qd1_hd z_reg_27_ ( .D(n1251), .CK(i_CLK), .Q(n1343) );
  fd1qd1_hd z_reg_25_ ( .D(n1249), .CK(i_CLK), .Q(n1341) );
  fd1qd1_hd z_reg_23_ ( .D(n1247), .CK(i_CLK), .Q(n1339) );
  fd1qd1_hd z_reg_30_ ( .D(n1254), .CK(i_CLK), .Q(n1346) );
  fd1qd1_hd z_reg_28_ ( .D(n1252), .CK(i_CLK), .Q(n1344) );
  fd1qd1_hd z_reg_26_ ( .D(n1250), .CK(i_CLK), .Q(n1342) );
  fd1qd1_hd z_reg_24_ ( .D(n1248), .CK(i_CLK), .Q(n1340) );
  fd1qd1_hd z_m_reg_20_ ( .D(n1219), .CK(i_CLK), .Q(n1372) );
  fd1qd1_hd z_m_reg_16_ ( .D(n1215), .CK(i_CLK), .Q(n1368) );
  fd1qd1_hd z_m_reg_12_ ( .D(n1211), .CK(i_CLK), .Q(n1364) );
  fd1qd1_hd z_m_reg_18_ ( .D(n1217), .CK(i_CLK), .Q(n1370) );
  fd1qd1_hd z_m_reg_14_ ( .D(n1213), .CK(i_CLK), .Q(n1366) );
  fd1qd1_hd z_m_reg_10_ ( .D(n1209), .CK(i_CLK), .Q(n1362) );
  fd1qd1_hd z_m_reg_19_ ( .D(n1218), .CK(i_CLK), .Q(n1371) );
  fd1qd1_hd z_m_reg_15_ ( .D(n1214), .CK(i_CLK), .Q(n1367) );
  fd1qd1_hd z_m_reg_11_ ( .D(n1210), .CK(i_CLK), .Q(n1363) );
  fd1qd1_hd z_m_reg_21_ ( .D(n1220), .CK(i_CLK), .Q(n1373) );
  fd1qd1_hd z_m_reg_17_ ( .D(n1216), .CK(i_CLK), .Q(n1369) );
  fd1qd1_hd z_m_reg_13_ ( .D(n1212), .CK(i_CLK), .Q(n1365) );
  fd1qd1_hd z_m_reg_9_ ( .D(n1208), .CK(i_CLK), .Q(n1361) );
  fd1qd1_hd z_m_reg_22_ ( .D(n1221), .CK(i_CLK), .Q(n1374) );
  fd1qd1_hd z_m_reg_8_ ( .D(n1207), .CK(i_CLK), .Q(n1360) );
  fd1qd1_hd z_m_reg_4_ ( .D(n1203), .CK(i_CLK), .Q(n1356) );
  fd1qd1_hd z_m_reg_0_ ( .D(n1199), .CK(i_CLK), .Q(n1352) );
  fd1qd1_hd z_m_reg_2_ ( .D(n1201), .CK(i_CLK), .Q(n1354) );
  fd1qd1_hd z_m_reg_6_ ( .D(n1205), .CK(i_CLK), .Q(n1358) );
  fd1qd1_hd z_m_reg_7_ ( .D(n1206), .CK(i_CLK), .Q(n1359) );
  fd1qd1_hd z_m_reg_23_ ( .D(n1198), .CK(i_CLK), .Q(n1375) );
  fd1qd1_hd z_m_reg_3_ ( .D(n1202), .CK(i_CLK), .Q(n1355) );
  fd1qd1_hd z_m_reg_1_ ( .D(n1200), .CK(i_CLK), .Q(n1353) );
  fd1qd1_hd z_m_reg_5_ ( .D(n1204), .CK(i_CLK), .Q(n1357) );
  fd1qd1_hd b_e_reg_9_ ( .D(n1112), .CK(i_CLK), .Q(n1452) );
  fd1qd1_hd b_e_reg_8_ ( .D(n1126), .CK(i_CLK), .Q(n1451) );
  fd1qd1_hd z_e_reg_9_ ( .D(n1188), .CK(i_CLK), .Q(n1385) );
  fd1qd1_hd z_e_reg_8_ ( .D(n1197), .CK(i_CLK), .Q(n1384) );
  fd1qd1_hd z_e_reg_4_ ( .D(n1193), .CK(i_CLK), .Q(n1380) );
  fd1qd1_hd z_e_reg_2_ ( .D(n1191), .CK(i_CLK), .Q(n1378) );
  fd1qd1_hd z_e_reg_3_ ( .D(n1192), .CK(i_CLK), .Q(n1379) );
  fd1qd1_hd z_e_reg_7_ ( .D(n1196), .CK(i_CLK), .Q(n1383) );
  fd1qd1_hd a_e_reg_9_ ( .D(n1127), .CK(i_CLK), .Q(n1489) );
  fd1qd1_hd z_e_reg_6_ ( .D(n1195), .CK(i_CLK), .Q(n1382) );
  fd1qd1_hd z_e_reg_1_ ( .D(n1190), .CK(i_CLK), .Q(n1377) );
  fd1qd1_hd a_e_reg_8_ ( .D(n1136), .CK(i_CLK), .Q(n1488) );
  fd1qd1_hd z_e_reg_5_ ( .D(n1194), .CK(i_CLK), .Q(n1381) );
  fd1qd1_hd b_e_reg_6_ ( .D(n1124), .CK(i_CLK), .Q(n1449) );
  fd1qd1_hd a_e_reg_5_ ( .D(n1133), .CK(i_CLK), .Q(n1485) );
  fd1qd1_hd state_reg_3_ ( .D(n1111), .CK(i_CLK), .Q(n[1557]) );
  fd1qd1_hd state_reg_2_ ( .D(n1116), .CK(i_CLK), .Q(n[1556]) );
  fd1qd1_hd state_reg_1_ ( .D(n1115), .CK(i_CLK), .Q(n[1555]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n1123), .CK(i_CLK), .Q(n1448) );
  fd1qd1_hd a_e_reg_7_ ( .D(n1135), .CK(i_CLK), .Q(n1487) );
  fd1qd1_hd a_e_reg_1_ ( .D(n1129), .CK(i_CLK), .Q(n1481) );
  fd1qd1_hd b_e_reg_1_ ( .D(n1119), .CK(i_CLK), .Q(n1444) );
  fd1qd1_hd state_reg_0_ ( .D(n1114), .CK(i_CLK), .Q(n[1554]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n1128), .CK(i_CLK), .Q(n1480) );
  fd1qd1_hd a_e_reg_2_ ( .D(n1130), .CK(i_CLK), .Q(n1482) );
  fd1qd1_hd b_e_reg_7_ ( .D(n1125), .CK(i_CLK), .Q(n1450) );
  fd1qd1_hd b_e_reg_4_ ( .D(n1122), .CK(i_CLK), .Q(n1447) );
  fd1qd1_hd a_e_reg_4_ ( .D(n1132), .CK(i_CLK), .Q(n1484) );
  fd1qd1_hd a_e_reg_6_ ( .D(n1134), .CK(i_CLK), .Q(n1486) );
  fd1qd1_hd b_e_reg_2_ ( .D(n1120), .CK(i_CLK), .Q(n1445) );
  fd1qd1_hd b_m_reg_25_ ( .D(n1113), .CK(i_CLK), .Q(n1441) );
  fd1qd1_hd a_m_reg_24_ ( .D(n1162), .CK(i_CLK), .Q(n1477) );
  fd1qd1_hd b_m_reg_24_ ( .D(n1187), .CK(i_CLK), .Q(n1440) );
  fd1qd1_hd b_m_reg_21_ ( .D(n1184), .CK(i_CLK), .Q(n1437) );
  fd1qd1_hd a_m_reg_23_ ( .D(n1161), .CK(i_CLK), .Q(n1476) );
  fd1qd1_hd b_m_reg_15_ ( .D(n1178), .CK(i_CLK), .Q(n1431) );
  fd1qd1_hd b_m_reg_16_ ( .D(n1179), .CK(i_CLK), .Q(n1432) );
  fd1qd1_hd b_m_reg_13_ ( .D(n1176), .CK(i_CLK), .Q(n1429) );
  fd1qd1_hd b_m_reg_18_ ( .D(n1181), .CK(i_CLK), .Q(n1434) );
  fd1qd1_hd b_m_reg_19_ ( .D(n1182), .CK(i_CLK), .Q(n1435) );
  fd1qd1_hd b_m_reg_17_ ( .D(n1180), .CK(i_CLK), .Q(n1433) );
  fd1qd1_hd a_m_reg_21_ ( .D(n1159), .CK(i_CLK), .Q(n1474) );
  fd1qd1_hd b_m_reg_14_ ( .D(n1177), .CK(i_CLK), .Q(n1430) );
  fd1qd1_hd a_m_reg_19_ ( .D(n1157), .CK(i_CLK), .Q(n1472) );
  fd1qd1_hd a_m_reg_22_ ( .D(n1160), .CK(i_CLK), .Q(n1475) );
  fd1qd1_hd b_m_reg_23_ ( .D(n1186), .CK(i_CLK), .Q(n1439) );
  fd1qd1_hd a_m_reg_20_ ( .D(n1158), .CK(i_CLK), .Q(n1473) );
  fd1qd1_hd b_m_reg_7_ ( .D(n1170), .CK(i_CLK), .Q(n1423) );
  fd1qd1_hd b_m_reg_22_ ( .D(n1185), .CK(i_CLK), .Q(n1438) );
  fd1qd1_hd b_m_reg_20_ ( .D(n1183), .CK(i_CLK), .Q(n1436) );
  fd1qd1_hd a_m_reg_0_ ( .D(n1138), .CK(i_CLK), .Q(n1453) );
  fd1qd1_hd a_m_reg_1_ ( .D(n1139), .CK(i_CLK), .Q(n1454) );
  fd1qd1_hd a_m_reg_2_ ( .D(n1140), .CK(i_CLK), .Q(n1455) );
  fd1qd1_hd a_m_reg_7_ ( .D(n1145), .CK(i_CLK), .Q(n1460) );
  fd1qd1_hd b_m_reg_0_ ( .D(n1163), .CK(i_CLK), .Q(n1416) );
  fd1qd1_hd a_m_reg_5_ ( .D(n1143), .CK(i_CLK), .Q(n1458) );
  fd1qd1_hd a_m_reg_3_ ( .D(n1141), .CK(i_CLK), .Q(n1456) );
  fd1qd1_hd b_m_reg_3_ ( .D(n1166), .CK(i_CLK), .Q(n1419) );
  fd1qd1_hd b_m_reg_6_ ( .D(n1169), .CK(i_CLK), .Q(n1422) );
  fd1qd1_hd b_m_reg_4_ ( .D(n1167), .CK(i_CLK), .Q(n1420) );
  fd1qd1_hd b_m_reg_1_ ( .D(n1164), .CK(i_CLK), .Q(n1417) );
  fd1qd1_hd b_m_reg_2_ ( .D(n1165), .CK(i_CLK), .Q(n1418) );
  fd1qd1_hd b_m_reg_5_ ( .D(n1168), .CK(i_CLK), .Q(n1421) );
  fd1qd1_hd a_m_reg_4_ ( .D(n1142), .CK(i_CLK), .Q(n1457) );
  fd1qd1_hd a_m_reg_6_ ( .D(n1144), .CK(i_CLK), .Q(n1459) );
  fad1_hd DP_OP_43J1_124_6938_U28 ( .A(n1083), .B(n77), .CI(n1082), .CO(n1055), 
        .S(n1315) );
  fad1_hd DP_OP_43J1_124_6938_U25 ( .A(n1079), .B(n1086), .CI(n1053), .CO(
        n1052), .S(n1312) );
  fad1_hd DP_OP_43J1_124_6938_U23 ( .A(n1077), .B(n1088), .CI(n1051), .CO(
        n1050), .S(n1310) );
  fad1_hd DP_OP_43J1_124_6938_U27 ( .A(n1081), .B(n1084), .CI(n1055), .CO(
        n1054), .S(n1314) );
  fad1_hd DP_OP_43J1_124_6938_U26 ( .A(n1080), .B(n1085), .CI(n1054), .CO(
        n1053), .S(n1313) );
  fad1_hd DP_OP_43J1_124_6938_U24 ( .A(n1078), .B(n1087), .CI(n1052), .CO(
        n1051), .S(n1311) );
  fad1_hd DP_OP_43J1_124_6938_U22 ( .A(n1076), .B(n1089), .CI(n1050), .CO(
        n1049), .S(n1309) );
  fad1_hd DP_OP_43J1_124_6938_U21 ( .A(n1075), .B(n1090), .CI(n1049), .CO(
        n1048), .S(n1308) );
  fad1_hd DP_OP_43J1_124_6938_U2 ( .A(n1056), .B(n1109), .CI(n1030), .CO(n1029), .S(n1289) );
  fad1_hd DP_OP_43J1_124_6938_U3 ( .A(n1057), .B(n1108), .CI(n1031), .CO(n1030), .S(n1290) );
  fad1_hd DP_OP_43J1_124_6938_U4 ( .A(n1058), .B(n1107), .CI(n1032), .CO(n1031), .S(n1291) );
  fad1_hd DP_OP_43J1_124_6938_U15 ( .A(n1069), .B(n1096), .CI(n1043), .CO(
        n1042), .S(n1302) );
  fad1_hd DP_OP_43J1_124_6938_U16 ( .A(n1070), .B(n1095), .CI(n1044), .CO(
        n1043), .S(n1303) );
  fad1_hd DP_OP_43J1_124_6938_U17 ( .A(n1071), .B(n1094), .CI(n1045), .CO(
        n1044), .S(n1304) );
  fad1_hd DP_OP_43J1_124_6938_U18 ( .A(n1072), .B(n1093), .CI(n1046), .CO(
        n1045), .S(n1305) );
  fad1_hd DP_OP_43J1_124_6938_U19 ( .A(n1073), .B(n1092), .CI(n1047), .CO(
        n1046), .S(n1306) );
  fad1_hd DP_OP_43J1_124_6938_U20 ( .A(n1074), .B(n1091), .CI(n1048), .CO(
        n1047), .S(n1307) );
  fad1_hd DP_OP_43J1_124_6938_U14 ( .A(n1068), .B(n1097), .CI(n1042), .CO(
        n1041), .S(n1301) );
  fad1_hd DP_OP_43J1_124_6938_U13 ( .A(n1067), .B(n1098), .CI(n1041), .CO(
        n1040), .S(n1300) );
  fad1_hd DP_OP_43J1_124_6938_U12 ( .A(n1066), .B(n1099), .CI(n1040), .CO(
        n1039), .S(n1299) );
  fad1_hd DP_OP_43J1_124_6938_U11 ( .A(n1065), .B(n1100), .CI(n1039), .CO(
        n1038), .S(n1298) );
  fad1_hd DP_OP_43J1_124_6938_U10 ( .A(n1064), .B(n1101), .CI(n1038), .CO(
        n1037), .S(n1297) );
  fad1_hd DP_OP_43J1_124_6938_U9 ( .A(n1063), .B(n1102), .CI(n1037), .CO(n1036), .S(n1296) );
  fad1_hd DP_OP_43J1_124_6938_U8 ( .A(n1062), .B(n1103), .CI(n1036), .CO(n1035), .S(n1295) );
  fad1_hd DP_OP_43J1_124_6938_U7 ( .A(n1061), .B(n1104), .CI(n1035), .CO(n1034), .S(n1294) );
  fad1_hd DP_OP_43J1_124_6938_U6 ( .A(n1060), .B(n1105), .CI(n1034), .CO(n1033), .S(n1293) );
  fad1_hd DP_OP_43J1_124_6938_U5 ( .A(n1059), .B(n1106), .CI(n1033), .CO(n1032), .S(n1292) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n1117), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd o_Z_STB_reg ( .D(n1110), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd sticky_reg ( .D(n1223), .CK(i_CLK), .Q(n1349) );
  fd1qd1_hd round_bit_reg ( .D(n1222), .CK(i_CLK), .Q(n1350) );
  fd1qd1_hd a_m_reg_17_ ( .D(n1155), .CK(i_CLK), .Q(n1470) );
  fd1qd1_hd a_m_reg_16_ ( .D(n1154), .CK(i_CLK), .Q(n1469) );
  fd1qd1_hd b_m_reg_8_ ( .D(n1171), .CK(i_CLK), .Q(n1424) );
  fd1qd1_hd b_m_reg_12_ ( .D(n1175), .CK(i_CLK), .Q(n1428) );
  fd1qd1_hd b_m_reg_11_ ( .D(n1174), .CK(i_CLK), .Q(n1427) );
  fd1qd1_hd b_m_reg_10_ ( .D(n1173), .CK(i_CLK), .Q(n1426) );
  fd1qd1_hd b_m_reg_9_ ( .D(n1172), .CK(i_CLK), .Q(n1425) );
  fd1qd1_hd a_m_reg_14_ ( .D(n1152), .CK(i_CLK), .Q(n1467) );
  fd1qd1_hd a_m_reg_13_ ( .D(n1151), .CK(i_CLK), .Q(n1466) );
  fd1qd1_hd a_m_reg_15_ ( .D(n1153), .CK(i_CLK), .Q(n1468) );
  fd1qd1_hd a_m_reg_18_ ( .D(n1156), .CK(i_CLK), .Q(n1471) );
  fd1qd1_hd a_m_reg_12_ ( .D(n1150), .CK(i_CLK), .Q(n1465) );
  fd1qd1_hd a_m_reg_11_ ( .D(n1149), .CK(i_CLK), .Q(n1464) );
  fd1qd1_hd a_m_reg_10_ ( .D(n1148), .CK(i_CLK), .Q(n1463) );
  fd1qd1_hd a_m_reg_9_ ( .D(n1147), .CK(i_CLK), .Q(n1462) );
  fd1qd1_hd a_m_reg_8_ ( .D(n1146), .CK(i_CLK), .Q(n1461) );
  fd1qd1_hd a_m_reg_25_ ( .D(n1137), .CK(i_CLK), .Q(n1478) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(n1339), .E(n16), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(n1333), .E(n16), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(n1329), .E(n5), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(n1316), .E(n200), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n9), .CK(i_CLK), .Q(n1513) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n11), .CK(i_CLK), .Q(n1550) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(n1347), .E(n15), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(n1346), .E(n15), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(n1331), .E(n14), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(n1328), .E(n202), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n19), .CK(i_CLK), .Q(n1505) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n3), .CK(i_CLK), .Q(n1495) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n9), .CK(i_CLK), .Q(n1551) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n8), .CK(i_CLK), .Q(n1532) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n3), .CK(i_CLK), .Q(n1521) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n3), .CK(i_CLK), .Q(n1508) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n19), .CK(i_CLK), .Q(n1502) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n9), .CK(i_CLK), .Q(n1500) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n206), .CK(i_CLK), .Q(n1499) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n206), .CK(i_CLK), .Q(n1497) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n9), .CK(i_CLK), .Q(n1493) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n6), .CK(i_CLK), .Q(n1490) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n18), .CK(i_CLK), .Q(n1547) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n18), .CK(i_CLK), .Q(n1533) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n11), .CK(i_CLK), .Q(n1531) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n10), .CK(i_CLK), .Q(n1530) );
  fd1eqd1_hd b_s_reg ( .D(n1521), .E(n181), .CK(i_CLK), .Q(n1414) );
  fd1eqd1_hd a_s_reg ( .D(n1553), .E(n181), .CK(i_CLK), .Q(n1415) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(n1332), .E(n202), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(n1330), .E(n5), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(n1318), .E(n16), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(n1345), .E(n5), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(n1343), .E(n202), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(n1342), .E(n200), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(n1341), .E(n15), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(n1322), .E(n14), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(n1321), .E(n5), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n7), .CK(i_CLK), .Q(n1516) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n17), .CK(i_CLK), .Q(n1553) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n10), .CK(i_CLK), .Q(n1544) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n19), .CK(i_CLK), .Q(n1535) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n6), .CK(i_CLK), .Q(n1520) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n18), .CK(i_CLK), .Q(n1519) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n9), .CK(i_CLK), .Q(n1518) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n206), .CK(i_CLK), .Q(n1517) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n6), .CK(i_CLK), .Q(n1515) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n11), .CK(i_CLK), .Q(n1514) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n8), .CK(i_CLK), .Q(n1512) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n8), .CK(i_CLK), .Q(n1511) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n7), .CK(i_CLK), .Q(n1510) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n206), .CK(i_CLK), .Q(n1509) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n9), .CK(i_CLK), .Q(n1507) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n19), .CK(i_CLK), .Q(n1506) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n18), .CK(i_CLK), .Q(n1504) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n7), .CK(i_CLK), .Q(n1503) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n3), .CK(i_CLK), .Q(n1501) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n17), .CK(i_CLK), .Q(n1498) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n11), .CK(i_CLK), .Q(n1496) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n10), .CK(i_CLK), .Q(n1494) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n11), .CK(i_CLK), .Q(n1492) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n7), .CK(i_CLK), .Q(n1491) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n10), .CK(i_CLK), .Q(n1552) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n6), .CK(i_CLK), .Q(n1549) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n17), .CK(i_CLK), .Q(n1548) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n8), .CK(i_CLK), .Q(n1546) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n18), .CK(i_CLK), .Q(n1545) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n7), .CK(i_CLK), .Q(n1543) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n17), .CK(i_CLK), .Q(n1542) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n11), .CK(i_CLK), .Q(n1541) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n7), .CK(i_CLK), .Q(n1540) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n10), .CK(i_CLK), .Q(n1539) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n18), .CK(i_CLK), .Q(n1538) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n3), .CK(i_CLK), .Q(n1537) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n10), .CK(i_CLK), .Q(n1536) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n8), .CK(i_CLK), .Q(n1534) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n19), .CK(i_CLK), .Q(n1529) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n8), .CK(i_CLK), .Q(n1528) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n17), .CK(i_CLK), .Q(n1527) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n206), .CK(i_CLK), .Q(n1526) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n3), .CK(i_CLK), .Q(n1525) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n17), .CK(i_CLK), .Q(n1524) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n6), .CK(i_CLK), .Q(n1523) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n19), .CK(i_CLK), .Q(n1522) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(n1340), .E(n5), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(n1324), .E(n200), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(n1319), .E(n16), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(n1344), .E(n14), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(n1338), .E(n14), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(n1337), .E(n200), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(n1336), .E(n15), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(n1335), .E(n16), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(n1334), .E(n16), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(n1327), .E(n5), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(n1326), .E(n200), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(n1325), .E(n15), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(n1323), .E(n15), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(n1320), .E(n14), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(n1317), .E(n202), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd guard_reg ( .D(n1256), .E(n1257), .CK(i_CLK), .Q(n1351) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n56), .E(n1276), .CK(i_CLK), .Q(n1442) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n57), .E(n1277), .CK(i_CLK), .Q(n1479) );
  fd1eqd1_hd z_s_reg ( .D(n1287), .E(n13), .CK(i_CLK), .Q(n1348) );
  fd1eqd1_hd sum_reg_0_ ( .D(n1315), .E(n204), .CK(i_CLK), .Q(n1386) );
  fd1eqd1_hd sum_reg_1_ ( .D(n1314), .E(n4), .CK(i_CLK), .Q(n1387) );
  fd1eqd1_hd sum_reg_2_ ( .D(n1313), .E(n12), .CK(i_CLK), .Q(n1388) );
  fd1eqd1_hd sum_reg_3_ ( .D(n1312), .E(n205), .CK(i_CLK), .Q(n1389) );
  fd1eqd1_hd sum_reg_4_ ( .D(n1311), .E(n4), .CK(i_CLK), .Q(n1390) );
  fd1eqd1_hd sum_reg_5_ ( .D(n1310), .E(n12), .CK(i_CLK), .Q(n1391) );
  fd1eqd1_hd sum_reg_6_ ( .D(n1309), .E(n13), .CK(i_CLK), .Q(n1392) );
  fd1eqd1_hd sum_reg_7_ ( .D(n1308), .E(n204), .CK(i_CLK), .Q(n1393) );
  fd1eqd1_hd sum_reg_8_ ( .D(n1307), .E(n12), .CK(i_CLK), .Q(n1394) );
  fd1eqd1_hd sum_reg_9_ ( .D(n1306), .E(n13), .CK(i_CLK), .Q(n1395) );
  fd1eqd1_hd sum_reg_10_ ( .D(n1305), .E(n4), .CK(i_CLK), .Q(n1396) );
  fd1eqd1_hd sum_reg_11_ ( .D(n1304), .E(n4), .CK(i_CLK), .Q(n1397) );
  fd1eqd1_hd sum_reg_12_ ( .D(n1303), .E(n13), .CK(i_CLK), .Q(n1398) );
  fd1eqd1_hd sum_reg_13_ ( .D(n1302), .E(n205), .CK(i_CLK), .Q(n1399) );
  fd1eqd1_hd sum_reg_14_ ( .D(n1301), .E(n205), .CK(i_CLK), .Q(n1400) );
  fd1eqd1_hd sum_reg_15_ ( .D(n1300), .E(n12), .CK(i_CLK), .Q(n1401) );
  fd1eqd1_hd sum_reg_16_ ( .D(n1299), .E(n205), .CK(i_CLK), .Q(n1402) );
  fd1eqd1_hd sum_reg_17_ ( .D(n1298), .E(n203), .CK(i_CLK), .Q(n1403) );
  fd1eqd1_hd sum_reg_18_ ( .D(n1297), .E(n205), .CK(i_CLK), .Q(n1404) );
  fd1eqd1_hd sum_reg_19_ ( .D(n1296), .E(n13), .CK(i_CLK), .Q(n1405) );
  fd1eqd1_hd sum_reg_20_ ( .D(n1295), .E(n203), .CK(i_CLK), .Q(n1406) );
  fd1eqd1_hd sum_reg_21_ ( .D(n1294), .E(n204), .CK(i_CLK), .Q(n1407) );
  fd1eqd1_hd sum_reg_22_ ( .D(n1293), .E(n4), .CK(i_CLK), .Q(n1408) );
  fd1eqd1_hd sum_reg_23_ ( .D(n1292), .E(n204), .CK(i_CLK), .Q(n1409) );
  fd1eqd1_hd sum_reg_24_ ( .D(n1291), .E(n204), .CK(i_CLK), .Q(n1410) );
  fd1eqd1_hd sum_reg_25_ ( .D(n1290), .E(n4), .CK(i_CLK), .Q(n1411) );
  fd1eqd1_hd sum_reg_26_ ( .D(n1289), .E(n12), .CK(i_CLK), .Q(n1412) );
  fd1eqd1_hd sum_reg_27_ ( .D(n1288), .E(n203), .CK(i_CLK), .Q(n1413) );
  clknd2d1_hd U523 ( .A(n781), .B(n780), .Y(n783) );
  clknd2d1_hd U524 ( .A(n770), .B(n769), .Y(n804) );
  clknd2d1_hd U525 ( .A(n59), .B(n950), .Y(n769) );
  clknd2d1_hd U526 ( .A(n1437), .B(n981), .Y(n776) );
  clknd2d1_hd U527 ( .A(n237), .B(n236), .Y(n252) );
  clknd2d1_hd U528 ( .A(n1448), .B(n914), .Y(n237) );
  clknd2d1_hd U529 ( .A(n1447), .B(n916), .Y(n236) );
  clknd2d1_hd U530 ( .A(n1449), .B(n919), .Y(n246) );
  clknd2d1_hd U531 ( .A(n1444), .B(n908), .Y(n245) );
  clknd2d1_hd U532 ( .A(n1275), .B(n[1556]), .Y(n558) );
  clknd2d1_hd U533 ( .A(n825), .B(n547), .Y(n527) );
  clknd2d1_hd U534 ( .A(n1478), .B(n992), .Y(n816) );
  clknd2d1_hd U535 ( .A(n1450), .B(n328), .Y(n209) );
  clknd2d1_hd U536 ( .A(n244), .B(n66), .Y(n526) );
  clknd2d1_hd U537 ( .A(n247), .B(n241), .Y(n242) );
  nid1_hd U538 ( .A(n1012), .Y(n192) );
  clknd2d1_hd U539 ( .A(n253), .B(n49), .Y(n525) );
  clknd2d1_hd U540 ( .A(n244), .B(n253), .Y(n313) );
  clknd2d1_hd U541 ( .A(n49), .B(n508), .Y(n564) );
  clknd2d1_hd U542 ( .A(n1257), .B(n896), .Y(n659) );
  clknd2d1_hd U543 ( .A(n359), .B(n343), .Y(n221) );
  clknd2d1_hd U544 ( .A(n1383), .B(n1384), .Y(n559) );
  nid1_hd U545 ( .A(n180), .Y(n179) );
  nid2_hd U546 ( .A(n1010), .Y(n180) );
  ivd1_hd U547 ( .A(n170), .Y(n163) );
  ivd1_hd U548 ( .A(n179), .Y(n164) );
  nid1_hd U549 ( .A(n169), .Y(n173) );
  nid1_hd U550 ( .A(n178), .Y(n170) );
  nid1_hd U551 ( .A(n179), .Y(n175) );
  nid1_hd U552 ( .A(n180), .Y(n178) );
  nid1_hd U553 ( .A(n169), .Y(n174) );
  ivd1_hd U554 ( .A(n179), .Y(n165) );
  nid1_hd U555 ( .A(n178), .Y(n171) );
  nid1_hd U556 ( .A(n1006), .Y(n99) );
  nid1_hd U557 ( .A(n180), .Y(n176) );
  nid1_hd U558 ( .A(n1006), .Y(n145) );
  nid1_hd U559 ( .A(n178), .Y(n172) );
  nid1_hd U560 ( .A(n172), .Y(n177) );
  ivd1_hd U561 ( .A(n171), .Y(n161) );
  nid1_hd U562 ( .A(n179), .Y(n169) );
  nid1_hd U563 ( .A(n1272), .Y(n1019) );
  ivd1_hd U564 ( .A(n1479), .Y(n998) );
  nid1_hd U565 ( .A(n763), .Y(n154) );
  clknd2d1_hd U566 ( .A(n73), .B(n135), .Y(n739) );
  clknd2d1_hd U567 ( .A(n72), .B(n151), .Y(n763) );
  nid1_hd U568 ( .A(n202), .Y(n201) );
  nid1_hd U569 ( .A(n123), .Y(n151) );
  nid1_hd U570 ( .A(n763), .Y(n152) );
  nid1_hd U571 ( .A(n144), .Y(n138) );
  nid1_hd U572 ( .A(n739), .Y(n144) );
  nid1_hd U573 ( .A(n144), .Y(n139) );
  nid1_hd U574 ( .A(n152), .Y(n155) );
  nid1_hd U575 ( .A(n152), .Y(n153) );
  nid1_hd U576 ( .A(n144), .Y(n137) );
  clknd2d1_hd U577 ( .A(n357), .B(n1515), .Y(n349) );
  clknd2d1_hd U578 ( .A(n273), .B(n271), .Y(n268) );
  nid1_hd U579 ( .A(n1012), .Y(n191) );
  clknd2d1_hd U580 ( .A(n344), .B(n341), .Y(n338) );
  clknd2d1_hd U581 ( .A(n300), .B(n1547), .Y(n292) );
  clknd2d1_hd U582 ( .A(n306), .B(n302), .Y(n303) );
  clknd2d1_hd U583 ( .A(n508), .B(n66), .Y(n510) );
  clknd2d1_hd U584 ( .A(n67), .B(n509), .Y(n920) );
  clknd2d1_hd U585 ( .A(n57), .B(n534), .Y(n511) );
  clknd2d1_hd U586 ( .A(n358), .B(n360), .Y(n354) );
  clknd2d1_hd U587 ( .A(n301), .B(n303), .Y(n296) );
  clknd2d1_hd U588 ( .A(n57), .B(n301), .Y(n307) );
  clknd2d1_hd U589 ( .A(n94), .B(n333), .Y(n327) );
  clknd2d1_hd U590 ( .A(n54), .B(n328), .Y(n326) );
  clknd2d1_hd U591 ( .A(n1660), .B(n1268), .Y(n1269) );
  clknd2d1_hd U592 ( .A(n1484), .B(n277), .Y(n272) );
  clknd2d1_hd U593 ( .A(n306), .B(n914), .Y(n271) );
  clknd2d1_hd U594 ( .A(n278), .B(n1550), .Y(n274) );
  clknd2d1_hd U595 ( .A(n335), .B(n1518), .Y(n330) );
  clknd2d1_hd U596 ( .A(n329), .B(n326), .Y(n323) );
  clknd2d1_hd U597 ( .A(n1486), .B(n262), .Y(n764) );
  clknd2d1_hd U598 ( .A(n267), .B(n260), .Y(n766) );
  clknd2d1_hd U599 ( .A(n66), .B(n889), .Y(n918) );
  clknd2d1_hd U600 ( .A(n92), .B(n319), .Y(n921) );
  clknd2d1_hd U601 ( .A(n322), .B(n317), .Y(n923) );
  clknd2d1_hd U602 ( .A(n660), .B(n685), .Y(n666) );
  clknd2d1_hd U603 ( .A(n63), .B(n711), .Y(n707) );
  clknd2d1_hd U604 ( .A(n931), .B(n1413), .Y(n894) );
  clknd2d1_hd U605 ( .A(n65), .B(n698), .Y(n691) );
  clknd2d1_hd U606 ( .A(n61), .B(n65), .Y(n684) );
  clknd2d1_hd U607 ( .A(n936), .B(n60), .Y(n567) );
  nid1_hd U608 ( .A(n705), .Y(n142) );
  clknd2d1_hd U609 ( .A(n635), .B(n685), .Y(n642) );
  clknd2d1_hd U610 ( .A(n612), .B(n65), .Y(n618) );
  clknd2d1_hd U611 ( .A(n589), .B(n65), .Y(n595) );
  clknd2d1_hd U612 ( .A(n569), .B(n685), .Y(n708) );
  nid1_hd U613 ( .A(n159), .Y(n156) );
  nid1_hd U614 ( .A(n932), .Y(n159) );
  nid1_hd U615 ( .A(n705), .Y(n141) );
  nid1_hd U616 ( .A(n932), .Y(n157) );
  nid1_hd U617 ( .A(n159), .Y(n158) );
  nid1_hd U618 ( .A(n705), .Y(n140) );
  clknd2d1_hd U619 ( .A(n873), .B(n872), .Y(n871) );
  clknd2d1_hd U620 ( .A(n827), .B(n826), .Y(n888) );
  clknd2d1_hd U621 ( .A(n859), .B(n835), .Y(n877) );
  clknd2d1_hd U622 ( .A(n884), .B(n861), .Y(n860) );
  clknd2d1_hd U623 ( .A(n876), .B(n841), .Y(n851) );
  clknd2d1_hd U624 ( .A(n880), .B(n879), .Y(n878) );
  clknd2d1_hd U625 ( .A(n850), .B(n828), .Y(n866) );
  clknd2d1_hd U626 ( .A(n854), .B(n853), .Y(n852) );
  nid1_hd U627 ( .A(n199), .Y(n196) );
  clknd2d1_hd U628 ( .A(n885), .B(n869), .Y(n844) );
  clknd2d1_hd U629 ( .A(n56), .B(n870), .Y(n548) );
  nid1_hd U630 ( .A(n199), .Y(n195) );
  clknd2d1_hd U631 ( .A(n1415), .B(n550), .Y(n533) );
  clknd2d1_hd U632 ( .A(n1445), .B(n311), .Y(n342) );
  clknd2d1_hd U633 ( .A(n55), .B(n343), .Y(n341) );
  clknd2d1_hd U634 ( .A(n346), .B(n1516), .Y(n345) );
  clknd2d1_hd U635 ( .A(n55), .B(n359), .Y(n360) );
  nid1_hd U636 ( .A(n1012), .Y(n193) );
  clknd2d1_hd U637 ( .A(n1482), .B(n255), .Y(n286) );
  clknd2d1_hd U638 ( .A(n306), .B(n910), .Y(n285) );
  clknd2d1_hd U639 ( .A(n289), .B(n1548), .Y(n288) );
  nid1_hd U640 ( .A(n12), .Y(n203) );
  nid1_hd U641 ( .A(n203), .Y(n205) );
  nid1_hd U642 ( .A(n205), .Y(n204) );
  clknd2d1_hd U643 ( .A(n895), .B(n930), .Y(n1257) );
  ivd1_hd U644 ( .A(n1272), .Y(n18) );
  nid1_hd U645 ( .A(n6), .Y(n206) );
  nid1_hd U646 ( .A(n200), .Y(n202) );
  nid1_hd U647 ( .A(n14), .Y(n200) );
  clknd2d1_hd U648 ( .A(n21), .B(n1286), .Y(n935) );
  clknd2d1_hd U649 ( .A(n158), .B(n1387), .Y(n933) );
  clknd2d1_hd U650 ( .A(n95), .B(n262), .Y(n270) );
  clknd2d1_hd U651 ( .A(n274), .B(n263), .Y(n264) );
  clknd2d1_hd U652 ( .A(n95), .B(n277), .Y(n284) );
  clknd2d1_hd U653 ( .A(n55), .B(n333), .Y(n340) );
  clknd2d1_hd U654 ( .A(n304), .B(n303), .Y(n1128) );
  clknd2d1_hd U655 ( .A(n54), .B(n319), .Y(n325) );
  clknd2d1_hd U656 ( .A(n330), .B(n320), .Y(n321) );
  clknd2d1_hd U657 ( .A(n1489), .B(n203), .Y(n900) );
  clknd2d1_hd U658 ( .A(n1020), .B(n899), .Y(n898) );
  clknd2d1_hd U659 ( .A(n115), .B(n691), .Y(n693) );
  clknd2d1_hd U660 ( .A(n696), .B(n691), .Y(n686) );
  clknd2d1_hd U661 ( .A(n875), .B(n874), .Y(n1254) );
  clknd2d1_hd U662 ( .A(n552), .B(n551), .Y(n553) );
  clknd2d1_hd U663 ( .A(n542), .B(n541), .Y(n544) );
  clknd2d1_hd U664 ( .A(n507), .B(n360), .Y(n1118) );
  ivd1_hd U665 ( .A(n1019), .Y(n19) );
  ivd1_hd U666 ( .A(n1019), .Y(n3) );
  ivd1_hd U667 ( .A(n1016), .Y(n4) );
  ivd1_hd U668 ( .A(n1015), .Y(n5) );
  ivd1_hd U669 ( .A(n1019), .Y(n6) );
  ivd1_hd U670 ( .A(n1272), .Y(n7) );
  ivd1_hd U671 ( .A(n1272), .Y(n8) );
  ivd1_hd U672 ( .A(n1019), .Y(n9) );
  ivd1_hd U673 ( .A(n1272), .Y(n10) );
  ivd1_hd U674 ( .A(n1019), .Y(n11) );
  nid1_hd U675 ( .A(n918), .Y(n1016) );
  ivd1_hd U676 ( .A(n1016), .Y(n12) );
  ivd1_hd U677 ( .A(n1016), .Y(n13) );
  or2d1_hd U678 ( .A(n1275), .B(n526), .Y(n1015) );
  ivd1_hd U679 ( .A(n1015), .Y(n14) );
  ivd1_hd U680 ( .A(n1015), .Y(n15) );
  ivd1_hd U681 ( .A(n1015), .Y(n16) );
  ivd1_hd U682 ( .A(n1019), .Y(n17) );
  ivd1_hd U683 ( .A(n1439), .Y(n973) );
  xo2d1_hd U684 ( .A(n79), .B(n1011), .Y(n1065) );
  xo2d1_hd U685 ( .A(n78), .B(n967), .Y(n1067) );
  ao211d1_hd U686 ( .A(n820), .B(n819), .C(n818), .D(n145), .Y(n1010) );
  oa211d1_hd U687 ( .A(n1440), .B(n817), .C(n816), .D(n815), .Y(n819) );
  scg6d1_hd U688 ( .A(n39), .B(n817), .C(n937), .Y(n815) );
  ao211d1_hd U689 ( .A(n1476), .B(n973), .C(n814), .D(n813), .Y(n817) );
  ad4d1_hd U690 ( .A(n302), .B(n308), .C(n904), .D(n219), .Y(n550) );
  xo2d1_hd U691 ( .A(n78), .B(n1029), .Y(n1288) );
  xo2d1_hd U692 ( .A(n78), .B(n982), .Y(n1061) );
  xo2d1_hd U693 ( .A(n79), .B(n1004), .Y(n1060) );
  xo2d1_hd U694 ( .A(n78), .B(n994), .Y(n1057) );
  xo2d1_hd U695 ( .A(n77), .B(n978), .Y(n1062) );
  xo2d1_hd U696 ( .A(n77), .B(n975), .Y(n1059) );
  xo2d1_hd U697 ( .A(n78), .B(n991), .Y(n1080) );
  xo2d1_hd U698 ( .A(n79), .B(n963), .Y(n1078) );
  xo2d1_hd U699 ( .A(n78), .B(n997), .Y(n1075) );
  xo2d1_hd U700 ( .A(n77), .B(n986), .Y(n1076) );
  xo2d1_hd U701 ( .A(n79), .B(n958), .Y(n1072) );
  xo2d1_hd U702 ( .A(n77), .B(n970), .Y(n1069) );
  nid1_hd U703 ( .A(n844), .Y(n557) );
  scg6d1_hd U704 ( .A(n897), .B(n1013), .C(n70), .Y(n926) );
  or2d1_hd U705 ( .A(n1028), .B(n64), .Y(n701) );
  or2d1_hd U706 ( .A(n313), .B(n334), .Y(n515) );
  scg10d1_hd U707 ( .A(n302), .B(n301), .C(n193), .D(n1545), .Y(n304) );
  ad2d1_hd U708 ( .A(n56), .B(n358), .Y(n516) );
  scg10d1_hd U709 ( .A(n359), .B(n358), .C(n193), .D(n1513), .Y(n507) );
  ad2d1_hd U710 ( .A(n21), .B(n51), .Y(n697) );
  nid1_hd U711 ( .A(n737), .Y(n135) );
  nid1_hd U712 ( .A(n199), .Y(n198) );
  nid1_hd U713 ( .A(n194), .Y(n199) );
  nid1_hd U714 ( .A(n194), .Y(n197) );
  nid1_hd U715 ( .A(n1014), .Y(n194) );
  scg6d1_hd U716 ( .A(n72), .B(n254), .C(n189), .Y(n737) );
  ad3d1_hd U717 ( .A(n511), .B(n510), .C(n920), .Y(n1265) );
  scg2d1_hd U718 ( .A(n1375), .B(n121), .C(n201), .D(n1259), .Y(n1261) );
  nid1_hd U719 ( .A(n705), .Y(n143) );
  or2d1_hd U720 ( .A(n[1557]), .B(n526), .Y(n1273) );
  or2d1_hd U721 ( .A(n[1556]), .B(n525), .Y(n1012) );
  or2d1_hd U722 ( .A(n1275), .B(n920), .Y(n896) );
  or4d1_hd U723 ( .A(n1477), .B(n230), .C(n229), .D(n228), .Y(n529) );
  nr2bd1_hd U724 ( .AN(n823), .B(n824), .Y(n556) );
  scg2d1_hd U725 ( .A(n968), .B(n1466), .C(n954), .D(n799), .Y(n801) );
  or3d1_hd U726 ( .A(n67), .B(n49), .C(n558), .Y(n1018) );
  nid1_hd U727 ( .A(n1006), .Y(n100) );
  ad2d1_hd U728 ( .A(n1546), .B(n1545), .Y(n300) );
  ad2d1_hd U729 ( .A(n1514), .B(n1513), .Y(n357) );
  ad2d1_hd U730 ( .A(o_Z_STB), .B(i_Z_ACK), .Y(n1259) );
  ivd1_hd U731 ( .A(n1018), .Y(n20) );
  ivd1_hd U732 ( .A(n1018), .Y(n21) );
  ivd1_hd U733 ( .A(n516), .Y(n22) );
  ivd1_hd U734 ( .A(n516), .Y(n23) );
  ivd1_hd U735 ( .A(n1456), .Y(n24) );
  ivd1_hd U736 ( .A(n24), .Y(n25) );
  ivd1_hd U737 ( .A(n1469), .Y(n26) );
  ivd1_hd U738 ( .A(n26), .Y(n27) );
  ivd1_hd U739 ( .A(n1464), .Y(n30) );
  ivd1_hd U740 ( .A(n30), .Y(n31) );
  ivd1_hd U741 ( .A(n1430), .Y(n32) );
  ivd1_hd U742 ( .A(n32), .Y(n33) );
  ivd1_hd U743 ( .A(n1462), .Y(n34) );
  ivd1_hd U744 ( .A(n34), .Y(n35) );
  ivd1_hd U745 ( .A(n1434), .Y(n36) );
  ivd1_hd U746 ( .A(n36), .Y(n37) );
  ivd1_hd U747 ( .A(n1440), .Y(n38) );
  ivd1_hd U748 ( .A(n38), .Y(n39) );
  ivd1_hd U749 ( .A(n1357), .Y(n40) );
  ivd1_hd U750 ( .A(n40), .Y(n41) );
  ivd1_hd U751 ( .A(n1361), .Y(n42) );
  ivd1_hd U752 ( .A(n42), .Y(n43) );
  ivd1_hd U753 ( .A(n1365), .Y(n44) );
  ivd1_hd U754 ( .A(n44), .Y(n45) );
  ivd1_hd U755 ( .A(n1369), .Y(n46) );
  ivd1_hd U756 ( .A(n46), .Y(n47) );
  ivd1_hd U757 ( .A(n[1555]), .Y(n48) );
  ivd1_hd U758 ( .A(n[1555]), .Y(n49) );
  ivd1_hd U759 ( .A(n704), .Y(n50) );
  ivd1_hd U760 ( .A(n50), .Y(n51) );
  ivd1_hd U761 ( .A(n701), .Y(n52) );
  ivd1_hd U762 ( .A(n701), .Y(n53) );
  ivd1_hd U763 ( .A(n515), .Y(n54) );
  ivd1_hd U764 ( .A(n515), .Y(n55) );
  ivd1_hd U765 ( .A(n1273), .Y(n56) );
  ivd1_hd U766 ( .A(n1273), .Y(n57) );
  ivd1_hd U767 ( .A(n1435), .Y(n58) );
  ivd1_hd U768 ( .A(n58), .Y(n59) );
  ivd1_hd U769 ( .A(n1352), .Y(n60) );
  ivd1_hd U770 ( .A(n60), .Y(n61) );
  ivd1_hd U771 ( .A(n1373), .Y(n62) );
  ivd1_hd U772 ( .A(n62), .Y(n63) );
  ivd1_hd U773 ( .A(n51), .Y(n64) );
  ivd1_hd U774 ( .A(n119), .Y(n65) );
  ivd1_hd U775 ( .A(n[1554]), .Y(n66) );
  ivd1_hd U776 ( .A(n[1554]), .Y(n67) );
  ivd1_hd U777 ( .A(n896), .Y(n68) );
  ivd1_hd U778 ( .A(n896), .Y(n69) );
  ivd1_hd U779 ( .A(n928), .Y(n70) );
  ivd1_hd U780 ( .A(n928), .Y(n71) );
  ivd1_hd U781 ( .A(n313), .Y(n72) );
  ivd1_hd U782 ( .A(n313), .Y(n73) );
  ivd1_hd U783 ( .A(n697), .Y(n74) );
  ivd1_hd U784 ( .A(n697), .Y(n75) );
  ivd1_hd U785 ( .A(n697), .Y(n76) );
  ivd1_hd U786 ( .A(n99), .Y(n77) );
  ivd1_hd U787 ( .A(n100), .Y(n78) );
  ivd1_hd U788 ( .A(n1006), .Y(n79) );
  ivd1_hd U789 ( .A(n557), .Y(n80) );
  ivd1_hd U790 ( .A(n557), .Y(n81) );
  ivd1_hd U791 ( .A(n557), .Y(n82) );
  ivd1_hd U792 ( .A(n557), .Y(n83) );
  ivd1_hd U793 ( .A(n556), .Y(n84) );
  ivd1_hd U794 ( .A(n84), .Y(n85) );
  ivd1_hd U795 ( .A(n84), .Y(n86) );
  ivd1_hd U796 ( .A(n84), .Y(n87) );
  ivd1_hd U797 ( .A(n926), .Y(n88) );
  ivd1_hd U798 ( .A(n926), .Y(n89) );
  nid1_hd U799 ( .A(n307), .Y(n90) );
  nid1_hd U800 ( .A(n887), .Y(n91) );
  nid1_hd U801 ( .A(n1449), .Y(n92) );
  nid1_hd U802 ( .A(n1447), .Y(n94) );
  ivd1_hd U803 ( .A(n765), .Y(n95) );
  nid1_hd U804 ( .A(n1444), .Y(n96) );
  ivd1_hd U805 ( .A(n13), .Y(n97) );
  nid1_hd U806 ( .A(n692), .Y(n98) );
  xo2d1_hd U807 ( .A(n988), .B(n100), .Y(n1058) );
  xo2d1_hd U808 ( .A(n1005), .B(n99), .Y(n1063) );
  xo2d1_hd U809 ( .A(n979), .B(n145), .Y(n1064) );
  xo2d1_hd U810 ( .A(n1007), .B(n100), .Y(n1066) );
  xo2d1_hd U811 ( .A(n964), .B(n99), .Y(n1068) );
  xo2d1_hd U812 ( .A(n959), .B(n145), .Y(n1070) );
  xo2d1_hd U813 ( .A(n955), .B(n100), .Y(n1071) );
  xo2d1_hd U814 ( .A(n960), .B(n99), .Y(n1073) );
  xo2d1_hd U815 ( .A(n971), .B(n145), .Y(n1074) );
  xo2d1_hd U816 ( .A(n972), .B(n100), .Y(n1077) );
  xo2d1_hd U817 ( .A(n983), .B(n99), .Y(n1079) );
  xo2d1_hd U818 ( .A(n987), .B(n145), .Y(n1081) );
  xo2d1_hd U819 ( .A(n1001), .B(n100), .Y(n1082) );
  ivd1_hd U820 ( .A(n548), .Y(n101) );
  ivd1_hd U821 ( .A(n548), .Y(n102) );
  ivd1_hd U822 ( .A(n548), .Y(n105) );
  ivd1_hd U823 ( .A(n548), .Y(n109) );
  ivd1_hd U824 ( .A(n52), .Y(n113) );
  ivd1_hd U825 ( .A(n52), .Y(n114) );
  ivd1_hd U826 ( .A(n52), .Y(n115) );
  ivd1_hd U827 ( .A(n846), .Y(n116) );
  ad2d1_hd U828 ( .A(n51), .B(n68), .Y(n685) );
  ivd1_hd U829 ( .A(n685), .Y(n117) );
  ivd1_hd U830 ( .A(n685), .Y(n118) );
  ivd1_hd U831 ( .A(n685), .Y(n119) );
  or2d1_hd U832 ( .A(n48), .B(n510), .Y(n1017) );
  ivd1_hd U833 ( .A(n1017), .Y(n120) );
  ivd1_hd U834 ( .A(n1017), .Y(n121) );
  ivd1_hd U835 ( .A(n1017), .Y(n122) );
  ivd1_hd U836 ( .A(n170), .Y(n162) );
  ivd1_hd U837 ( .A(n169), .Y(n168) );
  ivd1_hd U838 ( .A(n169), .Y(n166) );
  ivd1_hd U839 ( .A(n172), .Y(n160) );
  ivd1_hd U840 ( .A(n169), .Y(n167) );
  nr2d1_hd U841 ( .A(n1273), .B(n196), .Y(n885) );
  scg20d1_hd U842 ( .A(n1273), .B(n534), .C(n827), .Y(n1014) );
  nd2bd1_hd U843 ( .AN(n1257), .B(n568), .Y(n704) );
  scg6d1_hd U844 ( .A(n520), .B(n524), .C(n189), .Y(n123) );
  ivd1_hd U845 ( .A(n193), .Y(n189) );
  ivd1_hd U846 ( .A(n867), .Y(n887) );
  nr2bd1_hd U847 ( .AN(n530), .B(n527), .Y(n870) );
  ivd1_hd U848 ( .A(n74), .Y(n692) );
  ivd1_hd U849 ( .A(n120), .Y(n1028) );
  ivd1_hd U850 ( .A(n558), .Y(n508) );
  ivd1_hd U851 ( .A(n151), .Y(n147) );
  ivd1_hd U852 ( .A(n135), .Y(n133) );
  ivd1_hd U853 ( .A(n135), .Y(n126) );
  ivd1_hd U854 ( .A(n135), .Y(n131) );
  ivd1_hd U855 ( .A(n123), .Y(n148) );
  ivd1_hd U856 ( .A(n191), .Y(n181) );
  ivd1_hd U857 ( .A(n151), .Y(n146) );
  ivd1_hd U858 ( .A(n151), .Y(n149) );
  ivd1_hd U859 ( .A(n824), .Y(n827) );
  ivd1_hd U860 ( .A(n894), .Y(n932) );
  ivd1_hd U861 ( .A(n931), .Y(n930) );
  nr2d1_hd U862 ( .A(n66), .B(n564), .Y(n931) );
  ivd1_hd U863 ( .A(n564), .Y(n889) );
  nr2d1_hd U864 ( .A(n313), .B(n280), .Y(n306) );
  ivd1_hd U865 ( .A(n301), .Y(n280) );
  ivd1_hd U866 ( .A(n358), .Y(n334) );
  ivd1_hd U867 ( .A(n830), .Y(n547) );
  ivd1_hd U868 ( .A(n1441), .Y(n992) );
  ivd1_hd U869 ( .A(n1478), .Y(n993) );
  ivd1_hd U870 ( .A(n191), .Y(n185) );
  ivd1_hd U871 ( .A(n737), .Y(n125) );
  ivd1_hd U872 ( .A(n192), .Y(n188) );
  ivd1_hd U873 ( .A(n192), .Y(n187) );
  ivd1_hd U874 ( .A(n192), .Y(n186) );
  ivd1_hd U875 ( .A(n192), .Y(n183) );
  ivd1_hd U876 ( .A(n192), .Y(n182) );
  ivd1_hd U877 ( .A(n191), .Y(n184) );
  ivd1_hd U878 ( .A(n885), .Y(n846) );
  nr2d1_hd U879 ( .A(n1413), .B(n930), .Y(n705) );
  ivd1_hd U880 ( .A(n1371), .Y(n594) );
  ivd1_hd U881 ( .A(n1367), .Y(n617) );
  ivd1_hd U882 ( .A(n1385), .Y(n902) );
  ivd1_hd U883 ( .A(n[1557]), .Y(n1275) );
  ivd1_hd U884 ( .A(n306), .Y(n765) );
  oa21d1_hd U885 ( .A(n256), .B(n511), .C(n150), .Y(n301) );
  ivd1_hd U886 ( .A(n191), .Y(n190) );
  oa21d1_hd U887 ( .A(n312), .B(n511), .C(n134), .Y(n358) );
  ivd1_hd U888 ( .A(n1485), .Y(n914) );
  ivd1_hd U889 ( .A(n1487), .Y(n906) );
  ivd1_hd U890 ( .A(n1446), .Y(n343) );
  ivd1_hd U891 ( .A(n1484), .Y(n916) );
  ivd1_hd U892 ( .A(n1482), .Y(n912) );
  ivd1_hd U893 ( .A(n1483), .Y(n910) );
  ivd1_hd U894 ( .A(n1480), .Y(n302) );
  nr2d1_hd U895 ( .A(n312), .B(n528), .Y(n530) );
  ivd1_hd U896 ( .A(n1443), .Y(n359) );
  ivd1_hd U897 ( .A(n1477), .Y(n937) );
  ivd1_hd U898 ( .A(n1438), .Y(n1002) );
  ivd1_hd U899 ( .A(n1429), .Y(n968) );
  ivd1_hd U900 ( .A(n1426), .Y(n956) );
  ivd1_hd U901 ( .A(n1455), .Y(n990) );
  ivd1_hd U902 ( .A(n1454), .Y(n945) );
  ivd1_hd U903 ( .A(n1418), .Y(n989) );
  ivd1_hd U904 ( .A(n1423), .Y(n995) );
  ivd1_hd U905 ( .A(n1422), .Y(n984) );
  ivd1_hd U906 ( .A(n1431), .Y(n965) );
  ivd1_hd U907 ( .A(n1436), .Y(n976) );
  ivd1_hd U908 ( .A(n1437), .Y(n980) );
  ivd1_hd U909 ( .A(n1475), .Y(n1003) );
  ivd1_hd U910 ( .A(n1476), .Y(n974) );
  ivd1_hd U911 ( .A(n1415), .Y(n821) );
  nd3d1_hd U912 ( .A(n1271), .B(i_AB_STB), .C(o_AB_ACK), .Y(n1272) );
  nr2d1_hd U913 ( .A(n[1557]), .B(n920), .Y(n1271) );
  ivd1_hd U914 ( .A(n888), .Y(n843) );
  ivd1_hd U915 ( .A(n1353), .Y(n698) );
  ivd1_hd U916 ( .A(n1375), .Y(n711) );
  ivd1_hd U917 ( .A(n1350), .Y(n936) );
  ivd1_hd U918 ( .A(n1372), .Y(n588) );
  ivd1_hd U919 ( .A(n1368), .Y(n605) );
  ivd1_hd U920 ( .A(n1363), .Y(n641) );
  ivd1_hd U921 ( .A(n1364), .Y(n628) );
  ivd1_hd U922 ( .A(n1359), .Y(n665) );
  ivd1_hd U923 ( .A(n1360), .Y(n652) );
  ivd1_hd U924 ( .A(n1355), .Y(n690) );
  ivd1_hd U925 ( .A(n1356), .Y(n676) );
  ivd1_hd U926 ( .A(n1374), .Y(n891) );
  nr2bd1_hd U927 ( .AN(n1377), .B(n929), .Y(n858) );
  ivd1_hd U928 ( .A(n1376), .Y(n929) );
  scg17d1_hd U929 ( .A(n1488), .B(n768), .C(n767), .D(n766), .Y(n1136) );
  scg17d1_hd U930 ( .A(n1451), .B(n925), .C(n924), .D(n923), .Y(n1126) );
  ivd1_hd U931 ( .A(n1552), .Y(n260) );
  nr2d1_hd U932 ( .A(n254), .B(n313), .Y(n520) );
  ivd1_hd U933 ( .A(n1520), .Y(n317) );
  ao22d1_hd U934 ( .A(n1489), .B(n518), .C(n243), .D(n242), .Y(n254) );
  ivd1_hd U935 ( .A(n1481), .Y(n908) );
  ivd1_hd U936 ( .A(n1450), .Y(n922) );
  ivd1_hd U937 ( .A(n1486), .Y(n919) );
  ivd1_hd U938 ( .A(n1452), .Y(n518) );
  nr2d1_hd U939 ( .A(n530), .B(n527), .Y(n534) );
  nr2d1_hd U940 ( .A(n256), .B(n529), .Y(n830) );
  nr4d1_hd U941 ( .A(n1451), .B(n1452), .C(n222), .D(n221), .Y(n549) );
  ivd1_hd U942 ( .A(n1488), .Y(n904) );
  ivd1_hd U943 ( .A(n1489), .Y(n308) );
  ivd1_hd U944 ( .A(n1448), .Y(n328) );
  nr2d1_hd U945 ( .A(n[1557]), .B(n67), .Y(n253) );
  nr2d1_hd U946 ( .A(n[1556]), .B(n48), .Y(n244) );
  ivd1_hd U947 ( .A(n1416), .Y(n941) );
  ivd1_hd U948 ( .A(n1417), .Y(n946) );
  ivd1_hd U949 ( .A(n1421), .Y(n943) );
  ivd1_hd U950 ( .A(n1424), .Y(n939) );
  ivd1_hd U951 ( .A(n1466), .Y(n969) );
  ivd1_hd U952 ( .A(n1468), .Y(n966) );
  ivd1_hd U953 ( .A(n1467), .Y(n951) );
  ivd1_hd U954 ( .A(n1428), .Y(n954) );
  ivd1_hd U955 ( .A(n1459), .Y(n985) );
  ivd1_hd U956 ( .A(n1458), .Y(n942) );
  ivd1_hd U957 ( .A(n1457), .Y(n962) );
  ivd1_hd U958 ( .A(n1420), .Y(n961) );
  ivd1_hd U959 ( .A(n1453), .Y(n940) );
  ivd1_hd U960 ( .A(n1419), .Y(n944) );
  ivd1_hd U961 ( .A(n1460), .Y(n996) );
  ivd1_hd U962 ( .A(n1461), .Y(n938) );
  ivd1_hd U963 ( .A(n1425), .Y(n952) );
  ivd1_hd U964 ( .A(n1463), .Y(n957) );
  ivd1_hd U965 ( .A(n1427), .Y(n949) );
  ivd1_hd U966 ( .A(n1465), .Y(n953) );
  ivd1_hd U967 ( .A(n1470), .Y(n1009) );
  ivd1_hd U968 ( .A(n1433), .Y(n1008) );
  ivd1_hd U969 ( .A(n1432), .Y(n947) );
  ivd1_hd U970 ( .A(n1471), .Y(n948) );
  ivd1_hd U971 ( .A(n1472), .Y(n950) );
  ivd1_hd U972 ( .A(n1473), .Y(n977) );
  ivd1_hd U973 ( .A(n1474), .Y(n981) );
  ivd1_hd U974 ( .A(n1442), .Y(n999) );
  ivd1_hd U975 ( .A(n1414), .Y(n822) );
  nd4d1_hd U976 ( .A(n49), .B(n1274), .C(n[1554]), .D(n[1557]), .Y(n824) );
  ivd1_hd U977 ( .A(n[1556]), .Y(n1274) );
  nr2d1_hd U978 ( .A(n[1555]), .B(n[1556]), .Y(n509) );
  nr2d1_hd U979 ( .A(n1442), .B(n998), .Y(n818) );
  ao22d1_hd U980 ( .A(n1441), .B(n993), .C(n1442), .D(n998), .Y(n820) );
  oa22d1_hd U981 ( .A(n822), .B(n821), .C(n1415), .D(n1414), .Y(n1006) );
  nr2d1_hd U982 ( .A(n549), .B(n547), .Y(n869) );
  oa21d1_hd U983 ( .A(n1383), .B(n1384), .C(n902), .Y(n823) );
  nd2bd1_hd U984 ( .AN(n252), .B(n251), .Y(n524) );
  ivd1_hd U985 ( .A(n151), .Y(n150) );
  ivd1_hd U986 ( .A(n135), .Y(n134) );
  nd4d1_hd U987 ( .A(n1487), .B(n910), .C(n912), .D(n916), .Y(n207) );
  nr4d1_hd U988 ( .A(n1486), .B(n1481), .C(n1485), .D(n207), .Y(n219) );
  nd4d1_hd U989 ( .A(n1480), .B(n219), .C(n1489), .D(n1488), .Y(n256) );
  nr2d1_hd U990 ( .A(n1446), .B(n359), .Y(n210) );
  ivd1_hd U991 ( .A(n1444), .Y(n310) );
  ivd1_hd U992 ( .A(n1449), .Y(n831) );
  ivd1_hd U993 ( .A(n1445), .Y(n837) );
  ivd1_hd U994 ( .A(n1447), .Y(n845) );
  nd4d1_hd U995 ( .A(n310), .B(n831), .C(n837), .D(n845), .Y(n208) );
  nr2d1_hd U996 ( .A(n209), .B(n208), .Y(n220) );
  nd4d1_hd U997 ( .A(n1451), .B(n1452), .C(n210), .D(n220), .Y(n312) );
  nr4d1_hd U998 ( .A(n1439), .B(n1438), .C(n39), .D(n1441), .Y(n218) );
  nr4d1_hd U999 ( .A(n1435), .B(n1434), .C(n1437), .D(n1436), .Y(n217) );
  nr4d1_hd U1000 ( .A(n1428), .B(n1431), .C(n1430), .D(n1432), .Y(n216) );
  nr4d1_hd U1001 ( .A(n1417), .B(n1416), .C(n1418), .D(n1433), .Y(n211) );
  nd3d1_hd U1002 ( .A(n211), .B(n944), .C(n961), .Y(n214) );
  nd4d1_hd U1003 ( .A(n949), .B(n956), .C(n939), .D(n968), .Y(n213) );
  nd4d1_hd U1004 ( .A(n943), .B(n984), .C(n995), .D(n952), .Y(n212) );
  nr4d1_hd U1005 ( .A(n1442), .B(n214), .C(n213), .D(n212), .Y(n215) );
  nd4d1_hd U1006 ( .A(n218), .B(n217), .C(n216), .D(n215), .Y(n528) );
  ivd1_hd U1007 ( .A(n220), .Y(n222) );
  nr2d1_hd U1008 ( .A(n550), .B(n549), .Y(n825) );
  nd3d1_hd U1009 ( .A(n974), .B(n1003), .C(n993), .Y(n230) );
  nr4d1_hd U1010 ( .A(n1455), .B(n1456), .C(n1457), .D(n1458), .Y(n223) );
  nd4d1_hd U1011 ( .A(n223), .B(n945), .C(n940), .D(n998), .Y(n229) );
  nr4d1_hd U1012 ( .A(n1463), .B(n1464), .C(n1466), .D(n1465), .Y(n227) );
  nr4d1_hd U1013 ( .A(n1459), .B(n1460), .C(n35), .D(n1461), .Y(n226) );
  nr4d1_hd U1014 ( .A(n1472), .B(n1470), .C(n1471), .D(n1473), .Y(n225) );
  nr4d1_hd U1015 ( .A(n1468), .B(n1467), .C(n27), .D(n1474), .Y(n224) );
  nd4d1_hd U1016 ( .A(n227), .B(n226), .C(n225), .D(n224), .Y(n228) );
  ivd1_hd U1017 ( .A(n1451), .Y(n514) );
  ao22d1_hd U1018 ( .A(n1488), .B(n514), .C(n1452), .D(n308), .Y(n243) );
  ao22d1_hd U1019 ( .A(n1451), .B(n904), .C(n1450), .D(n906), .Y(n247) );
  ao211d1_hd U1020 ( .A(n1444), .B(n908), .C(n1443), .D(n302), .Y(n232) );
  oa22d1_hd U1021 ( .A(n1444), .B(n908), .C(n1445), .D(n912), .Y(n231) );
  nr2d1_hd U1022 ( .A(n232), .B(n231), .Y(n234) );
  ao22d1_hd U1023 ( .A(n912), .B(n1445), .C(n910), .D(n1446), .Y(n248) );
  ivd1_hd U1024 ( .A(n248), .Y(n233) );
  oa22d1_hd U1025 ( .A(n1447), .B(n916), .C(n234), .D(n233), .Y(n235) );
  ao21d1_hd U1026 ( .A(n1483), .B(n343), .C(n235), .Y(n238) );
  oa22d1_hd U1027 ( .A(n1448), .B(n914), .C(n238), .D(n252), .Y(n239) );
  ao22d1_hd U1028 ( .A(n1487), .B(n922), .C(n246), .D(n239), .Y(n240) );
  oa21d1_hd U1029 ( .A(n919), .B(n1449), .C(n240), .Y(n241) );
  nr2d1_hd U1030 ( .A(n1452), .B(n308), .Y(n250) );
  nd4d1_hd U1031 ( .A(n248), .B(n247), .C(n246), .D(n245), .Y(n249) );
  ao211d1_hd U1032 ( .A(n1443), .B(n302), .C(n250), .D(n249), .Y(n251) );
  scg16d1_hd U1033 ( .A(n256), .B(n511), .C(n149), .Y(n1277) );
  scg16d1_hd U1034 ( .A(n312), .B(n511), .C(n133), .Y(n1276) );
  nr2d1_hd U1035 ( .A(n302), .B(n908), .Y(n255) );
  nr2d1_hd U1036 ( .A(n910), .B(n286), .Y(n277) );
  nr2d1_hd U1037 ( .A(n914), .B(n272), .Y(n262) );
  ao21d1_hd U1038 ( .A(n72), .B(n764), .C(n280), .Y(n305) );
  nr2d1_hd U1039 ( .A(n193), .B(n260), .Y(n258) );
  ivd1_hd U1040 ( .A(n292), .Y(n289) );
  ivd1_hd U1041 ( .A(n1549), .Y(n279) );
  nr2d1_hd U1042 ( .A(n288), .B(n279), .Y(n278) );
  ivd1_hd U1043 ( .A(n1551), .Y(n263) );
  nr2d1_hd U1044 ( .A(n274), .B(n263), .Y(n259) );
  nr2d1_hd U1045 ( .A(n765), .B(n764), .Y(n257) );
  ao22d1_hd U1046 ( .A(n258), .B(n259), .C(n257), .D(n906), .Y(n261) );
  nr2d1_hd U1047 ( .A(n259), .B(n192), .Y(n267) );
  oa211d1_hd U1048 ( .A(n305), .B(n906), .C(n261), .D(n766), .Y(n1135) );
  ao21d1_hd U1049 ( .A(n73), .B(n272), .C(n280), .Y(n273) );
  ao22d1_hd U1050 ( .A(n1486), .B(n268), .C(n267), .D(n264), .Y(n269) );
  oa211d1_hd U1051 ( .A(n1486), .B(n270), .C(n269), .D(n307), .Y(n1134) );
  oa22d1_hd U1052 ( .A(n273), .B(n914), .C(n272), .D(n271), .Y(n276) );
  oa211d1_hd U1053 ( .A(n278), .B(n1550), .C(n190), .D(n274), .Y(n275) );
  nd3bd1_hd U1054 ( .AN(n276), .B(n90), .C(n275), .Y(n1133) );
  ao211d1_hd U1055 ( .A(n288), .B(n279), .C(n278), .D(n191), .Y(n282) );
  ao21d1_hd U1056 ( .A(n73), .B(n286), .C(n280), .Y(n287) );
  ao21d1_hd U1057 ( .A(n287), .B(n285), .C(n916), .Y(n281) );
  nr2d1_hd U1058 ( .A(n282), .B(n281), .Y(n283) );
  oa211d1_hd U1059 ( .A(n1484), .B(n284), .C(n283), .D(n307), .Y(n1132) );
  oa22d1_hd U1060 ( .A(n287), .B(n910), .C(n286), .D(n285), .Y(n291) );
  oa211d1_hd U1061 ( .A(n289), .B(n1548), .C(n190), .D(n288), .Y(n290) );
  nd3bd1_hd U1062 ( .AN(n291), .B(n90), .C(n290), .Y(n1131) );
  nr2d1_hd U1063 ( .A(n1481), .B(n765), .Y(n297) );
  oa21d1_hd U1064 ( .A(n297), .B(n296), .C(n1482), .Y(n295) );
  nd4d1_hd U1065 ( .A(n1481), .B(n1480), .C(n95), .D(n912), .Y(n294) );
  oa211d1_hd U1066 ( .A(n300), .B(n1547), .C(n190), .D(n292), .Y(n293) );
  nd4d1_hd U1067 ( .A(n90), .B(n295), .C(n294), .D(n293), .Y(n1130) );
  oa21d1_hd U1068 ( .A(n1546), .B(n1545), .C(n190), .Y(n299) );
  ao22d1_hd U1069 ( .A(n1480), .B(n297), .C(n1481), .D(n296), .Y(n298) );
  oa211d1_hd U1070 ( .A(n300), .B(n299), .C(n298), .D(n307), .Y(n1129) );
  oa21d1_hd U1071 ( .A(n1487), .B(n765), .C(n305), .Y(n768) );
  ao21d1_hd U1072 ( .A(n95), .B(n904), .C(n768), .Y(n309) );
  oa211d1_hd U1073 ( .A(n309), .B(n308), .C(n766), .D(n90), .Y(n1127) );
  nr2d1_hd U1074 ( .A(n310), .B(n359), .Y(n311) );
  nr2d1_hd U1075 ( .A(n343), .B(n342), .Y(n333) );
  nr2d1_hd U1076 ( .A(n328), .B(n327), .Y(n319) );
  ao21d1_hd U1077 ( .A(n73), .B(n921), .C(n334), .Y(n513) );
  nr2d1_hd U1078 ( .A(n193), .B(n317), .Y(n315) );
  ivd1_hd U1079 ( .A(n349), .Y(n346) );
  ivd1_hd U1080 ( .A(n1517), .Y(n336) );
  nr2d1_hd U1081 ( .A(n345), .B(n336), .Y(n335) );
  ivd1_hd U1082 ( .A(n1519), .Y(n320) );
  nr2d1_hd U1083 ( .A(n330), .B(n320), .Y(n316) );
  nr2d1_hd U1084 ( .A(n515), .B(n921), .Y(n314) );
  ao22d1_hd U1085 ( .A(n315), .B(n316), .C(n314), .D(n922), .Y(n318) );
  nr2d1_hd U1086 ( .A(n316), .B(n193), .Y(n322) );
  oa211d1_hd U1087 ( .A(n513), .B(n922), .C(n318), .D(n923), .Y(n1125) );
  ao21d1_hd U1088 ( .A(n72), .B(n327), .C(n334), .Y(n329) );
  ao22d1_hd U1089 ( .A(n92), .B(n323), .C(n322), .D(n321), .Y(n324) );
  oa211d1_hd U1090 ( .A(n92), .B(n325), .C(n324), .D(n22), .Y(n1124) );
  oa22d1_hd U1091 ( .A(n329), .B(n328), .C(n327), .D(n326), .Y(n332) );
  oa211d1_hd U1092 ( .A(n335), .B(n1518), .C(n190), .D(n330), .Y(n331) );
  nd3bd1_hd U1093 ( .AN(n332), .B(n23), .C(n331), .Y(n1123) );
  ao21d1_hd U1094 ( .A(n72), .B(n342), .C(n334), .Y(n344) );
  ao211d1_hd U1095 ( .A(n345), .B(n336), .C(n335), .D(n191), .Y(n337) );
  ao21d1_hd U1096 ( .A(n338), .B(n94), .C(n337), .Y(n339) );
  oa211d1_hd U1097 ( .A(n94), .B(n340), .C(n339), .D(n23), .Y(n1122) );
  oa22d1_hd U1098 ( .A(n344), .B(n343), .C(n342), .D(n341), .Y(n348) );
  oa211d1_hd U1099 ( .A(n346), .B(n1516), .C(n189), .D(n345), .Y(n347) );
  nd3bd1_hd U1100 ( .AN(n348), .B(n22), .C(n347), .Y(n1121) );
  nr2d1_hd U1101 ( .A(n96), .B(n515), .Y(n353) );
  oa21d1_hd U1102 ( .A(n353), .B(n354), .C(n1445), .Y(n352) );
  nd4d1_hd U1103 ( .A(n96), .B(n1443), .C(n55), .D(n837), .Y(n351) );
  oa211d1_hd U1104 ( .A(n357), .B(n1515), .C(n189), .D(n349), .Y(n350) );
  nd4d1_hd U1105 ( .A(n22), .B(n352), .C(n351), .D(n350), .Y(n1120) );
  oa21d1_hd U1106 ( .A(n1514), .B(n1513), .C(n190), .Y(n356) );
  ao22d1_hd U1107 ( .A(n96), .B(n354), .C(n1443), .D(n353), .Y(n355) );
  oa211d1_hd U1108 ( .A(n357), .B(n356), .C(n355), .D(n22), .Y(n1119) );
  nr3d1_hd U1109 ( .A(n73), .B(n121), .C(n889), .Y(n1270) );
  ao22d1_hd U1110 ( .A(n1441), .B(n125), .C(n188), .D(n1512), .Y(n512) );
  oa21d1_hd U1111 ( .A(n999), .B(n137), .C(n512), .Y(n1113) );
  oa21d1_hd U1112 ( .A(n1450), .B(n515), .C(n513), .Y(n925) );
  ao21d1_hd U1113 ( .A(n54), .B(n514), .C(n925), .Y(n519) );
  oa211d1_hd U1114 ( .A(n519), .B(n518), .C(n923), .D(n23), .Y(n1112) );
  ivd1_hd U1115 ( .A(n520), .Y(n523) );
  nr4d1_hd U1116 ( .A(n1381), .B(n1382), .C(n1380), .D(n1378), .Y(n521) );
  nd2bd1_hd U1117 ( .AN(n1379), .B(n521), .Y(n560) );
  nr2d1_hd U1118 ( .A(n560), .B(n858), .Y(n522) );
  oa21d1_hd U1119 ( .A(n559), .B(n522), .C(n1385), .Y(n562) );
  oa22d1_hd U1120 ( .A(n524), .B(n523), .C(n1028), .D(n562), .Y(n1262) );
  scg12d1_hd U1121 ( .A(n1273), .B(n525), .C(n827), .Y(n1266) );
  nr2d1_hd U1122 ( .A(n201), .B(o_Z_STB), .Y(n1258) );
  ao22d1_hd U1123 ( .A(n550), .B(n529), .C(n549), .D(n528), .Y(n551) );
  ao21d1_hd U1124 ( .A(n530), .B(n821), .C(n547), .Y(n531) );
  oa21d1_hd U1125 ( .A(n549), .B(n531), .C(n1414), .Y(n532) );
  oa211d1_hd U1126 ( .A(n549), .B(n533), .C(n551), .D(n532), .Y(n535) );
  ao22d1_hd U1127 ( .A(n57), .B(n535), .C(n195), .D(n1347), .Y(n546) );
  ivd1_hd U1128 ( .A(n1354), .Y(n683) );
  nd4d1_hd U1129 ( .A(n683), .B(n676), .C(n690), .D(n40), .Y(n536) );
  nr4d1_hd U1130 ( .A(n63), .B(n61), .C(n1353), .D(n536), .Y(n542) );
  ivd1_hd U1131 ( .A(n1366), .Y(n611) );
  nd4d1_hd U1132 ( .A(n42), .B(n628), .C(n641), .D(n611), .Y(n540) );
  ivd1_hd U1133 ( .A(n1358), .Y(n658) );
  ivd1_hd U1134 ( .A(n1362), .Y(n634) );
  nd4d1_hd U1135 ( .A(n658), .B(n652), .C(n665), .D(n634), .Y(n539) );
  nd4d1_hd U1136 ( .A(n891), .B(n46), .C(n588), .D(n594), .Y(n538) );
  ivd1_hd U1137 ( .A(n1370), .Y(n582) );
  nd4d1_hd U1138 ( .A(n44), .B(n605), .C(n617), .D(n582), .Y(n537) );
  nr4d1_hd U1139 ( .A(n540), .B(n539), .C(n538), .D(n537), .Y(n541) );
  nr4d1_hd U1140 ( .A(n1376), .B(n560), .C(n902), .D(n559), .Y(n543) );
  nd3d1_hd U1141 ( .A(n1377), .B(n543), .C(n711), .Y(n826) );
  oa211d1_hd U1142 ( .A(n544), .B(n826), .C(n827), .D(n1348), .Y(n545) );
  oa211d1_hd U1143 ( .A(n548), .B(n821), .C(n546), .D(n545), .Y(n1255) );
  ao22d1_hd U1144 ( .A(n1478), .B(n105), .C(n1374), .D(n85), .Y(n555) );
  nd3d1_hd U1145 ( .A(n550), .B(n549), .C(n77), .Y(n552) );
  ao22d1_hd U1146 ( .A(n195), .B(n1338), .C(n885), .D(n553), .Y(n554) );
  oa211d1_hd U1147 ( .A(n992), .B(n844), .C(n555), .D(n554), .Y(n1246) );
  scg4d1_hd U1148 ( .A(n1440), .B(n80), .C(n199), .D(n1337), .E(n1373), .F(n86), .G(n101), .H(n1477), .Y(n1245) );
  scg4d1_hd U1149 ( .A(n1476), .B(n105), .C(n1014), .D(n1336), .E(n1372), .F(
        n556), .G(n1439), .H(n82), .Y(n1244) );
  scg4d1_hd U1150 ( .A(n1475), .B(n109), .C(n1014), .D(n1335), .E(n1371), .F(
        n85), .G(n1438), .H(n83), .Y(n1243) );
  scg4d1_hd U1151 ( .A(n1474), .B(n101), .C(n1014), .D(n1334), .E(n1370), .F(
        n86), .G(n1437), .H(n80), .Y(n1242) );
  scg4d1_hd U1152 ( .A(n1473), .B(n102), .C(n1014), .D(n1333), .E(n47), .F(n87), .G(n1436), .H(n81), .Y(n1241) );
  scg4d1_hd U1153 ( .A(n1472), .B(n105), .C(n197), .D(n1332), .E(n1368), .F(
        n556), .G(n59), .H(n82), .Y(n1240) );
  scg4d1_hd U1154 ( .A(n1471), .B(n109), .C(n198), .D(n1331), .E(n1367), .F(
        n85), .G(n1434), .H(n83), .Y(n1239) );
  scg4d1_hd U1155 ( .A(n1433), .B(n81), .C(n198), .D(n1330), .E(n1366), .F(n87), .G(n102), .H(n1470), .Y(n1238) );
  scg4d1_hd U1156 ( .A(n1469), .B(n101), .C(n198), .D(n1329), .E(n45), .F(n86), 
        .G(n1432), .H(n80), .Y(n1237) );
  scg4d1_hd U1157 ( .A(n1468), .B(n102), .C(n198), .D(n1328), .E(n1364), .F(
        n87), .G(n1431), .H(n81), .Y(n1236) );
  scg4d1_hd U1158 ( .A(n1467), .B(n105), .C(n198), .D(n1327), .E(n1363), .F(
        n556), .G(n1430), .H(n82), .Y(n1235) );
  scg4d1_hd U1159 ( .A(n1466), .B(n109), .C(n198), .D(n1326), .E(n1362), .F(
        n85), .G(n1429), .H(n83), .Y(n1234) );
  scg4d1_hd U1160 ( .A(n1465), .B(n101), .C(n197), .D(n1325), .E(n43), .F(n86), 
        .G(n1428), .H(n80), .Y(n1233) );
  scg4d1_hd U1161 ( .A(n1427), .B(n82), .C(n197), .D(n1324), .E(n1360), .F(
        n556), .G(n105), .H(n1464), .Y(n1232) );
  scg4d1_hd U1162 ( .A(n1463), .B(n102), .C(n197), .D(n1323), .E(n1359), .F(
        n87), .G(n1426), .H(n81), .Y(n1231) );
  scg4d1_hd U1163 ( .A(n1462), .B(n105), .C(n197), .D(n1322), .E(n1358), .F(
        n556), .G(n1425), .H(n82), .Y(n1230) );
  scg4d1_hd U1164 ( .A(n1461), .B(n109), .C(n197), .D(n1321), .E(n41), .F(n85), 
        .G(n1424), .H(n83), .Y(n1229) );
  scg4d1_hd U1165 ( .A(n1423), .B(n83), .C(n199), .D(n1320), .E(n1356), .F(n85), .G(n109), .H(n1460), .Y(n1228) );
  scg4d1_hd U1166 ( .A(n1459), .B(n101), .C(n194), .D(n1319), .E(n1355), .F(
        n86), .G(n1422), .H(n80), .Y(n1227) );
  scg4d1_hd U1167 ( .A(n1421), .B(n80), .C(n194), .D(n1318), .E(n1354), .F(n86), .G(n101), .H(n1458), .Y(n1226) );
  scg4d1_hd U1168 ( .A(n1457), .B(n102), .C(n194), .D(n1317), .E(n1353), .F(
        n87), .G(n1420), .H(n81), .Y(n1225) );
  scg4d1_hd U1169 ( .A(n1419), .B(n81), .C(n194), .D(n1316), .E(n1352), .F(n87), .G(n102), .H(n1456), .Y(n1224) );
  scg20d1_hd U1170 ( .A(n1377), .B(n560), .C(n559), .Y(n561) );
  nr2d1_hd U1171 ( .A(n561), .B(n902), .Y(n1286) );
  nr2d1_hd U1172 ( .A(n1375), .B(n1028), .Y(n563) );
  ao22d1_hd U1173 ( .A(n20), .B(n1286), .C(n563), .D(n562), .Y(n895) );
  ao22d1_hd U1174 ( .A(n140), .B(n1387), .C(n156), .D(n1388), .Y(n566) );
  nd3d1_hd U1175 ( .A(n20), .B(n1351), .C(n1257), .Y(n565) );
  oa211d1_hd U1176 ( .A(n936), .B(n1257), .C(n566), .D(n565), .Y(n1222) );
  oa211d1_hd U1177 ( .A(n1349), .B(n567), .C(n1351), .D(n68), .Y(n568) );
  ao22d1_hd U1178 ( .A(n140), .B(n1411), .C(n159), .D(n1412), .Y(n572) );
  nd3d1_hd U1179 ( .A(n61), .B(n1353), .C(n1354), .Y(n671) );
  nr3d1_hd U1180 ( .A(n671), .B(n676), .C(n690), .Y(n660) );
  nd3d1_hd U1181 ( .A(n660), .B(n41), .C(n1358), .Y(n647) );
  nr3d1_hd U1182 ( .A(n647), .B(n652), .C(n665), .Y(n635) );
  nd3d1_hd U1183 ( .A(n635), .B(n1362), .C(n43), .Y(n623) );
  nr3d1_hd U1184 ( .A(n623), .B(n628), .C(n641), .Y(n612) );
  nd3d1_hd U1185 ( .A(n612), .B(n1366), .C(n45), .Y(n600) );
  nr3d1_hd U1186 ( .A(n600), .B(n605), .C(n617), .Y(n589) );
  nd3d1_hd U1187 ( .A(n589), .B(n1370), .C(n47), .Y(n577) );
  nr3d1_hd U1188 ( .A(n577), .B(n588), .C(n594), .Y(n569) );
  oa21d1_hd U1189 ( .A(n1374), .B(n708), .C(n113), .Y(n570) );
  ivd1_hd U1190 ( .A(n569), .Y(n890) );
  oa21d1_hd U1191 ( .A(n64), .B(n890), .C(n659), .Y(n573) );
  oa21d1_hd U1192 ( .A(n1373), .B(n119), .C(n573), .Y(n706) );
  ao22d1_hd U1193 ( .A(n63), .B(n570), .C(n1374), .D(n706), .Y(n571) );
  oa211d1_hd U1194 ( .A(n711), .B(n75), .C(n572), .D(n571), .Y(n1221) );
  ao22d1_hd U1195 ( .A(n140), .B(n1410), .C(n1411), .D(n156), .Y(n576) );
  ao22d1_hd U1196 ( .A(n63), .B(n573), .C(n708), .D(n62), .Y(n574) );
  ao21d1_hd U1197 ( .A(n53), .B(n1372), .C(n574), .Y(n575) );
  oa211d1_hd U1198 ( .A(n891), .B(n74), .C(n576), .D(n575), .Y(n1220) );
  nr2d1_hd U1199 ( .A(n577), .B(n117), .Y(n585) );
  ao21d1_hd U1200 ( .A(n585), .B(n588), .C(n52), .Y(n581) );
  ao22d1_hd U1201 ( .A(n140), .B(n1409), .C(n932), .D(n1410), .Y(n580) );
  ao21d1_hd U1202 ( .A(n68), .B(n577), .C(n64), .Y(n583) );
  oa21d1_hd U1203 ( .A(n1371), .B(n117), .C(n583), .Y(n578) );
  ao22d1_hd U1204 ( .A(n1373), .B(n98), .C(n1372), .D(n578), .Y(n579) );
  oa211d1_hd U1205 ( .A(n581), .B(n594), .C(n580), .D(n579), .Y(n1219) );
  ao22d1_hd U1206 ( .A(n140), .B(n1408), .C(n159), .D(n1409), .Y(n587) );
  oa22d1_hd U1207 ( .A(n583), .B(n594), .C(n114), .D(n582), .Y(n584) );
  ao21d1_hd U1208 ( .A(n585), .B(n594), .C(n584), .Y(n586) );
  oa211d1_hd U1209 ( .A(n588), .B(n76), .C(n587), .D(n586), .Y(n1218) );
  ao22d1_hd U1210 ( .A(n140), .B(n1407), .C(n932), .D(n1408), .Y(n593) );
  scg14d1_hd U1211 ( .A(n51), .B(n589), .C(n659), .Y(n596) );
  oa21d1_hd U1212 ( .A(n47), .B(n118), .C(n596), .Y(n591) );
  oa21d1_hd U1213 ( .A(n1370), .B(n595), .C(n115), .Y(n590) );
  ao22d1_hd U1214 ( .A(n1370), .B(n591), .C(n47), .D(n590), .Y(n592) );
  oa211d1_hd U1215 ( .A(n594), .B(n75), .C(n593), .D(n592), .Y(n1217) );
  ao22d1_hd U1216 ( .A(n705), .B(n1406), .C(n932), .D(n1407), .Y(n599) );
  ao22d1_hd U1217 ( .A(n47), .B(n596), .C(n595), .D(n46), .Y(n597) );
  ao21d1_hd U1218 ( .A(n1370), .B(n98), .C(n597), .Y(n598) );
  oa211d1_hd U1219 ( .A(n114), .B(n605), .C(n599), .D(n598), .Y(n1216) );
  nr2d1_hd U1220 ( .A(n600), .B(n118), .Y(n608) );
  ao21d1_hd U1221 ( .A(n608), .B(n605), .C(n52), .Y(n604) );
  ao22d1_hd U1222 ( .A(n143), .B(n1405), .C(n932), .D(n1406), .Y(n603) );
  ao21d1_hd U1223 ( .A(n68), .B(n600), .C(n64), .Y(n606) );
  oa21d1_hd U1224 ( .A(n1367), .B(n118), .C(n606), .Y(n601) );
  ao22d1_hd U1225 ( .A(n1368), .B(n601), .C(n1369), .D(n692), .Y(n602) );
  oa211d1_hd U1226 ( .A(n604), .B(n617), .C(n603), .D(n602), .Y(n1215) );
  ao22d1_hd U1227 ( .A(n143), .B(n1404), .C(n159), .D(n1405), .Y(n610) );
  oa22d1_hd U1228 ( .A(n606), .B(n617), .C(n605), .D(n75), .Y(n607) );
  ao21d1_hd U1229 ( .A(n608), .B(n617), .C(n607), .Y(n609) );
  oa211d1_hd U1230 ( .A(n113), .B(n611), .C(n610), .D(n609), .Y(n1214) );
  ao22d1_hd U1231 ( .A(n143), .B(n1403), .C(n158), .D(n1404), .Y(n616) );
  scg14d1_hd U1232 ( .A(n51), .B(n612), .C(n659), .Y(n619) );
  oa21d1_hd U1233 ( .A(n45), .B(n119), .C(n619), .Y(n614) );
  oa21d1_hd U1234 ( .A(n1366), .B(n618), .C(n114), .Y(n613) );
  ao22d1_hd U1235 ( .A(n1366), .B(n614), .C(n45), .D(n613), .Y(n615) );
  oa211d1_hd U1236 ( .A(n617), .B(n74), .C(n616), .D(n615), .Y(n1213) );
  ao22d1_hd U1237 ( .A(n705), .B(n1402), .C(n158), .D(n1403), .Y(n622) );
  ao22d1_hd U1238 ( .A(n45), .B(n619), .C(n618), .D(n44), .Y(n620) );
  ao21d1_hd U1239 ( .A(n1366), .B(n98), .C(n620), .Y(n621) );
  oa211d1_hd U1240 ( .A(n115), .B(n628), .C(n622), .D(n621), .Y(n1212) );
  nr2d1_hd U1241 ( .A(n623), .B(n119), .Y(n631) );
  ao21d1_hd U1242 ( .A(n631), .B(n628), .C(n53), .Y(n627) );
  ao22d1_hd U1243 ( .A(n143), .B(n1401), .C(n158), .D(n1402), .Y(n626) );
  ao21d1_hd U1244 ( .A(n69), .B(n623), .C(n64), .Y(n629) );
  oa21d1_hd U1245 ( .A(n1363), .B(n119), .C(n629), .Y(n624) );
  ao22d1_hd U1246 ( .A(n1364), .B(n624), .C(n1365), .D(n692), .Y(n625) );
  oa211d1_hd U1247 ( .A(n627), .B(n641), .C(n626), .D(n625), .Y(n1211) );
  ao22d1_hd U1248 ( .A(n141), .B(n1400), .C(n159), .D(n1401), .Y(n633) );
  oa22d1_hd U1249 ( .A(n629), .B(n641), .C(n628), .D(n76), .Y(n630) );
  ao21d1_hd U1250 ( .A(n631), .B(n641), .C(n630), .Y(n632) );
  oa211d1_hd U1251 ( .A(n114), .B(n634), .C(n633), .D(n632), .Y(n1210) );
  ao22d1_hd U1252 ( .A(n141), .B(n1399), .C(n157), .D(n1400), .Y(n640) );
  scg14d1_hd U1253 ( .A(n704), .B(n635), .C(n659), .Y(n643) );
  oa21d1_hd U1254 ( .A(n43), .B(n117), .C(n643), .Y(n638) );
  oa21d1_hd U1255 ( .A(n1362), .B(n642), .C(n113), .Y(n637) );
  ao22d1_hd U1256 ( .A(n1362), .B(n638), .C(n43), .D(n637), .Y(n639) );
  oa211d1_hd U1257 ( .A(n641), .B(n76), .C(n640), .D(n639), .Y(n1209) );
  ao22d1_hd U1258 ( .A(n141), .B(n1398), .C(n157), .D(n1399), .Y(n646) );
  ao22d1_hd U1259 ( .A(n43), .B(n643), .C(n642), .D(n42), .Y(n644) );
  ao21d1_hd U1260 ( .A(n1362), .B(n98), .C(n644), .Y(n645) );
  oa211d1_hd U1261 ( .A(n113), .B(n652), .C(n646), .D(n645), .Y(n1208) );
  nr2d1_hd U1262 ( .A(n647), .B(n117), .Y(n655) );
  ao21d1_hd U1263 ( .A(n655), .B(n652), .C(n52), .Y(n651) );
  ao22d1_hd U1264 ( .A(n141), .B(n1397), .C(n157), .D(n1398), .Y(n650) );
  ao21d1_hd U1265 ( .A(n68), .B(n647), .C(n50), .Y(n653) );
  oa21d1_hd U1266 ( .A(n1359), .B(n117), .C(n653), .Y(n648) );
  ao22d1_hd U1267 ( .A(n1360), .B(n648), .C(n1361), .D(n692), .Y(n649) );
  oa211d1_hd U1268 ( .A(n651), .B(n665), .C(n650), .D(n649), .Y(n1207) );
  ao22d1_hd U1269 ( .A(n141), .B(n1396), .C(n157), .D(n1397), .Y(n657) );
  oa22d1_hd U1270 ( .A(n653), .B(n665), .C(n652), .D(n76), .Y(n654) );
  ao21d1_hd U1271 ( .A(n655), .B(n665), .C(n654), .Y(n656) );
  oa211d1_hd U1272 ( .A(n115), .B(n658), .C(n657), .D(n656), .Y(n1206) );
  ao22d1_hd U1273 ( .A(n141), .B(n1395), .C(n157), .D(n1396), .Y(n664) );
  oa21d1_hd U1274 ( .A(n1358), .B(n666), .C(n115), .Y(n662) );
  scg14d1_hd U1275 ( .A(n704), .B(n660), .C(n659), .Y(n667) );
  oa21d1_hd U1276 ( .A(n41), .B(n119), .C(n667), .Y(n661) );
  ao22d1_hd U1277 ( .A(n1357), .B(n662), .C(n1358), .D(n661), .Y(n663) );
  oa211d1_hd U1278 ( .A(n665), .B(n75), .C(n664), .D(n663), .Y(n1205) );
  ao22d1_hd U1279 ( .A(n142), .B(n1394), .C(n157), .D(n1395), .Y(n670) );
  ao22d1_hd U1280 ( .A(n41), .B(n667), .C(n666), .D(n40), .Y(n668) );
  ao21d1_hd U1281 ( .A(n1358), .B(n98), .C(n668), .Y(n669) );
  oa211d1_hd U1282 ( .A(n114), .B(n676), .C(n670), .D(n669), .Y(n1204) );
  nr2d1_hd U1283 ( .A(n671), .B(n118), .Y(n680) );
  ao21d1_hd U1284 ( .A(n680), .B(n676), .C(n53), .Y(n675) );
  ao22d1_hd U1285 ( .A(n142), .B(n1393), .C(n158), .D(n1394), .Y(n674) );
  ao21d1_hd U1286 ( .A(n69), .B(n671), .C(n64), .Y(n678) );
  oa21d1_hd U1287 ( .A(n1355), .B(n118), .C(n678), .Y(n672) );
  ao22d1_hd U1288 ( .A(n1356), .B(n672), .C(n41), .D(n692), .Y(n673) );
  oa211d1_hd U1289 ( .A(n675), .B(n690), .C(n674), .D(n673), .Y(n1203) );
  ao22d1_hd U1290 ( .A(n142), .B(n1392), .C(n156), .D(n1393), .Y(n682) );
  oa22d1_hd U1291 ( .A(n678), .B(n690), .C(n676), .D(n74), .Y(n679) );
  ao21d1_hd U1292 ( .A(n680), .B(n690), .C(n679), .Y(n681) );
  oa211d1_hd U1293 ( .A(n113), .B(n683), .C(n682), .D(n681), .Y(n1202) );
  ao22d1_hd U1294 ( .A(n142), .B(n1391), .C(n156), .D(n1392), .Y(n689) );
  oa21d1_hd U1295 ( .A(n1354), .B(n684), .C(n114), .Y(n687) );
  nr2d1_hd U1296 ( .A(n61), .B(n118), .Y(n700) );
  nr2d1_hd U1297 ( .A(n50), .B(n700), .Y(n696) );
  ao22d1_hd U1298 ( .A(n1353), .B(n687), .C(n1354), .D(n686), .Y(n688) );
  oa211d1_hd U1299 ( .A(n690), .B(n74), .C(n689), .D(n688), .Y(n1201) );
  ao22d1_hd U1300 ( .A(n142), .B(n1390), .C(n156), .D(n1391), .Y(n695) );
  ao22d1_hd U1301 ( .A(n61), .B(n693), .C(n1354), .D(n692), .Y(n694) );
  oa211d1_hd U1302 ( .A(n696), .B(n698), .C(n695), .D(n694), .Y(n1200) );
  ao22d1_hd U1303 ( .A(n142), .B(n1389), .C(n156), .D(n1390), .Y(n703) );
  nr2d1_hd U1304 ( .A(n698), .B(n75), .Y(n699) );
  ao211d1_hd U1305 ( .A(n53), .B(n1351), .C(n700), .D(n699), .Y(n702) );
  oa211d1_hd U1306 ( .A(n60), .B(n704), .C(n703), .D(n702), .Y(n1199) );
  scg4d1_hd U1307 ( .A(n120), .B(n1350), .C(n20), .D(n1352), .E(n143), .F(
        n1388), .G(n1389), .H(n158), .Y(n1256) );
  ao21d1_hd U1308 ( .A(n65), .B(n891), .C(n706), .Y(n712) );
  oa21d1_hd U1309 ( .A(n708), .B(n707), .C(n113), .Y(n709) );
  ao22d1_hd U1310 ( .A(n931), .B(n1412), .C(n1374), .D(n709), .Y(n710) );
  oa211d1_hd U1311 ( .A(n712), .B(n711), .C(n710), .D(n894), .Y(n1198) );
  ao22d1_hd U1312 ( .A(n39), .B(n125), .C(n188), .D(n1511), .Y(n713) );
  oa21d1_hd U1313 ( .A(n992), .B(n137), .C(n713), .Y(n1187) );
  ao22d1_hd U1314 ( .A(n1439), .B(n125), .C(n188), .D(n1510), .Y(n714) );
  oa21d1_hd U1315 ( .A(n38), .B(n137), .C(n714), .Y(n1186) );
  ao22d1_hd U1316 ( .A(n1438), .B(n125), .C(n188), .D(n1509), .Y(n715) );
  oa21d1_hd U1317 ( .A(n973), .B(n137), .C(n715), .Y(n1185) );
  ao22d1_hd U1318 ( .A(n1437), .B(n126), .C(n188), .D(n1508), .Y(n716) );
  oa21d1_hd U1319 ( .A(n1002), .B(n137), .C(n716), .Y(n1184) );
  ao22d1_hd U1320 ( .A(n1436), .B(n125), .C(n187), .D(n1507), .Y(n717) );
  oa21d1_hd U1321 ( .A(n980), .B(n137), .C(n717), .Y(n1183) );
  ao22d1_hd U1322 ( .A(n1435), .B(n126), .C(n188), .D(n1506), .Y(n719) );
  oa21d1_hd U1323 ( .A(n976), .B(n139), .C(n719), .Y(n1182) );
  ao22d1_hd U1324 ( .A(n37), .B(n126), .C(n187), .D(n1505), .Y(n720) );
  oa21d1_hd U1325 ( .A(n58), .B(n144), .C(n720), .Y(n1181) );
  ao22d1_hd U1326 ( .A(n1433), .B(n126), .C(n187), .D(n1504), .Y(n722) );
  oa21d1_hd U1327 ( .A(n36), .B(n144), .C(n722), .Y(n1180) );
  ao22d1_hd U1328 ( .A(n1432), .B(n126), .C(n187), .D(n1503), .Y(n723) );
  oa21d1_hd U1329 ( .A(n1008), .B(n139), .C(n723), .Y(n1179) );
  ao22d1_hd U1330 ( .A(n1431), .B(n126), .C(n187), .D(n1502), .Y(n724) );
  oa21d1_hd U1331 ( .A(n947), .B(n139), .C(n724), .Y(n1178) );
  ao22d1_hd U1332 ( .A(n1430), .B(n131), .C(n186), .D(n1501), .Y(n725) );
  oa21d1_hd U1333 ( .A(n965), .B(n139), .C(n725), .Y(n1177) );
  ao22d1_hd U1334 ( .A(n1429), .B(n131), .C(n187), .D(n1500), .Y(n726) );
  oa21d1_hd U1335 ( .A(n32), .B(n144), .C(n726), .Y(n1176) );
  ao22d1_hd U1336 ( .A(n1428), .B(n131), .C(n186), .D(n1499), .Y(n727) );
  oa21d1_hd U1337 ( .A(n968), .B(n739), .C(n727), .Y(n1175) );
  ao22d1_hd U1338 ( .A(n1427), .B(n131), .C(n186), .D(n1498), .Y(n729) );
  oa21d1_hd U1339 ( .A(n954), .B(n739), .C(n729), .Y(n1174) );
  ao22d1_hd U1340 ( .A(n1426), .B(n131), .C(n186), .D(n1497), .Y(n730) );
  oa21d1_hd U1341 ( .A(n949), .B(n739), .C(n730), .Y(n1173) );
  ao22d1_hd U1342 ( .A(n1425), .B(n131), .C(n186), .D(n1496), .Y(n731) );
  oa21d1_hd U1343 ( .A(n956), .B(n739), .C(n731), .Y(n1172) );
  ao22d1_hd U1344 ( .A(n1424), .B(n133), .C(n186), .D(n1495), .Y(n732) );
  oa21d1_hd U1345 ( .A(n952), .B(n739), .C(n732), .Y(n1171) );
  ao22d1_hd U1346 ( .A(n1423), .B(n133), .C(n185), .D(n1494), .Y(n733) );
  oa21d1_hd U1347 ( .A(n939), .B(n138), .C(n733), .Y(n1170) );
  ao22d1_hd U1348 ( .A(n1422), .B(n133), .C(n185), .D(n1493), .Y(n734) );
  oa21d1_hd U1349 ( .A(n995), .B(n138), .C(n734), .Y(n1169) );
  ao22d1_hd U1350 ( .A(n1421), .B(n133), .C(n185), .D(n1492), .Y(n735) );
  oa21d1_hd U1351 ( .A(n984), .B(n138), .C(n735), .Y(n1168) );
  ao22d1_hd U1352 ( .A(n1420), .B(n133), .C(n185), .D(n1491), .Y(n736) );
  oa21d1_hd U1353 ( .A(n943), .B(n138), .C(n736), .Y(n1167) );
  ao22d1_hd U1354 ( .A(n1419), .B(n125), .C(n185), .D(n1490), .Y(n738) );
  oa21d1_hd U1355 ( .A(n961), .B(n138), .C(n738), .Y(n1166) );
  oa22d1_hd U1356 ( .A(n989), .B(n737), .C(n944), .D(n138), .Y(n1165) );
  oa22d1_hd U1357 ( .A(n946), .B(n737), .C(n989), .D(n139), .Y(n1164) );
  oa22d1_hd U1358 ( .A(n189), .B(n941), .C(n946), .D(n139), .Y(n1163) );
  ao22d1_hd U1359 ( .A(n1477), .B(n149), .C(n184), .D(n1543), .Y(n740) );
  oa21d1_hd U1360 ( .A(n993), .B(n153), .C(n740), .Y(n1162) );
  ao22d1_hd U1361 ( .A(n1476), .B(n149), .C(n184), .D(n1542), .Y(n741) );
  oa21d1_hd U1362 ( .A(n937), .B(n155), .C(n741), .Y(n1161) );
  ao22d1_hd U1363 ( .A(n1475), .B(n149), .C(n184), .D(n1541), .Y(n742) );
  oa21d1_hd U1364 ( .A(n974), .B(n155), .C(n742), .Y(n1160) );
  ao22d1_hd U1365 ( .A(n1474), .B(n149), .C(n184), .D(n1540), .Y(n743) );
  oa21d1_hd U1366 ( .A(n1003), .B(n155), .C(n743), .Y(n1159) );
  ao22d1_hd U1367 ( .A(n1473), .B(n149), .C(n184), .D(n1539), .Y(n744) );
  oa21d1_hd U1368 ( .A(n981), .B(n155), .C(n744), .Y(n1158) );
  ao22d1_hd U1369 ( .A(n1472), .B(n148), .C(n184), .D(n1538), .Y(n745) );
  oa21d1_hd U1370 ( .A(n977), .B(n155), .C(n745), .Y(n1157) );
  ao22d1_hd U1371 ( .A(n1471), .B(n148), .C(n183), .D(n1537), .Y(n746) );
  oa21d1_hd U1372 ( .A(n950), .B(n152), .C(n746), .Y(n1156) );
  ao22d1_hd U1373 ( .A(n1470), .B(n148), .C(n183), .D(n1536), .Y(n747) );
  oa21d1_hd U1374 ( .A(n948), .B(n763), .C(n747), .Y(n1155) );
  ao22d1_hd U1375 ( .A(n27), .B(n148), .C(n185), .D(n1535), .Y(n748) );
  oa21d1_hd U1376 ( .A(n1009), .B(n763), .C(n748), .Y(n1154) );
  ao22d1_hd U1377 ( .A(n1468), .B(n148), .C(n183), .D(n1534), .Y(n749) );
  oa21d1_hd U1378 ( .A(n26), .B(n152), .C(n749), .Y(n1153) );
  ao22d1_hd U1379 ( .A(n1467), .B(n147), .C(n183), .D(n1533), .Y(n750) );
  oa21d1_hd U1380 ( .A(n966), .B(n763), .C(n750), .Y(n1152) );
  ao22d1_hd U1381 ( .A(n1466), .B(n147), .C(n183), .D(n1532), .Y(n751) );
  oa21d1_hd U1382 ( .A(n951), .B(n763), .C(n751), .Y(n1151) );
  ao22d1_hd U1383 ( .A(n1465), .B(n147), .C(n182), .D(n1531), .Y(n752) );
  oa21d1_hd U1384 ( .A(n969), .B(n154), .C(n752), .Y(n1150) );
  ao22d1_hd U1385 ( .A(n1464), .B(n147), .C(n182), .D(n1530), .Y(n753) );
  oa21d1_hd U1386 ( .A(n953), .B(n154), .C(n753), .Y(n1149) );
  ao22d1_hd U1387 ( .A(n1463), .B(n147), .C(n182), .D(n1529), .Y(n754) );
  oa21d1_hd U1388 ( .A(n30), .B(n154), .C(n754), .Y(n1148) );
  ao22d1_hd U1389 ( .A(n35), .B(n147), .C(n182), .D(n1528), .Y(n755) );
  oa21d1_hd U1390 ( .A(n957), .B(n154), .C(n755), .Y(n1147) );
  ao22d1_hd U1391 ( .A(n1461), .B(n146), .C(n182), .D(n1527), .Y(n756) );
  oa21d1_hd U1392 ( .A(n34), .B(n154), .C(n756), .Y(n1146) );
  ao22d1_hd U1393 ( .A(n1460), .B(n146), .C(n182), .D(n1526), .Y(n757) );
  oa21d1_hd U1394 ( .A(n938), .B(n153), .C(n757), .Y(n1145) );
  ao22d1_hd U1395 ( .A(n1459), .B(n146), .C(n181), .D(n1525), .Y(n758) );
  oa21d1_hd U1396 ( .A(n996), .B(n153), .C(n758), .Y(n1144) );
  ao22d1_hd U1397 ( .A(n1458), .B(n146), .C(n181), .D(n1524), .Y(n759) );
  oa21d1_hd U1398 ( .A(n985), .B(n153), .C(n759), .Y(n1143) );
  ao22d1_hd U1399 ( .A(n1457), .B(n146), .C(n183), .D(n1523), .Y(n760) );
  oa21d1_hd U1400 ( .A(n942), .B(n153), .C(n760), .Y(n1142) );
  ao22d1_hd U1401 ( .A(n1456), .B(n146), .C(n181), .D(n1522), .Y(n761) );
  oa21d1_hd U1402 ( .A(n962), .B(n153), .C(n761), .Y(n1141) );
  oa22d1_hd U1403 ( .A(n990), .B(n123), .C(n24), .D(n155), .Y(n1140) );
  oa22d1_hd U1404 ( .A(n945), .B(n151), .C(n990), .D(n152), .Y(n1139) );
  oa22d1_hd U1405 ( .A(n189), .B(n940), .C(n945), .D(n152), .Y(n1138) );
  ao22d1_hd U1406 ( .A(n1478), .B(n148), .C(n181), .D(n1544), .Y(n762) );
  oa21d1_hd U1407 ( .A(n998), .B(n154), .C(n762), .Y(n1137) );
  nr4d1_hd U1408 ( .A(n1488), .B(n906), .C(n765), .D(n764), .Y(n767) );
  ao211d1_hd U1409 ( .A(n1439), .B(n974), .C(n1438), .D(n1003), .Y(n814) );
  nr2d1_hd U1410 ( .A(n1473), .B(n976), .Y(n808) );
  ao211d1_hd U1411 ( .A(n59), .B(n950), .C(n1434), .D(n948), .Y(n773) );
  ao22d1_hd U1412 ( .A(n27), .B(n947), .C(n1470), .D(n1008), .Y(n771) );
  ao22d1_hd U1413 ( .A(n1433), .B(n1009), .C(n37), .D(n948), .Y(n770) );
  oa22d1_hd U1414 ( .A(n59), .B(n950), .C(n771), .D(n804), .Y(n772) );
  nr2d1_hd U1415 ( .A(n773), .B(n772), .Y(n774) );
  oa22d1_hd U1416 ( .A(n1436), .B(n977), .C(n808), .D(n774), .Y(n775) );
  ao22d1_hd U1417 ( .A(n1474), .B(n980), .C(n776), .D(n775), .Y(n811) );
  nr2d1_hd U1418 ( .A(n1468), .B(n965), .Y(n777) );
  nr2d1_hd U1419 ( .A(n777), .B(n33), .Y(n778) );
  ao22d1_hd U1420 ( .A(n1468), .B(n965), .C(n1467), .D(n778), .Y(n806) );
  ao211d1_hd U1421 ( .A(n1427), .B(n30), .C(n1426), .D(n957), .Y(n796) );
  nr2d1_hd U1422 ( .A(n35), .B(n952), .Y(n791) );
  nr2d1_hd U1423 ( .A(n791), .B(n1424), .Y(n779) );
  ao22d1_hd U1424 ( .A(n35), .B(n952), .C(n1461), .D(n779), .Y(n794) );
  ao22d1_hd U1425 ( .A(n1459), .B(n984), .C(n1460), .D(n995), .Y(n789) );
  ao22d1_hd U1426 ( .A(n1455), .B(n989), .C(n25), .D(n944), .Y(n784) );
  ao22d1_hd U1427 ( .A(n1417), .B(n945), .C(n1418), .D(n990), .Y(n781) );
  oa211d1_hd U1428 ( .A(n1417), .B(n945), .C(n1416), .D(n940), .Y(n780) );
  oa22d1_hd U1429 ( .A(n25), .B(n944), .C(n1457), .D(n961), .Y(n782) );
  ao21d1_hd U1430 ( .A(n784), .B(n783), .C(n782), .Y(n787) );
  oa22d1_hd U1431 ( .A(n1420), .B(n962), .C(n1421), .D(n942), .Y(n786) );
  ao22d1_hd U1432 ( .A(n1421), .B(n942), .C(n1422), .D(n985), .Y(n785) );
  oa21d1_hd U1433 ( .A(n787), .B(n786), .C(n785), .Y(n788) );
  ao22d1_hd U1434 ( .A(n1423), .B(n996), .C(n789), .D(n788), .Y(n790) );
  scg17d1_hd U1435 ( .A(n938), .B(n1424), .C(n791), .D(n790), .Y(n793) );
  oa22d1_hd U1436 ( .A(n1463), .B(n956), .C(n31), .D(n949), .Y(n792) );
  ao21d1_hd U1437 ( .A(n794), .B(n793), .C(n792), .Y(n795) );
  ao211d1_hd U1438 ( .A(n31), .B(n949), .C(n796), .D(n795), .Y(n797) );
  nr2d1_hd U1439 ( .A(n1466), .B(n968), .Y(n798) );
  ao211d1_hd U1440 ( .A(n1428), .B(n953), .C(n797), .D(n798), .Y(n802) );
  nr2d1_hd U1441 ( .A(n953), .B(n798), .Y(n799) );
  ao22d1_hd U1442 ( .A(n33), .B(n951), .C(n1431), .D(n966), .Y(n800) );
  oa21d1_hd U1443 ( .A(n802), .B(n801), .C(n800), .Y(n805) );
  oa22d1_hd U1444 ( .A(n1474), .B(n980), .C(n27), .D(n947), .Y(n803) );
  ao211d1_hd U1445 ( .A(n806), .B(n805), .C(n804), .D(n803), .Y(n807) );
  nd2bd1_hd U1446 ( .AN(n808), .B(n807), .Y(n810) );
  oa22d1_hd U1447 ( .A(n1475), .B(n1002), .C(n1476), .D(n973), .Y(n809) );
  ao21d1_hd U1448 ( .A(n811), .B(n810), .C(n809), .Y(n813) );
  ao22d1_hd U1449 ( .A(n169), .B(n822), .C(n821), .D(n160), .Y(n1287) );
  oa22d1_hd U1450 ( .A(n825), .B(n846), .C(n824), .D(n823), .Y(n867) );
  nr2d1_hd U1451 ( .A(n1377), .B(n1376), .Y(n859) );
  ivd1_hd U1452 ( .A(n1378), .Y(n835) );
  nr2d1_hd U1453 ( .A(n1379), .B(n877), .Y(n876) );
  ivd1_hd U1454 ( .A(n1380), .Y(n841) );
  nr2d1_hd U1455 ( .A(n1381), .B(n851), .Y(n850) );
  ivd1_hd U1456 ( .A(n1382), .Y(n828) );
  oa21d1_hd U1457 ( .A(n850), .B(n828), .C(n866), .Y(n829) );
  ao22d1_hd U1458 ( .A(n196), .B(n1345), .C(n843), .D(n829), .Y(n834) );
  nr2d1_hd U1459 ( .A(n1485), .B(n1448), .Y(n854) );
  ao22d1_hd U1460 ( .A(n1480), .B(n870), .C(n1443), .D(n830), .Y(n884) );
  nr2d1_hd U1461 ( .A(n1481), .B(n96), .Y(n861) );
  nr3d1_hd U1462 ( .A(n1482), .B(n1445), .C(n860), .Y(n880) );
  nr2d1_hd U1463 ( .A(n1483), .B(n1446), .Y(n879) );
  nr3d1_hd U1464 ( .A(n1484), .B(n94), .C(n878), .Y(n853) );
  nr3d1_hd U1465 ( .A(n1486), .B(n92), .C(n852), .Y(n872) );
  oa22d1_hd U1466 ( .A(n919), .B(n846), .C(n831), .D(n844), .Y(n832) );
  ao22d1_hd U1467 ( .A(n116), .B(n872), .C(n852), .D(n832), .Y(n833) );
  nd3d1_hd U1468 ( .A(n91), .B(n834), .C(n833), .Y(n1253) );
  oa21d1_hd U1469 ( .A(n859), .B(n835), .C(n877), .Y(n836) );
  ao22d1_hd U1470 ( .A(n196), .B(n1341), .C(n843), .D(n836), .Y(n840) );
  oa22d1_hd U1471 ( .A(n912), .B(n846), .C(n837), .D(n844), .Y(n838) );
  ao22d1_hd U1472 ( .A(n116), .B(n880), .C(n860), .D(n838), .Y(n839) );
  nd3d1_hd U1473 ( .A(n91), .B(n840), .C(n839), .Y(n1249) );
  oa21d1_hd U1474 ( .A(n876), .B(n841), .C(n851), .Y(n842) );
  ao22d1_hd U1475 ( .A(n196), .B(n1343), .C(n843), .D(n842), .Y(n849) );
  oa22d1_hd U1476 ( .A(n916), .B(n846), .C(n845), .D(n844), .Y(n847) );
  ao22d1_hd U1477 ( .A(n116), .B(n853), .C(n878), .D(n847), .Y(n848) );
  nd3d1_hd U1478 ( .A(n91), .B(n849), .C(n848), .Y(n1251) );
  ao21d1_hd U1479 ( .A(n1381), .B(n851), .C(n850), .Y(n857) );
  oa21d1_hd U1480 ( .A(n854), .B(n853), .C(n852), .Y(n855) );
  ao22d1_hd U1481 ( .A(n195), .B(n1344), .C(n885), .D(n855), .Y(n856) );
  oa211d1_hd U1482 ( .A(n857), .B(n888), .C(n887), .D(n856), .Y(n1252) );
  nr2d1_hd U1483 ( .A(n859), .B(n858), .Y(n864) );
  oa21d1_hd U1484 ( .A(n884), .B(n861), .C(n860), .Y(n862) );
  ao22d1_hd U1485 ( .A(n196), .B(n1340), .C(n885), .D(n862), .Y(n863) );
  oa211d1_hd U1486 ( .A(n864), .B(n888), .C(n887), .D(n863), .Y(n1248) );
  nr2d1_hd U1487 ( .A(n1383), .B(n866), .Y(n865) );
  ao211d1_hd U1488 ( .A(n1383), .B(n866), .C(n888), .D(n865), .Y(n868) );
  ao211d1_hd U1489 ( .A(n195), .B(n1346), .C(n868), .D(n867), .Y(n875) );
  ao22d1_hd U1490 ( .A(n1487), .B(n870), .C(n1450), .D(n869), .Y(n873) );
  oa211d1_hd U1491 ( .A(n873), .B(n872), .C(n116), .D(n871), .Y(n874) );
  ao21d1_hd U1492 ( .A(n1379), .B(n877), .C(n876), .Y(n883) );
  oa21d1_hd U1493 ( .A(n880), .B(n879), .C(n878), .Y(n881) );
  ao22d1_hd U1494 ( .A(n195), .B(n1342), .C(n885), .D(n881), .Y(n882) );
  oa211d1_hd U1495 ( .A(n883), .B(n888), .C(n887), .D(n882), .Y(n1250) );
  ao22d1_hd U1496 ( .A(n195), .B(n1339), .C(n116), .D(n884), .Y(n886) );
  oa211d1_hd U1497 ( .A(n1376), .B(n888), .C(n91), .D(n886), .Y(n1247) );
  nr4d1_hd U1498 ( .A(n62), .B(n896), .C(n891), .D(n890), .Y(n892) );
  nd3d1_hd U1499 ( .A(n1375), .B(n1351), .C(n892), .Y(n893) );
  nd4d1_hd U1500 ( .A(n895), .B(n918), .C(n894), .D(n893), .Y(n928) );
  ao22d1_hd U1501 ( .A(n1385), .B(n122), .C(n1028), .D(n902), .Y(n899) );
  nr2d1_hd U1502 ( .A(n122), .B(n931), .Y(n897) );
  nr2d1_hd U1503 ( .A(n21), .B(n69), .Y(n1013) );
  oa211d1_hd U1504 ( .A(n1020), .B(n899), .C(n89), .D(n898), .Y(n901) );
  oa211d1_hd U1505 ( .A(n928), .B(n902), .C(n901), .D(n900), .Y(n1188) );
  ao22d1_hd U1506 ( .A(n1384), .B(n71), .C(n88), .D(n1278), .Y(n903) );
  oa21d1_hd U1507 ( .A(n904), .B(n918), .C(n903), .Y(n1197) );
  ao22d1_hd U1508 ( .A(n1383), .B(n70), .C(n89), .D(n1279), .Y(n905) );
  oa21d1_hd U1509 ( .A(n906), .B(n918), .C(n905), .Y(n1196) );
  ao22d1_hd U1510 ( .A(n1377), .B(n71), .C(n88), .D(n1285), .Y(n907) );
  oa21d1_hd U1511 ( .A(n908), .B(n918), .C(n907), .Y(n1190) );
  ao22d1_hd U1512 ( .A(n1379), .B(n71), .C(n89), .D(n1283), .Y(n909) );
  oa21d1_hd U1513 ( .A(n910), .B(n97), .C(n909), .Y(n1192) );
  ao22d1_hd U1514 ( .A(n1378), .B(n70), .C(n89), .D(n1284), .Y(n911) );
  oa21d1_hd U1515 ( .A(n912), .B(n97), .C(n911), .Y(n1191) );
  ao22d1_hd U1516 ( .A(n1381), .B(n70), .C(n88), .D(n1281), .Y(n913) );
  oa21d1_hd U1517 ( .A(n914), .B(n97), .C(n913), .Y(n1194) );
  ao22d1_hd U1518 ( .A(n1380), .B(n71), .C(n88), .D(n1282), .Y(n915) );
  oa21d1_hd U1519 ( .A(n916), .B(n97), .C(n915), .Y(n1193) );
  ao22d1_hd U1520 ( .A(n1382), .B(n70), .C(n89), .D(n1280), .Y(n917) );
  oa21d1_hd U1521 ( .A(n919), .B(n97), .C(n917), .Y(n1195) );
  nr4d1_hd U1522 ( .A(n1451), .B(n922), .C(n515), .D(n921), .Y(n924) );
  ao22d1_hd U1523 ( .A(n1480), .B(n203), .C(n88), .D(n929), .Y(n927) );
  oa21d1_hd U1524 ( .A(n929), .B(n928), .C(n927), .Y(n1189) );
  ao22d1_hd U1525 ( .A(n931), .B(n1386), .C(n1349), .D(n930), .Y(n934) );
  oa211d1_hd U1526 ( .A(n936), .B(n935), .C(n934), .D(n933), .Y(n1223) );
  oa21d1_hd U1527 ( .A(n145), .B(n999), .C(n998), .Y(n1109) );
  ao22d1_hd U1528 ( .A(n179), .B(n992), .C(n993), .D(n160), .Y(n1108) );
  ao22d1_hd U1529 ( .A(n180), .B(n38), .C(n937), .D(n160), .Y(n1107) );
  ao22d1_hd U1530 ( .A(n179), .B(n980), .C(n981), .D(n160), .Y(n1104) );
  ao22d1_hd U1531 ( .A(n180), .B(n1002), .C(n1003), .D(n160), .Y(n1105) );
  ao22d1_hd U1532 ( .A(n171), .B(n973), .C(n974), .D(n160), .Y(n1106) );
  ao22d1_hd U1533 ( .A(n170), .B(n995), .C(n996), .D(n161), .Y(n1090) );
  ao22d1_hd U1534 ( .A(n171), .B(n939), .C(n938), .D(n161), .Y(n1091) );
  ao22d1_hd U1535 ( .A(n172), .B(n941), .C(n940), .D(n161), .Y(n1083) );
  ao22d1_hd U1536 ( .A(n178), .B(n984), .C(n985), .D(n161), .Y(n1089) );
  ao22d1_hd U1537 ( .A(n178), .B(n943), .C(n942), .D(n161), .Y(n1088) );
  ao22d1_hd U1538 ( .A(n178), .B(n961), .C(n962), .D(n161), .Y(n1087) );
  ao22d1_hd U1539 ( .A(n171), .B(n944), .C(n24), .D(n162), .Y(n1086) );
  ao22d1_hd U1540 ( .A(n172), .B(n946), .C(n945), .D(n162), .Y(n1084) );
  ao22d1_hd U1541 ( .A(n172), .B(n989), .C(n990), .D(n162), .Y(n1085) );
  ao22d1_hd U1542 ( .A(n171), .B(n1008), .C(n1009), .D(n162), .Y(n1100) );
  ao22d1_hd U1543 ( .A(n171), .B(n947), .C(n26), .D(n162), .Y(n1099) );
  ao22d1_hd U1544 ( .A(n170), .B(n976), .C(n977), .D(n162), .Y(n1103) );
  ao22d1_hd U1545 ( .A(n172), .B(n36), .C(n948), .D(n163), .Y(n1101) );
  ao22d1_hd U1546 ( .A(n170), .B(n949), .C(n30), .D(n163), .Y(n1094) );
  ao22d1_hd U1547 ( .A(n170), .B(n58), .C(n950), .D(n163), .Y(n1102) );
  ao22d1_hd U1548 ( .A(n173), .B(n965), .C(n966), .D(n163), .Y(n1098) );
  ao22d1_hd U1549 ( .A(n173), .B(n32), .C(n951), .D(n163), .Y(n1097) );
  ao22d1_hd U1550 ( .A(n173), .B(n956), .C(n957), .D(n163), .Y(n1093) );
  ao22d1_hd U1551 ( .A(n173), .B(n968), .C(n969), .D(n164), .Y(n1096) );
  ao22d1_hd U1552 ( .A(n173), .B(n952), .C(n34), .D(n164), .Y(n1092) );
  ao22d1_hd U1553 ( .A(n173), .B(n954), .C(n953), .D(n164), .Y(n1095) );
  ao22d1_hd U1554 ( .A(n174), .B(n1464), .C(n1427), .D(n164), .Y(n955) );
  ao22d1_hd U1555 ( .A(n174), .B(n957), .C(n956), .D(n164), .Y(n958) );
  ao22d1_hd U1556 ( .A(n174), .B(n1465), .C(n1428), .D(n164), .Y(n959) );
  ao22d1_hd U1557 ( .A(n174), .B(n35), .C(n1425), .D(n165), .Y(n960) );
  ao22d1_hd U1558 ( .A(n174), .B(n962), .C(n961), .D(n165), .Y(n963) );
  ao22d1_hd U1559 ( .A(n174), .B(n1467), .C(n1430), .D(n165), .Y(n964) );
  ao22d1_hd U1560 ( .A(n175), .B(n966), .C(n965), .D(n165), .Y(n967) );
  ao22d1_hd U1561 ( .A(n175), .B(n969), .C(n968), .D(n165), .Y(n970) );
  ao22d1_hd U1562 ( .A(n175), .B(n1461), .C(n1424), .D(n165), .Y(n971) );
  ao22d1_hd U1563 ( .A(n175), .B(n1458), .C(n1421), .D(n166), .Y(n972) );
  ao22d1_hd U1564 ( .A(n175), .B(n974), .C(n973), .D(n166), .Y(n975) );
  ao22d1_hd U1565 ( .A(n175), .B(n977), .C(n976), .D(n166), .Y(n978) );
  ao22d1_hd U1566 ( .A(n176), .B(n1471), .C(n37), .D(n166), .Y(n979) );
  ao22d1_hd U1567 ( .A(n176), .B(n981), .C(n980), .D(n166), .Y(n982) );
  ao22d1_hd U1568 ( .A(n176), .B(n25), .C(n1419), .D(n166), .Y(n983) );
  ao22d1_hd U1569 ( .A(n176), .B(n985), .C(n984), .D(n167), .Y(n986) );
  ao22d1_hd U1570 ( .A(n176), .B(n1454), .C(n1417), .D(n167), .Y(n987) );
  ao22d1_hd U1571 ( .A(n176), .B(n1477), .C(n1440), .D(n167), .Y(n988) );
  ao22d1_hd U1572 ( .A(n177), .B(n990), .C(n989), .D(n167), .Y(n991) );
  ao22d1_hd U1573 ( .A(n177), .B(n993), .C(n992), .D(n167), .Y(n994) );
  ao22d1_hd U1574 ( .A(n177), .B(n996), .C(n995), .D(n167), .Y(n997) );
  nr2d1_hd U1575 ( .A(n998), .B(n999), .Y(n1000) );
  ao22d1_hd U1576 ( .A(n79), .B(n1000), .C(n999), .D(n99), .Y(n1056) );
  ao22d1_hd U1577 ( .A(n177), .B(n1453), .C(n1416), .D(n168), .Y(n1001) );
  ao22d1_hd U1578 ( .A(n177), .B(n1003), .C(n1002), .D(n168), .Y(n1004) );
  ao22d1_hd U1579 ( .A(n177), .B(n1472), .C(n59), .D(n168), .Y(n1005) );
  ao22d1_hd U1580 ( .A(n1010), .B(n27), .C(n1432), .D(n168), .Y(n1007) );
  ao22d1_hd U1581 ( .A(n180), .B(n1009), .C(n1008), .D(n168), .Y(n1011) );
endmodule


module float_multiplier_1 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, 
        i_Z_ACK, i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N34, b_s, round_bit, sticky, z_s, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, C82_DATA2_1, C82_DATA2_2,
         C82_DATA2_3, C82_DATA2_4, C82_DATA2_5, C82_DATA2_6, C81_DATA2_1,
         C81_DATA2_2, C81_DATA2_3, C81_DATA2_4, C81_DATA2_5, C81_DATA2_6,
         net908, n10, n14, n36, n104, n105, n138, n141, n146, n148, n151, n155,
         n156, n157, n158, n160, n161, n171, n172, n173, n174, n177, n179,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358,
         DP_OP_116J2_127_7148_n3, DP_OP_116J2_127_7148_n4,
         DP_OP_116J2_127_7148_n5, DP_OP_116J2_127_7148_n6,
         DP_OP_116J2_127_7148_n7, DP_OP_116J2_127_7148_n8,
         DP_OP_113J2_124_6892_n3, DP_OP_113J2_124_6892_n4,
         DP_OP_113J2_124_6892_n5, DP_OP_113J2_124_6892_n6,
         DP_OP_113J2_124_6892_n7, DP_OP_113J2_124_6892_n8, C1_Z_6, C1_Z_5,
         C1_Z_4, C1_Z_3, C1_Z_2, C1_Z_1, DP_OP_125J2_130_6300_n42,
         DP_OP_125J2_130_6300_n41, DP_OP_125J2_130_6300_n40,
         DP_OP_125J2_130_6300_n39, DP_OP_125J2_130_6300_n38,
         DP_OP_125J2_130_6300_n37, DP_OP_125J2_130_6300_n36,
         DP_OP_125J2_130_6300_n35, DP_OP_125J2_130_6300_n34,
         DP_OP_125J2_130_6300_n32, DP_OP_125J2_130_6300_n31,
         DP_OP_125J2_130_6300_n30, DP_OP_125J2_130_6300_n29,
         DP_OP_125J2_130_6300_n28, DP_OP_125J2_130_6300_n27,
         DP_OP_125J2_130_6300_n26, DP_OP_125J2_130_6300_n25,
         DP_OP_125J2_130_6300_n20, DP_OP_125J2_130_6300_n19,
         DP_OP_125J2_130_6300_n18, DP_OP_125J2_130_6300_n17,
         DP_OP_125J2_130_6300_n16, DP_OP_125J2_130_6300_n15,
         DP_OP_125J2_130_6300_n14, DP_OP_125J2_130_6300_n13,
         DP_OP_125J2_130_6300_n12, DP_OP_125J2_130_6300_n9,
         DP_OP_125J2_130_6300_n8, DP_OP_125J2_130_6300_n7,
         DP_OP_125J2_130_6300_n6, DP_OP_125J2_130_6300_n5,
         DP_OP_125J2_130_6300_n4, DP_OP_125J2_130_6300_n3,
         DP_OP_125J2_130_6300_n2, n381, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1332, n1544, n1613, n1614, n1624, n1627, n1628,
         n1629, n3276, n3277, n3278, n3279, intadd_5_A_11_, intadd_5_A_10_,
         intadd_5_A_9_, intadd_5_A_8_, intadd_5_A_7_, intadd_5_A_6_,
         intadd_5_A_5_, intadd_5_A_4_, intadd_5_A_3_, intadd_5_A_2_,
         intadd_5_A_1_, intadd_5_A_0_, intadd_5_B_11_, intadd_5_B_10_,
         intadd_5_B_9_, intadd_5_B_8_, intadd_5_B_7_, intadd_5_B_6_,
         intadd_5_B_5_, intadd_5_B_4_, intadd_5_B_3_, intadd_5_B_2_,
         intadd_5_B_1_, intadd_5_B_0_, intadd_5_CI, intadd_5_SUM_11_,
         intadd_5_SUM_10_, intadd_5_SUM_9_, intadd_5_SUM_8_, intadd_5_SUM_7_,
         intadd_5_SUM_6_, intadd_5_SUM_5_, intadd_5_SUM_4_, intadd_5_SUM_3_,
         intadd_5_SUM_2_, intadd_5_SUM_1_, intadd_5_SUM_0_, intadd_5_n12,
         intadd_5_n11, intadd_5_n10, intadd_5_n9, intadd_5_n8, intadd_5_n7,
         intadd_5_n6, intadd_5_n5, intadd_5_n4, intadd_5_n3, intadd_5_n2,
         intadd_5_n1, intadd_7_A_10_, intadd_7_A_9_, intadd_7_A_8_,
         intadd_7_A_7_, intadd_7_A_6_, intadd_7_A_5_, intadd_7_A_4_,
         intadd_7_A_3_, intadd_7_A_2_, intadd_7_A_1_, intadd_7_A_0_,
         intadd_7_B_10_, intadd_7_B_9_, intadd_7_B_8_, intadd_7_B_7_,
         intadd_7_B_6_, intadd_7_B_5_, intadd_7_B_4_, intadd_7_B_3_,
         intadd_7_B_2_, intadd_7_B_1_, intadd_7_B_0_, intadd_7_CI,
         intadd_7_SUM_10_, intadd_7_SUM_9_, intadd_7_SUM_8_, intadd_7_SUM_7_,
         intadd_7_SUM_6_, intadd_7_SUM_5_, intadd_7_SUM_4_, intadd_7_SUM_3_,
         intadd_7_SUM_2_, intadd_7_SUM_1_, intadd_7_SUM_0_, intadd_7_n11,
         intadd_7_n10, intadd_7_n9, intadd_7_n8, intadd_7_n7, intadd_7_n6,
         intadd_7_n5, intadd_7_n4, intadd_7_n3, intadd_7_n2, intadd_7_n1,
         intadd_8_A_8_, intadd_8_A_7_, intadd_8_A_6_, intadd_8_A_5_,
         intadd_8_A_3_, intadd_8_A_2_, intadd_8_A_1_, intadd_8_B_8_,
         intadd_8_B_7_, intadd_8_B_6_, intadd_8_B_5_, intadd_8_B_4_,
         intadd_8_B_3_, intadd_8_B_2_, intadd_8_B_1_, intadd_8_B_0_,
         intadd_8_CI, intadd_8_SUM_8_, intadd_8_SUM_7_, intadd_8_SUM_6_,
         intadd_8_SUM_5_, intadd_8_SUM_4_, intadd_8_SUM_0_, intadd_8_n9,
         intadd_8_n8, intadd_8_n7, intadd_8_n6, intadd_8_n5, intadd_8_n4,
         intadd_8_n3, intadd_8_n2, intadd_8_n1, intadd_9_A_7_, intadd_9_A_6_,
         intadd_9_A_5_, intadd_9_A_4_, intadd_9_A_3_, intadd_9_A_2_,
         intadd_9_A_1_, intadd_9_B_7_, intadd_9_B_6_, intadd_9_B_5_,
         intadd_9_B_4_, intadd_9_B_3_, intadd_9_B_2_, intadd_9_B_1_,
         intadd_9_CI, intadd_9_SUM_7_, intadd_9_SUM_6_, intadd_9_SUM_5_,
         intadd_9_SUM_4_, intadd_9_SUM_3_, intadd_9_SUM_2_, intadd_9_SUM_1_,
         intadd_9_SUM_0_, intadd_9_n8, intadd_9_n7, intadd_9_n6, intadd_9_n5,
         intadd_9_n4, intadd_9_n3, intadd_9_n2, intadd_9_n1, intadd_10_A_5_,
         intadd_10_A_4_, intadd_10_A_3_, intadd_10_A_2_, intadd_10_A_1_,
         intadd_10_A_0_, intadd_10_B_5_, intadd_10_B_4_, intadd_10_B_3_,
         intadd_10_B_2_, intadd_10_B_1_, intadd_10_B_0_, intadd_10_CI,
         intadd_10_SUM_5_, intadd_10_SUM_4_, intadd_10_SUM_3_,
         intadd_10_SUM_2_, intadd_10_SUM_1_, intadd_10_SUM_0_, intadd_10_n6,
         intadd_10_n5, intadd_10_n4, intadd_10_n3, intadd_10_n2, intadd_10_n1,
         intadd_11_A_4_, intadd_11_A_3_, intadd_11_A_2_, intadd_11_A_1_,
         intadd_11_A_0_, intadd_11_B_4_, intadd_11_B_3_, intadd_11_B_2_,
         intadd_11_B_1_, intadd_11_B_0_, intadd_11_CI, intadd_11_SUM_4_,
         intadd_11_SUM_3_, intadd_11_SUM_2_, intadd_11_SUM_1_,
         intadd_11_SUM_0_, intadd_11_n5, intadd_11_n4, intadd_11_n3,
         intadd_11_n2, intadd_11_n1, intadd_12_A_2_, intadd_12_A_1_,
         intadd_12_B_2_, intadd_12_B_1_, intadd_12_B_0_, intadd_12_CI,
         intadd_12_n3, intadd_12_n2, intadd_12_n1, intadd_13_A_2_,
         intadd_13_A_1_, intadd_13_A_0_, intadd_13_B_2_, intadd_13_B_1_,
         intadd_13_B_0_, intadd_13_CI, intadd_13_SUM_2_, intadd_13_SUM_1_,
         intadd_13_SUM_0_, intadd_13_n3, intadd_13_n2, intadd_13_n1,
         intadd_14_A_2_, intadd_14_A_1_, intadd_14_A_0_, intadd_14_B_2_,
         intadd_14_B_1_, intadd_14_B_0_, intadd_14_CI, intadd_14_SUM_2_,
         intadd_14_SUM_1_, intadd_14_SUM_0_, intadd_14_n3, intadd_14_n2,
         intadd_14_n1, intadd_15_A_0_, intadd_15_B_2_, intadd_15_B_1_,
         intadd_15_B_0_, intadd_15_SUM_2_, intadd_15_SUM_1_, intadd_15_SUM_0_,
         intadd_15_n3, intadd_15_n2, intadd_15_n1, intadd_16_B_2_,
         intadd_16_B_1_, intadd_16_B_0_, intadd_16_CI, intadd_16_SUM_2_,
         intadd_16_SUM_1_, intadd_16_SUM_0_, intadd_16_n3, intadd_16_n2,
         intadd_16_n1, intadd_17_A_2_, intadd_17_A_1_, intadd_17_A_0_,
         intadd_17_B_2_, intadd_17_B_1_, intadd_17_B_0_, intadd_17_CI,
         intadd_17_SUM_2_, intadd_17_SUM_1_, intadd_17_SUM_0_, intadd_17_n3,
         intadd_17_n2, intadd_17_n1, intadd_18_B_2_, intadd_18_B_1_,
         intadd_18_B_0_, intadd_18_CI, intadd_18_SUM_2_, intadd_18_SUM_1_,
         intadd_18_SUM_0_, intadd_18_n3, intadd_18_n2, intadd_18_n1,
         intadd_19_A_1_, intadd_19_A_0_, intadd_19_B_2_, intadd_19_CI,
         intadd_19_SUM_2_, intadd_19_SUM_1_, intadd_19_SUM_0_, intadd_19_n3,
         intadd_19_n2, intadd_19_n1, intadd_0_A_36_, intadd_0_A_35_,
         intadd_0_A_34_, intadd_0_A_33_, intadd_0_A_31_, intadd_0_A_30_,
         intadd_0_A_29_, intadd_0_A_27_, intadd_0_A_26_, intadd_0_A_24_,
         intadd_0_A_23_, intadd_0_A_21_, intadd_0_A_20_, intadd_0_A_19_,
         intadd_0_A_18_, intadd_0_A_17_, intadd_0_A_16_, intadd_0_A_15_,
         intadd_0_A_14_, intadd_0_A_13_, intadd_0_A_12_, intadd_0_A_11_,
         intadd_0_A_10_, intadd_0_A_9_, intadd_0_A_8_, intadd_0_A_7_,
         intadd_0_A_6_, intadd_0_A_5_, intadd_0_A_4_, intadd_0_A_3_,
         intadd_0_A_2_, intadd_0_A_1_, intadd_0_A_0_, intadd_0_B_36_,
         intadd_0_B_35_, intadd_0_B_34_, intadd_0_B_32_, intadd_0_B_31_,
         intadd_0_B_30_, intadd_0_B_28_, intadd_0_B_27_, intadd_0_B_25_,
         intadd_0_B_24_, intadd_0_B_22_, intadd_0_B_21_, intadd_0_B_20_,
         intadd_0_B_19_, intadd_0_B_18_, intadd_0_B_17_, intadd_0_B_16_,
         intadd_0_B_15_, intadd_0_B_14_, intadd_0_B_13_, intadd_0_B_12_,
         intadd_0_B_11_, intadd_0_B_10_, intadd_0_B_9_, intadd_0_B_8_,
         intadd_0_B_7_, intadd_0_B_6_, intadd_0_B_5_, intadd_0_B_4_,
         intadd_0_B_3_, intadd_0_B_2_, intadd_0_B_1_, intadd_0_B_0_,
         intadd_0_CI, intadd_0_SUM_16_, intadd_0_SUM_15_, intadd_0_SUM_14_,
         intadd_0_SUM_13_, intadd_0_SUM_12_, intadd_0_SUM_11_,
         intadd_0_SUM_10_, intadd_0_SUM_9_, intadd_0_SUM_8_, intadd_0_SUM_7_,
         intadd_0_SUM_6_, intadd_0_SUM_5_, intadd_0_SUM_4_, intadd_0_SUM_3_,
         intadd_0_SUM_2_, intadd_0_SUM_1_, intadd_0_SUM_0_, intadd_0_n37,
         intadd_0_n36, intadd_0_n35, intadd_0_n34, intadd_0_n33, intadd_0_n32,
         intadd_0_n31, intadd_0_n30, intadd_0_n29, intadd_0_n28, intadd_0_n27,
         intadd_0_n26, intadd_0_n25, intadd_0_n24, intadd_0_n23, intadd_0_n22,
         intadd_0_n21, intadd_0_n20, intadd_0_n19, intadd_0_n18, intadd_0_n17,
         intadd_0_n16, intadd_0_n15, intadd_0_n14, intadd_0_n13, intadd_0_n12,
         intadd_0_n11, intadd_0_n10, intadd_0_n9, intadd_0_n8, intadd_0_n7,
         intadd_0_n6, intadd_0_n5, intadd_0_n4, intadd_0_n3, intadd_0_n2,
         intadd_0_n1, intadd_1_A_21_, intadd_1_A_20_, intadd_1_A_19_,
         intadd_1_A_18_, intadd_1_A_17_, intadd_1_A_16_, intadd_1_A_15_,
         intadd_1_A_14_, intadd_1_A_13_, intadd_1_A_12_, intadd_1_A_11_,
         intadd_1_A_10_, intadd_1_A_9_, intadd_1_A_8_, intadd_1_A_7_,
         intadd_1_A_6_, intadd_1_A_5_, intadd_1_A_4_, intadd_1_A_3_,
         intadd_1_A_2_, intadd_1_A_1_, intadd_1_A_0_, intadd_1_B_22_,
         intadd_1_B_21_, intadd_1_B_20_, intadd_1_B_19_, intadd_1_B_18_,
         intadd_1_B_17_, intadd_1_B_16_, intadd_1_B_15_, intadd_1_B_14_,
         intadd_1_B_13_, intadd_1_B_12_, intadd_1_B_11_, intadd_1_B_10_,
         intadd_1_B_9_, intadd_1_B_8_, intadd_1_B_7_, intadd_1_B_6_,
         intadd_1_B_5_, intadd_1_B_4_, intadd_1_B_3_, intadd_1_B_2_,
         intadd_1_B_1_, intadd_1_B_0_, intadd_1_CI, intadd_1_SUM_22_,
         intadd_1_SUM_21_, intadd_1_SUM_20_, intadd_1_SUM_19_,
         intadd_1_SUM_18_, intadd_1_SUM_17_, intadd_1_SUM_16_,
         intadd_1_SUM_15_, intadd_1_SUM_14_, intadd_1_SUM_13_,
         intadd_1_SUM_12_, intadd_1_SUM_11_, intadd_1_SUM_10_, intadd_1_SUM_9_,
         intadd_1_SUM_8_, intadd_1_SUM_7_, intadd_1_SUM_6_, intadd_1_SUM_5_,
         intadd_1_SUM_4_, intadd_1_SUM_3_, intadd_1_SUM_2_, intadd_1_SUM_1_,
         intadd_1_SUM_0_, intadd_1_n23, intadd_1_n22, intadd_1_n21,
         intadd_1_n20, intadd_1_n19, intadd_1_n18, intadd_1_n17, intadd_1_n16,
         intadd_1_n15, intadd_1_n14, intadd_1_n13, intadd_1_n12, intadd_1_n11,
         intadd_1_n10, intadd_1_n9, intadd_1_n8, intadd_1_n7, intadd_1_n6,
         intadd_1_n5, intadd_1_n4, intadd_1_n3, intadd_1_n2, intadd_1_n1,
         intadd_2_A_18_, intadd_2_A_17_, intadd_2_A_16_, intadd_2_A_15_,
         intadd_2_A_14_, intadd_2_A_13_, intadd_2_A_12_, intadd_2_A_11_,
         intadd_2_A_10_, intadd_2_A_9_, intadd_2_A_8_, intadd_2_A_7_,
         intadd_2_A_6_, intadd_2_A_5_, intadd_2_A_4_, intadd_2_A_3_,
         intadd_2_A_2_, intadd_2_A_1_, intadd_2_A_0_, intadd_2_B_18_,
         intadd_2_B_17_, intadd_2_B_16_, intadd_2_B_15_, intadd_2_B_14_,
         intadd_2_B_13_, intadd_2_B_12_, intadd_2_B_11_, intadd_2_B_10_,
         intadd_2_B_9_, intadd_2_B_8_, intadd_2_B_7_, intadd_2_B_6_,
         intadd_2_B_5_, intadd_2_B_4_, intadd_2_B_3_, intadd_2_B_2_,
         intadd_2_B_1_, intadd_2_B_0_, intadd_2_CI, intadd_2_n19, intadd_2_n18,
         intadd_2_n17, intadd_2_n16, intadd_2_n15, intadd_2_n14, intadd_2_n13,
         intadd_2_n12, intadd_2_n11, intadd_2_n10, intadd_2_n9, intadd_2_n8,
         intadd_2_n7, intadd_2_n6, intadd_2_n5, intadd_2_n4, intadd_2_n3,
         intadd_2_n2, intadd_2_n1, intadd_3_A_17_, intadd_3_B_17_,
         intadd_3_B_16_, intadd_3_B_15_, intadd_3_B_13_, intadd_3_B_12_,
         intadd_3_B_11_, intadd_3_B_10_, intadd_3_B_9_, intadd_3_B_8_,
         intadd_3_B_7_, intadd_3_B_6_, intadd_3_B_5_, intadd_3_B_4_,
         intadd_3_B_3_, intadd_3_B_2_, intadd_3_B_1_, intadd_3_B_0_,
         intadd_3_CI, intadd_3_SUM_17_, intadd_3_SUM_16_, intadd_3_SUM_15_,
         intadd_3_SUM_14_, intadd_3_SUM_13_, intadd_3_SUM_12_,
         intadd_3_SUM_11_, intadd_3_SUM_10_, intadd_3_SUM_9_, intadd_3_SUM_8_,
         intadd_3_SUM_7_, intadd_3_SUM_6_, intadd_3_SUM_5_, intadd_3_SUM_4_,
         intadd_3_SUM_3_, intadd_3_SUM_2_, intadd_3_SUM_1_, intadd_3_SUM_0_,
         intadd_3_n18, intadd_3_n17, intadd_3_n16, intadd_3_n15, intadd_3_n14,
         intadd_3_n13, intadd_3_n12, intadd_3_n11, intadd_3_n10, intadd_3_n9,
         intadd_3_n8, intadd_3_n7, intadd_3_n6, intadd_3_n5, intadd_3_n4,
         intadd_3_n3, intadd_3_n2, intadd_3_n1, intadd_4_A_13_, intadd_4_A_12_,
         intadd_4_A_11_, intadd_4_A_10_, intadd_4_A_9_, intadd_4_A_8_,
         intadd_4_A_7_, intadd_4_A_6_, intadd_4_A_5_, intadd_4_A_4_,
         intadd_4_A_3_, intadd_4_A_2_, intadd_4_A_1_, intadd_4_A_0_,
         intadd_4_B_16_, intadd_4_B_15_, intadd_4_B_14_, intadd_4_B_13_,
         intadd_4_B_12_, intadd_4_B_11_, intadd_4_B_10_, intadd_4_B_9_,
         intadd_4_B_8_, intadd_4_B_7_, intadd_4_B_6_, intadd_4_B_5_,
         intadd_4_B_4_, intadd_4_B_3_, intadd_4_B_2_, intadd_4_B_1_,
         intadd_4_B_0_, intadd_4_CI, intadd_4_SUM_16_, intadd_4_SUM_15_,
         intadd_4_SUM_14_, intadd_4_SUM_13_, intadd_4_SUM_12_,
         intadd_4_SUM_11_, intadd_4_SUM_10_, intadd_4_SUM_9_, intadd_4_SUM_8_,
         intadd_4_SUM_7_, intadd_4_SUM_6_, intadd_4_SUM_5_, intadd_4_SUM_4_,
         intadd_4_SUM_3_, intadd_4_SUM_2_, intadd_4_SUM_1_, intadd_4_SUM_0_,
         intadd_4_n17, intadd_4_n16, intadd_4_n15, intadd_4_n14, intadd_4_n13,
         intadd_4_n12, intadd_4_n11, intadd_4_n10, intadd_4_n9, intadd_4_n8,
         intadd_4_n7, intadd_4_n6, intadd_4_n5, intadd_4_n4, intadd_4_n3,
         intadd_4_n2, intadd_4_n1, intadd_6_A_10_, intadd_6_A_8_,
         intadd_6_A_7_, intadd_6_A_6_, intadd_6_A_5_, intadd_6_A_3_,
         intadd_6_A_2_, intadd_6_A_1_, intadd_6_A_0_, intadd_6_B_9_,
         intadd_6_B_4_, intadd_6_B_2_, intadd_6_B_1_, intadd_6_B_0_,
         intadd_6_CI, intadd_6_n11, intadd_6_n10, intadd_6_n9, intadd_6_n8,
         intadd_6_n7, intadd_6_n6, intadd_6_n5, intadd_6_n4, intadd_6_n3,
         intadd_6_n2, intadd_6_n1, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11,
         n12, n13, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n139, n140, n142, n143, n144, n145, n147,
         n149, n150, n152, n153, n154, n159, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n175, n176, n178, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419;
  wire   [3:0] state;
  wire   [29:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [23:0] a_m;
  wire   [9:0] b_e;
  wire   [23:0] b_m;
  wire   [49:2] product;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ao211d1_hd U246 ( .A(n1544), .B(n155), .C(i_RST), .D(n501), .Y(n350) );
  oa22d1_hd U247 ( .A(n156), .B(n157), .C(n1628), .D(n158), .Y(n351) );
  oa22d1_hd U249 ( .A(n160), .B(n157), .C(n74), .D(n158), .Y(n352) );
  oa22d1_hd U250 ( .A(n161), .B(n157), .C(n1629), .D(n158), .Y(n353) );
  oa22d1_hd U267 ( .A(n171), .B(n157), .C(n1614), .D(n158), .Y(n357) );
  nd4d1_hd U269 ( .A(n160), .B(n172), .C(n173), .D(n174), .Y(n158) );
  ao211d1_hd U270 ( .A(n3279), .B(n36), .C(i_RST), .D(n500), .Y(n174) );
  ao211d1_hd U281 ( .A(n475), .B(n177), .C(i_RST), .D(n179), .Y(n358) );
  ivd1_hd U364 ( .A(i_RST), .Y(N34) );
  fad1_hd DP_OP_116J2_127_7148_U6 ( .A(n378), .B(n1213), .CI(
        DP_OP_116J2_127_7148_n4), .CO(DP_OP_116J2_127_7148_n3), .S(C82_DATA2_6) );
  fad1_hd DP_OP_116J2_127_7148_U7 ( .A(n379), .B(n1212), .CI(
        DP_OP_116J2_127_7148_n5), .CO(DP_OP_116J2_127_7148_n4), .S(C82_DATA2_5) );
  fad1_hd DP_OP_116J2_127_7148_U8 ( .A(n380), .B(n1211), .CI(
        DP_OP_116J2_127_7148_n6), .CO(DP_OP_116J2_127_7148_n5), .S(C82_DATA2_4) );
  fad1_hd DP_OP_116J2_127_7148_U9 ( .A(n378), .B(n1210), .CI(
        DP_OP_116J2_127_7148_n7), .CO(DP_OP_116J2_127_7148_n6), .S(C82_DATA2_3) );
  fad1_hd DP_OP_116J2_127_7148_U10 ( .A(n378), .B(n1209), .CI(
        DP_OP_116J2_127_7148_n8), .CO(DP_OP_116J2_127_7148_n7), .S(C82_DATA2_2) );
  fad1_hd DP_OP_116J2_127_7148_U11 ( .A(n379), .B(n1208), .CI(n1207), .CO(
        DP_OP_116J2_127_7148_n8), .S(C82_DATA2_1) );
  fad1_hd DP_OP_113J2_124_6892_U6 ( .A(n379), .B(C1_Z_6), .CI(
        DP_OP_113J2_124_6892_n4), .CO(DP_OP_113J2_124_6892_n3), .S(C81_DATA2_6) );
  fad1_hd DP_OP_113J2_124_6892_U7 ( .A(n380), .B(C1_Z_5), .CI(
        DP_OP_113J2_124_6892_n5), .CO(DP_OP_113J2_124_6892_n4), .S(C81_DATA2_5) );
  fad1_hd DP_OP_113J2_124_6892_U8 ( .A(n378), .B(C1_Z_4), .CI(
        DP_OP_113J2_124_6892_n6), .CO(DP_OP_113J2_124_6892_n5), .S(C81_DATA2_4) );
  fad1_hd DP_OP_113J2_124_6892_U9 ( .A(n379), .B(C1_Z_3), .CI(
        DP_OP_113J2_124_6892_n7), .CO(DP_OP_113J2_124_6892_n6), .S(C81_DATA2_3) );
  fad1_hd DP_OP_113J2_124_6892_U10 ( .A(n379), .B(C1_Z_2), .CI(
        DP_OP_113J2_124_6892_n8), .CO(DP_OP_113J2_124_6892_n7), .S(C81_DATA2_2) );
  fad1_hd DP_OP_113J2_124_6892_U11 ( .A(n380), .B(C1_Z_1), .CI(n1206), .CO(
        DP_OP_113J2_124_6892_n8), .S(C81_DATA2_1) );
  had1_hd DP_OP_125J2_130_6300_U32 ( .A(b_e[0]), .B(a_e[0]), .CO(
        DP_OP_125J2_130_6300_n20), .S(DP_OP_125J2_130_6300_n34) );
  fad1_hd DP_OP_125J2_130_6300_U31 ( .A(a_e[1]), .B(b_e[1]), .CI(
        DP_OP_125J2_130_6300_n20), .CO(DP_OP_125J2_130_6300_n19), .S(
        DP_OP_125J2_130_6300_n35) );
  fad1_hd DP_OP_125J2_130_6300_U30 ( .A(a_e[2]), .B(b_e[2]), .CI(
        DP_OP_125J2_130_6300_n19), .CO(DP_OP_125J2_130_6300_n18), .S(
        DP_OP_125J2_130_6300_n36) );
  fad1_hd DP_OP_125J2_130_6300_U29 ( .A(a_e[3]), .B(b_e[3]), .CI(
        DP_OP_125J2_130_6300_n18), .CO(DP_OP_125J2_130_6300_n17), .S(
        DP_OP_125J2_130_6300_n37) );
  fad1_hd DP_OP_125J2_130_6300_U28 ( .A(a_e[4]), .B(b_e[4]), .CI(
        DP_OP_125J2_130_6300_n17), .CO(DP_OP_125J2_130_6300_n16), .S(
        DP_OP_125J2_130_6300_n38) );
  fad1_hd DP_OP_125J2_130_6300_U27 ( .A(a_e[5]), .B(b_e[5]), .CI(
        DP_OP_125J2_130_6300_n16), .CO(DP_OP_125J2_130_6300_n15), .S(
        DP_OP_125J2_130_6300_n39) );
  fad1_hd DP_OP_125J2_130_6300_U26 ( .A(a_e[6]), .B(b_e[6]), .CI(
        DP_OP_125J2_130_6300_n15), .CO(DP_OP_125J2_130_6300_n14), .S(
        DP_OP_125J2_130_6300_n40) );
  fad1_hd DP_OP_125J2_130_6300_U25 ( .A(a_e[7]), .B(b_e[7]), .CI(
        DP_OP_125J2_130_6300_n14), .CO(DP_OP_125J2_130_6300_n13), .S(
        DP_OP_125J2_130_6300_n41) );
  fad1_hd DP_OP_125J2_130_6300_U24 ( .A(a_e[8]), .B(b_e[8]), .CI(
        DP_OP_125J2_130_6300_n13), .CO(DP_OP_125J2_130_6300_n12), .S(
        DP_OP_125J2_130_6300_n42) );
  fad1_hd DP_OP_125J2_130_6300_U10 ( .A(n1613), .B(n376), .CI(
        DP_OP_125J2_130_6300_n25), .CO(DP_OP_125J2_130_6300_n9), .S(N467) );
  fad1_hd DP_OP_125J2_130_6300_U9 ( .A(DP_OP_125J2_130_6300_n26), .B(n377), 
        .CI(DP_OP_125J2_130_6300_n9), .CO(DP_OP_125J2_130_6300_n8), .S(N468)
         );
  fad1_hd DP_OP_125J2_130_6300_U8 ( .A(DP_OP_125J2_130_6300_n27), .B(n376), 
        .CI(DP_OP_125J2_130_6300_n8), .CO(DP_OP_125J2_130_6300_n7), .S(N469)
         );
  fad1_hd DP_OP_125J2_130_6300_U7 ( .A(DP_OP_125J2_130_6300_n28), .B(n377), 
        .CI(DP_OP_125J2_130_6300_n7), .CO(DP_OP_125J2_130_6300_n6), .S(N470)
         );
  fad1_hd DP_OP_125J2_130_6300_U6 ( .A(DP_OP_125J2_130_6300_n29), .B(n376), 
        .CI(DP_OP_125J2_130_6300_n6), .CO(DP_OP_125J2_130_6300_n5), .S(N471)
         );
  fad1_hd DP_OP_125J2_130_6300_U5 ( .A(DP_OP_125J2_130_6300_n30), .B(n377), 
        .CI(DP_OP_125J2_130_6300_n5), .CO(DP_OP_125J2_130_6300_n4), .S(N472)
         );
  fad1_hd DP_OP_125J2_130_6300_U4 ( .A(DP_OP_125J2_130_6300_n31), .B(n376), 
        .CI(DP_OP_125J2_130_6300_n4), .CO(DP_OP_125J2_130_6300_n3), .S(N473)
         );
  fad1_hd DP_OP_125J2_130_6300_U3 ( .A(DP_OP_125J2_130_6300_n32), .B(n377), 
        .CI(DP_OP_125J2_130_6300_n3), .CO(DP_OP_125J2_130_6300_n2), .S(N474)
         );
  fds2d1_hd a_e_reg_7_ ( .CRN(n141), .D(n138), .CK(i_CLK), .Q(n10), .QN(a_e[7]) );
  fds2d1_hd b_e_reg_7_ ( .CRN(n151), .D(n148), .CK(i_CLK), .Q(n14), .QN(b_e[7]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n319), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n356), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n309), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n306), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n290), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n291), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n292), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n295), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n296), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n299), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n305), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n294), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd z_reg_28_ ( .D(n232), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n234), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_29_ ( .D(n231), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_24_ ( .D(n236), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n237), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n289), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n297), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n298), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n302), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n301), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n287), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd z_reg_27_ ( .D(n233), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n304), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n293), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n303), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n300), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd z_reg_17_ ( .D(n243), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n244), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_1_ ( .D(n259), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_0_ ( .D(n260), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_2_ ( .D(n258), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n288), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n326), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n317), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd z_reg_13_ ( .D(n247), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n248), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_9_ ( .D(n251), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n252), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_5_ ( .D(n255), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_4_ ( .D(n256), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_10_ ( .D(n250), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_7_ ( .D(n253), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n254), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_3_ ( .D(n257), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n327), .CK(i_CLK), .Q(b_e[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n318), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n325), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n316), .CK(i_CLK), .Q(a_e[2]) );
  fd1qd1_hd state_reg_3_ ( .D(n357), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd state_reg_2_ ( .D(n351), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_0_ ( .D(n353), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd state_reg_1_ ( .D(n352), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n315), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n324), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n323), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n314), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n282), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n322), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n313), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n281), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n285), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n312), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n321), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n262), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n276), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n264), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n280), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n268), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n272), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n261), .CK(i_CLK), .Q(z_m[22]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n270), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n266), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n274), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n278), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n269), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n265), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n277), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n273), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n275), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n267), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n279), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n271), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n263), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n286), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n320), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n311), .CK(i_CLK), .Q(a_e[8]) );
  clknd2d1_hd U552 ( .A(N34), .B(n158), .Y(n157) );
  fad1_hd intadd_5_U13 ( .A(intadd_5_A_0_), .B(intadd_5_B_0_), .CI(intadd_5_CI), .CO(intadd_5_n12), .S(intadd_5_SUM_0_) );
  fad1_hd intadd_5_U12 ( .A(intadd_5_A_1_), .B(intadd_5_B_1_), .CI(
        intadd_5_n12), .CO(intadd_5_n11), .S(intadd_5_SUM_1_) );
  fad1_hd intadd_5_U11 ( .A(intadd_5_A_2_), .B(intadd_5_B_2_), .CI(
        intadd_5_n11), .CO(intadd_5_n10), .S(intadd_5_SUM_2_) );
  fad1_hd intadd_5_U10 ( .A(intadd_5_A_3_), .B(intadd_5_B_3_), .CI(
        intadd_5_n10), .CO(intadd_5_n9), .S(intadd_5_SUM_3_) );
  fad1_hd intadd_5_U9 ( .A(intadd_5_A_4_), .B(intadd_5_B_4_), .CI(intadd_5_n9), 
        .CO(intadd_5_n8), .S(intadd_5_SUM_4_) );
  fad1_hd intadd_5_U8 ( .A(intadd_5_A_5_), .B(intadd_5_B_5_), .CI(intadd_5_n8), 
        .CO(intadd_5_n7), .S(intadd_5_SUM_5_) );
  fad1_hd intadd_5_U7 ( .A(intadd_5_A_6_), .B(intadd_5_B_6_), .CI(intadd_5_n7), 
        .CO(intadd_5_n6), .S(intadd_5_SUM_6_) );
  fad1_hd intadd_5_U6 ( .A(intadd_5_A_7_), .B(intadd_5_B_7_), .CI(intadd_5_n6), 
        .CO(intadd_5_n5), .S(intadd_5_SUM_7_) );
  fad1_hd intadd_5_U5 ( .A(intadd_5_A_8_), .B(intadd_5_B_8_), .CI(intadd_5_n5), 
        .CO(intadd_5_n4), .S(intadd_5_SUM_8_) );
  fad1_hd intadd_5_U4 ( .A(intadd_5_A_9_), .B(intadd_5_B_9_), .CI(intadd_5_n4), 
        .CO(intadd_5_n3), .S(intadd_5_SUM_9_) );
  fad1_hd intadd_5_U3 ( .A(intadd_5_A_10_), .B(intadd_5_B_10_), .CI(
        intadd_5_n3), .CO(intadd_5_n2), .S(intadd_5_SUM_10_) );
  fad1_hd intadd_5_U2 ( .A(intadd_5_A_11_), .B(intadd_5_B_11_), .CI(
        intadd_5_n2), .CO(intadd_5_n1), .S(intadd_5_SUM_11_) );
  fad1_hd intadd_7_U12 ( .A(intadd_7_A_0_), .B(intadd_7_B_0_), .CI(intadd_7_CI), .CO(intadd_7_n11), .S(intadd_7_SUM_0_) );
  fad1_hd intadd_7_U11 ( .A(intadd_7_A_1_), .B(intadd_7_B_1_), .CI(
        intadd_7_n11), .CO(intadd_7_n10), .S(intadd_7_SUM_1_) );
  fad1_hd intadd_7_U10 ( .A(intadd_7_A_2_), .B(intadd_7_B_2_), .CI(
        intadd_7_n10), .CO(intadd_7_n9), .S(intadd_7_SUM_2_) );
  fad1_hd intadd_7_U9 ( .A(intadd_7_A_3_), .B(intadd_7_B_3_), .CI(intadd_7_n9), 
        .CO(intadd_7_n8), .S(intadd_7_SUM_3_) );
  fad1_hd intadd_7_U8 ( .A(intadd_7_A_4_), .B(intadd_7_B_4_), .CI(intadd_7_n8), 
        .CO(intadd_7_n7), .S(intadd_7_SUM_4_) );
  fad1_hd intadd_7_U7 ( .A(intadd_7_A_5_), .B(intadd_7_B_5_), .CI(intadd_7_n7), 
        .CO(intadd_7_n6), .S(intadd_7_SUM_5_) );
  fad1_hd intadd_7_U6 ( .A(intadd_7_A_6_), .B(intadd_7_B_6_), .CI(intadd_7_n6), 
        .CO(intadd_7_n5), .S(intadd_7_SUM_6_) );
  fad1_hd intadd_7_U5 ( .A(intadd_7_A_7_), .B(intadd_7_B_7_), .CI(intadd_7_n5), 
        .CO(intadd_7_n4), .S(intadd_7_SUM_7_) );
  fad1_hd intadd_7_U4 ( .A(intadd_7_A_8_), .B(intadd_7_B_8_), .CI(intadd_7_n4), 
        .CO(intadd_7_n3), .S(intadd_7_SUM_8_) );
  fad1_hd intadd_7_U3 ( .A(intadd_7_A_9_), .B(intadd_7_B_9_), .CI(intadd_7_n3), 
        .CO(intadd_7_n2), .S(intadd_7_SUM_9_) );
  fad1_hd intadd_8_U10 ( .A(a_m[2]), .B(intadd_8_B_0_), .CI(intadd_8_CI), .CO(
        intadd_8_n9), .S(intadd_8_SUM_0_) );
  fad1_hd intadd_8_U9 ( .A(intadd_8_A_1_), .B(intadd_8_B_1_), .CI(intadd_8_n9), 
        .CO(intadd_8_n8), .S(intadd_7_A_6_) );
  fad1_hd intadd_8_U8 ( .A(intadd_8_A_2_), .B(intadd_8_B_2_), .CI(intadd_8_n8), 
        .CO(intadd_8_n7), .S(intadd_7_A_7_) );
  fad1_hd intadd_8_U7 ( .A(intadd_8_A_3_), .B(intadd_8_B_3_), .CI(intadd_8_n7), 
        .CO(intadd_8_n6), .S(intadd_7_A_8_) );
  fad1_hd intadd_8_U6 ( .A(intadd_12_n1), .B(intadd_8_B_4_), .CI(intadd_8_n6), 
        .CO(intadd_8_n5), .S(intadd_8_SUM_4_) );
  fad1_hd intadd_8_U5 ( .A(intadd_8_A_5_), .B(intadd_8_B_5_), .CI(intadd_8_n5), 
        .CO(intadd_8_n4), .S(intadd_8_SUM_5_) );
  fad1_hd intadd_8_U4 ( .A(intadd_8_A_6_), .B(intadd_8_B_6_), .CI(intadd_8_n4), 
        .CO(intadd_8_n3), .S(intadd_8_SUM_6_) );
  fad1_hd intadd_8_U3 ( .A(intadd_8_A_7_), .B(intadd_8_B_7_), .CI(intadd_8_n3), 
        .CO(intadd_8_n2), .S(intadd_8_SUM_7_) );
  fad1_hd intadd_9_U9 ( .A(a_m[5]), .B(n197), .CI(intadd_9_CI), .CO(
        intadd_9_n8), .S(intadd_9_SUM_0_) );
  fad1_hd intadd_9_U8 ( .A(intadd_9_A_1_), .B(intadd_9_B_1_), .CI(intadd_9_n8), 
        .CO(intadd_9_n7), .S(intadd_9_SUM_1_) );
  fad1_hd intadd_9_U7 ( .A(intadd_9_A_2_), .B(intadd_9_B_2_), .CI(intadd_9_n7), 
        .CO(intadd_9_n6), .S(intadd_9_SUM_2_) );
  fad1_hd intadd_9_U6 ( .A(intadd_9_A_3_), .B(intadd_9_B_3_), .CI(intadd_9_n6), 
        .CO(intadd_9_n5), .S(intadd_9_SUM_3_) );
  fad1_hd intadd_9_U5 ( .A(intadd_9_A_4_), .B(intadd_9_B_4_), .CI(intadd_9_n5), 
        .CO(intadd_9_n4), .S(intadd_9_SUM_4_) );
  fad1_hd intadd_9_U4 ( .A(intadd_9_A_5_), .B(intadd_9_B_5_), .CI(intadd_9_n4), 
        .CO(intadd_9_n3), .S(intadd_9_SUM_5_) );
  fad1_hd intadd_9_U3 ( .A(intadd_9_A_6_), .B(intadd_9_B_6_), .CI(intadd_9_n3), 
        .CO(intadd_9_n2), .S(intadd_9_SUM_6_) );
  fad1_hd intadd_9_U2 ( .A(intadd_9_A_7_), .B(intadd_9_B_7_), .CI(intadd_9_n2), 
        .CO(intadd_9_n1), .S(intadd_9_SUM_7_) );
  fad1_hd intadd_10_U7 ( .A(intadd_10_A_0_), .B(intadd_10_B_0_), .CI(
        intadd_10_CI), .CO(intadd_10_n6), .S(intadd_10_SUM_0_) );
  fad1_hd intadd_10_U6 ( .A(intadd_10_A_1_), .B(intadd_10_B_1_), .CI(
        intadd_10_n6), .CO(intadd_10_n5), .S(intadd_10_SUM_1_) );
  fad1_hd intadd_10_U5 ( .A(intadd_10_A_2_), .B(intadd_10_B_2_), .CI(
        intadd_10_n5), .CO(intadd_10_n4), .S(intadd_10_SUM_2_) );
  fad1_hd intadd_10_U4 ( .A(intadd_10_A_3_), .B(intadd_10_B_3_), .CI(
        intadd_10_n4), .CO(intadd_10_n3), .S(intadd_10_SUM_3_) );
  fad1_hd intadd_10_U3 ( .A(intadd_10_A_4_), .B(intadd_10_B_4_), .CI(
        intadd_10_n3), .CO(intadd_10_n2), .S(intadd_10_SUM_4_) );
  fad1_hd intadd_11_U6 ( .A(intadd_11_A_0_), .B(intadd_11_B_0_), .CI(
        intadd_11_CI), .CO(intadd_11_n5), .S(intadd_11_SUM_0_) );
  fad1_hd intadd_11_U5 ( .A(intadd_11_A_1_), .B(intadd_11_B_1_), .CI(
        intadd_11_n5), .CO(intadd_11_n4), .S(intadd_11_SUM_1_) );
  fad1_hd intadd_11_U4 ( .A(intadd_11_A_2_), .B(intadd_11_B_2_), .CI(
        intadd_11_n4), .CO(intadd_11_n3), .S(intadd_11_SUM_2_) );
  fad1_hd intadd_11_U3 ( .A(intadd_11_A_3_), .B(intadd_11_B_3_), .CI(
        intadd_11_n3), .CO(intadd_11_n2), .S(intadd_11_SUM_3_) );
  fad1_hd intadd_12_U4 ( .A(n196), .B(intadd_12_B_0_), .CI(intadd_12_CI), .CO(
        intadd_12_n3), .S(intadd_8_B_1_) );
  fad1_hd intadd_12_U3 ( .A(intadd_12_A_1_), .B(intadd_12_B_1_), .CI(
        intadd_12_n3), .CO(intadd_12_n2), .S(intadd_8_A_2_) );
  fad1_hd intadd_12_U2 ( .A(intadd_12_A_2_), .B(intadd_12_B_2_), .CI(
        intadd_12_n2), .CO(intadd_12_n1), .S(intadd_8_A_3_) );
  fad1_hd intadd_13_U4 ( .A(intadd_13_A_0_), .B(intadd_13_B_0_), .CI(
        intadd_13_CI), .CO(intadd_13_n3), .S(intadd_13_SUM_0_) );
  fad1_hd intadd_13_U3 ( .A(intadd_13_A_1_), .B(intadd_13_B_1_), .CI(
        intadd_13_n3), .CO(intadd_13_n2), .S(intadd_13_SUM_1_) );
  fad1_hd intadd_14_U3 ( .A(intadd_14_A_1_), .B(intadd_14_B_1_), .CI(
        intadd_14_n3), .CO(intadd_14_n2), .S(intadd_14_SUM_1_) );
  fad1_hd intadd_14_U2 ( .A(intadd_14_A_2_), .B(intadd_14_B_2_), .CI(
        intadd_14_n2), .CO(intadd_14_n1), .S(intadd_14_SUM_2_) );
  fad1_hd intadd_15_U4 ( .A(intadd_15_A_0_), .B(intadd_15_B_0_), .CI(
        intadd_10_SUM_1_), .CO(intadd_15_n3), .S(intadd_15_SUM_0_) );
  fad1_hd intadd_15_U3 ( .A(intadd_10_SUM_2_), .B(intadd_15_B_1_), .CI(
        intadd_15_n3), .CO(intadd_15_n2), .S(intadd_15_SUM_1_) );
  fad1_hd intadd_16_U4 ( .A(intadd_9_SUM_5_), .B(intadd_16_B_0_), .CI(
        intadd_16_CI), .CO(intadd_16_n3), .S(intadd_16_SUM_0_) );
  fad1_hd intadd_16_U3 ( .A(intadd_9_SUM_6_), .B(intadd_16_B_1_), .CI(
        intadd_16_n3), .CO(intadd_16_n2), .S(intadd_16_SUM_1_) );
  fad1_hd intadd_17_U4 ( .A(intadd_17_A_0_), .B(intadd_17_B_0_), .CI(
        intadd_17_CI), .CO(intadd_17_n3), .S(intadd_17_SUM_0_) );
  fad1_hd intadd_17_U3 ( .A(intadd_17_A_1_), .B(intadd_17_B_1_), .CI(
        intadd_17_n3), .CO(intadd_17_n2), .S(intadd_17_SUM_1_) );
  fad1_hd intadd_18_U4 ( .A(intadd_9_SUM_2_), .B(intadd_18_B_0_), .CI(
        intadd_18_CI), .CO(intadd_18_n3), .S(intadd_18_SUM_0_) );
  fad1_hd intadd_18_U3 ( .A(intadd_9_SUM_3_), .B(intadd_18_B_1_), .CI(
        intadd_18_n3), .CO(intadd_18_n2), .S(intadd_18_SUM_1_) );
  fad1_hd intadd_18_U2 ( .A(intadd_9_SUM_4_), .B(intadd_18_B_2_), .CI(
        intadd_18_n2), .CO(intadd_18_n1), .S(intadd_18_SUM_2_) );
  fad1_hd intadd_19_U4 ( .A(intadd_19_A_0_), .B(intadd_5_SUM_9_), .CI(
        intadd_19_CI), .CO(intadd_19_n3), .S(intadd_19_SUM_0_) );
  fad1_hd intadd_19_U3 ( .A(intadd_19_A_1_), .B(intadd_5_SUM_10_), .CI(
        intadd_19_n3), .CO(intadd_19_n2), .S(intadd_19_SUM_1_) );
  fad1_hd intadd_19_U2 ( .A(intadd_5_SUM_11_), .B(intadd_19_B_2_), .CI(
        intadd_19_n2), .CO(intadd_19_n1), .S(intadd_19_SUM_2_) );
  fad1_hd intadd_0_U38 ( .A(intadd_0_A_0_), .B(intadd_0_B_0_), .CI(intadd_0_CI), .CO(intadd_0_n37), .S(intadd_0_SUM_0_) );
  fad1_hd intadd_0_U37 ( .A(intadd_0_A_1_), .B(intadd_0_B_1_), .CI(
        intadd_0_n37), .CO(intadd_0_n36), .S(intadd_0_SUM_1_) );
  fad1_hd intadd_0_U36 ( .A(intadd_0_A_2_), .B(intadd_0_B_2_), .CI(
        intadd_0_n36), .CO(intadd_0_n35), .S(intadd_0_SUM_2_) );
  fad1_hd intadd_0_U35 ( .A(intadd_0_A_3_), .B(intadd_0_B_3_), .CI(
        intadd_0_n35), .CO(intadd_0_n34), .S(intadd_0_SUM_3_) );
  fad1_hd intadd_0_U34 ( .A(intadd_0_A_4_), .B(intadd_0_B_4_), .CI(
        intadd_0_n34), .CO(intadd_0_n33), .S(intadd_0_SUM_4_) );
  fad1_hd intadd_0_U33 ( .A(intadd_0_A_5_), .B(intadd_0_B_5_), .CI(
        intadd_0_n33), .CO(intadd_0_n32), .S(intadd_0_SUM_5_) );
  fad1_hd intadd_0_U32 ( .A(intadd_0_A_6_), .B(intadd_0_B_6_), .CI(
        intadd_0_n32), .CO(intadd_0_n31), .S(intadd_0_SUM_6_) );
  fad1_hd intadd_0_U31 ( .A(intadd_0_A_7_), .B(intadd_0_B_7_), .CI(
        intadd_0_n31), .CO(intadd_0_n30), .S(intadd_0_SUM_7_) );
  fad1_hd intadd_0_U30 ( .A(intadd_0_A_8_), .B(intadd_0_B_8_), .CI(
        intadd_0_n30), .CO(intadd_0_n29), .S(intadd_0_SUM_8_) );
  fad1_hd intadd_0_U29 ( .A(intadd_0_A_9_), .B(intadd_0_B_9_), .CI(
        intadd_0_n29), .CO(intadd_0_n28), .S(intadd_0_SUM_9_) );
  fad1_hd intadd_0_U28 ( .A(intadd_0_A_10_), .B(intadd_0_B_10_), .CI(
        intadd_0_n28), .CO(intadd_0_n27), .S(intadd_0_SUM_10_) );
  fad1_hd intadd_0_U27 ( .A(intadd_0_A_11_), .B(intadd_0_B_11_), .CI(
        intadd_0_n27), .CO(intadd_0_n26), .S(intadd_0_SUM_11_) );
  fad1_hd intadd_0_U26 ( .A(intadd_0_A_12_), .B(intadd_0_B_12_), .CI(
        intadd_0_n26), .CO(intadd_0_n25), .S(intadd_0_SUM_12_) );
  fad1_hd intadd_0_U25 ( .A(intadd_0_A_13_), .B(intadd_0_B_13_), .CI(
        intadd_0_n25), .CO(intadd_0_n24), .S(intadd_0_SUM_13_) );
  fad1_hd intadd_0_U24 ( .A(intadd_0_A_14_), .B(intadd_0_B_14_), .CI(
        intadd_0_n24), .CO(intadd_0_n23), .S(intadd_0_SUM_14_) );
  fad1_hd intadd_0_U23 ( .A(intadd_0_A_15_), .B(intadd_0_B_15_), .CI(
        intadd_0_n23), .CO(intadd_0_n22), .S(intadd_0_SUM_15_) );
  fad1_hd intadd_0_U22 ( .A(intadd_0_A_16_), .B(intadd_0_B_16_), .CI(
        intadd_0_n22), .CO(intadd_0_n21), .S(intadd_0_SUM_16_) );
  fad1_hd intadd_1_U24 ( .A(intadd_1_A_0_), .B(intadd_1_B_0_), .CI(intadd_1_CI), .CO(intadd_1_n23), .S(intadd_1_SUM_0_) );
  fad1_hd intadd_1_U23 ( .A(intadd_1_A_1_), .B(intadd_1_B_1_), .CI(
        intadd_1_n23), .CO(intadd_1_n22), .S(intadd_1_SUM_1_) );
  fad1_hd intadd_1_U22 ( .A(intadd_1_A_2_), .B(intadd_1_B_2_), .CI(
        intadd_1_n22), .CO(intadd_1_n21), .S(intadd_1_SUM_2_) );
  fad1_hd intadd_1_U21 ( .A(intadd_1_A_3_), .B(intadd_1_B_3_), .CI(
        intadd_1_n21), .CO(intadd_1_n20), .S(intadd_1_SUM_3_) );
  fad1_hd intadd_1_U20 ( .A(intadd_1_A_4_), .B(intadd_1_B_4_), .CI(
        intadd_1_n20), .CO(intadd_1_n19), .S(intadd_1_SUM_4_) );
  fad1_hd intadd_1_U19 ( .A(intadd_1_A_5_), .B(intadd_1_B_5_), .CI(
        intadd_1_n19), .CO(intadd_1_n18), .S(intadd_1_SUM_5_) );
  fad1_hd intadd_1_U18 ( .A(intadd_1_A_6_), .B(intadd_1_B_6_), .CI(
        intadd_1_n18), .CO(intadd_1_n17), .S(intadd_1_SUM_6_) );
  fad1_hd intadd_1_U17 ( .A(intadd_1_A_7_), .B(intadd_1_B_7_), .CI(
        intadd_1_n17), .CO(intadd_1_n16), .S(intadd_1_SUM_7_) );
  fad1_hd intadd_1_U16 ( .A(intadd_1_A_8_), .B(intadd_1_B_8_), .CI(
        intadd_1_n16), .CO(intadd_1_n15), .S(intadd_1_SUM_8_) );
  fad1_hd intadd_1_U15 ( .A(intadd_1_A_9_), .B(intadd_1_B_9_), .CI(
        intadd_1_n15), .CO(intadd_1_n14), .S(intadd_1_SUM_9_) );
  fad1_hd intadd_1_U14 ( .A(intadd_1_A_10_), .B(intadd_1_B_10_), .CI(
        intadd_1_n14), .CO(intadd_1_n13), .S(intadd_1_SUM_10_) );
  fad1_hd intadd_1_U13 ( .A(intadd_1_A_11_), .B(intadd_1_B_11_), .CI(
        intadd_1_n13), .CO(intadd_1_n12), .S(intadd_1_SUM_11_) );
  fad1_hd intadd_1_U12 ( .A(intadd_1_A_12_), .B(intadd_1_B_12_), .CI(
        intadd_1_n12), .CO(intadd_1_n11), .S(intadd_1_SUM_12_) );
  fad1_hd intadd_1_U11 ( .A(intadd_1_A_13_), .B(intadd_1_B_13_), .CI(
        intadd_1_n11), .CO(intadd_1_n10), .S(intadd_1_SUM_13_) );
  fad1_hd intadd_1_U10 ( .A(intadd_1_A_14_), .B(intadd_1_B_14_), .CI(
        intadd_1_n10), .CO(intadd_1_n9), .S(intadd_1_SUM_14_) );
  fad1_hd intadd_1_U9 ( .A(intadd_1_A_15_), .B(intadd_1_B_15_), .CI(
        intadd_1_n9), .CO(intadd_1_n8), .S(intadd_1_SUM_15_) );
  fad1_hd intadd_1_U8 ( .A(intadd_1_A_16_), .B(intadd_1_B_16_), .CI(
        intadd_1_n8), .CO(intadd_1_n7), .S(intadd_1_SUM_16_) );
  fad1_hd intadd_1_U7 ( .A(intadd_1_A_17_), .B(intadd_1_B_17_), .CI(
        intadd_1_n7), .CO(intadd_1_n6), .S(intadd_1_SUM_17_) );
  fad1_hd intadd_1_U6 ( .A(intadd_1_A_18_), .B(intadd_1_B_18_), .CI(
        intadd_1_n6), .CO(intadd_1_n5), .S(intadd_1_SUM_18_) );
  fad1_hd intadd_1_U5 ( .A(intadd_1_A_19_), .B(intadd_1_B_19_), .CI(
        intadd_1_n5), .CO(intadd_1_n4), .S(intadd_1_SUM_19_) );
  fad1_hd intadd_1_U4 ( .A(intadd_1_A_20_), .B(intadd_1_B_20_), .CI(
        intadd_1_n4), .CO(intadd_1_n3), .S(intadd_1_SUM_20_) );
  fad1_hd intadd_1_U2 ( .A(intadd_2_n1), .B(intadd_1_B_22_), .CI(intadd_1_n2), 
        .CO(intadd_1_n1), .S(intadd_1_SUM_22_) );
  fad1_hd intadd_2_U20 ( .A(intadd_2_A_0_), .B(intadd_2_B_0_), .CI(intadd_2_CI), .CO(intadd_2_n19), .S(intadd_1_A_3_) );
  fad1_hd intadd_2_U19 ( .A(intadd_2_A_1_), .B(intadd_2_B_1_), .CI(
        intadd_2_n19), .CO(intadd_2_n18), .S(intadd_1_A_4_) );
  fad1_hd intadd_2_U15 ( .A(intadd_2_A_5_), .B(intadd_2_B_5_), .CI(
        intadd_2_n15), .CO(intadd_2_n14), .S(intadd_1_A_8_) );
  fad1_hd intadd_2_U13 ( .A(intadd_2_A_7_), .B(intadd_2_B_7_), .CI(
        intadd_2_n13), .CO(intadd_2_n12), .S(intadd_1_A_10_) );
  fad1_hd intadd_2_U12 ( .A(intadd_2_A_8_), .B(intadd_2_B_8_), .CI(
        intadd_2_n12), .CO(intadd_2_n11), .S(intadd_1_A_11_) );
  fad1_hd intadd_2_U11 ( .A(intadd_2_A_9_), .B(intadd_2_B_9_), .CI(
        intadd_2_n11), .CO(intadd_2_n10), .S(intadd_1_A_12_) );
  fad1_hd intadd_2_U10 ( .A(intadd_2_A_10_), .B(intadd_2_B_10_), .CI(
        intadd_2_n10), .CO(intadd_2_n9), .S(intadd_1_B_13_) );
  fad1_hd intadd_2_U6 ( .A(intadd_2_A_14_), .B(intadd_2_B_14_), .CI(
        intadd_2_n6), .CO(intadd_2_n5), .S(intadd_1_B_17_) );
  fad1_hd intadd_2_U5 ( .A(intadd_2_A_15_), .B(intadd_2_B_15_), .CI(
        intadd_2_n5), .CO(intadd_2_n4), .S(intadd_1_B_18_) );
  fad1_hd intadd_2_U4 ( .A(intadd_2_A_16_), .B(intadd_2_B_16_), .CI(
        intadd_2_n4), .CO(intadd_2_n3), .S(intadd_1_B_19_) );
  fad1_hd intadd_4_U18 ( .A(intadd_4_A_0_), .B(intadd_4_B_0_), .CI(intadd_4_CI), .CO(intadd_4_n17), .S(intadd_4_SUM_0_) );
  fad1_hd intadd_4_U17 ( .A(intadd_4_A_1_), .B(intadd_4_B_1_), .CI(
        intadd_4_n17), .CO(intadd_4_n16), .S(intadd_4_SUM_1_) );
  fad1_hd intadd_4_U16 ( .A(intadd_4_A_2_), .B(intadd_4_B_2_), .CI(
        intadd_4_n16), .CO(intadd_4_n15), .S(intadd_4_SUM_2_) );
  fad1_hd intadd_4_U15 ( .A(intadd_4_A_3_), .B(intadd_4_B_3_), .CI(
        intadd_4_n15), .CO(intadd_4_n14), .S(intadd_4_SUM_3_) );
  fad1_hd intadd_4_U14 ( .A(intadd_4_A_4_), .B(intadd_4_B_4_), .CI(
        intadd_4_n14), .CO(intadd_4_n13), .S(intadd_4_SUM_4_) );
  fad1_hd intadd_4_U13 ( .A(intadd_4_A_5_), .B(intadd_4_B_5_), .CI(
        intadd_4_n13), .CO(intadd_4_n12), .S(intadd_4_SUM_5_) );
  fad1_hd intadd_4_U12 ( .A(intadd_4_A_6_), .B(intadd_4_B_6_), .CI(
        intadd_4_n12), .CO(intadd_4_n11), .S(intadd_4_SUM_6_) );
  fad1_hd intadd_4_U11 ( .A(intadd_4_A_7_), .B(intadd_4_B_7_), .CI(
        intadd_4_n11), .CO(intadd_4_n10), .S(intadd_4_SUM_7_) );
  fad1_hd intadd_4_U10 ( .A(intadd_4_A_8_), .B(intadd_4_B_8_), .CI(
        intadd_4_n10), .CO(intadd_4_n9), .S(intadd_4_SUM_8_) );
  fad1_hd intadd_4_U9 ( .A(intadd_4_A_9_), .B(intadd_4_B_9_), .CI(intadd_4_n9), 
        .CO(intadd_4_n8), .S(intadd_4_SUM_9_) );
  fad1_hd intadd_4_U8 ( .A(intadd_4_A_10_), .B(intadd_4_B_10_), .CI(
        intadd_4_n8), .CO(intadd_4_n7), .S(intadd_4_SUM_10_) );
  fad1_hd intadd_4_U7 ( .A(intadd_4_A_11_), .B(intadd_4_B_11_), .CI(
        intadd_4_n7), .CO(intadd_4_n6), .S(intadd_4_SUM_11_) );
  fad1_hd intadd_4_U6 ( .A(intadd_4_A_12_), .B(intadd_4_B_12_), .CI(
        intadd_4_n6), .CO(intadd_4_n5), .S(intadd_4_SUM_12_) );
  fad1_hd intadd_4_U5 ( .A(intadd_4_A_13_), .B(intadd_4_B_13_), .CI(
        intadd_4_n5), .CO(intadd_4_n4), .S(intadd_4_SUM_13_) );
  fad1_hd intadd_4_U4 ( .A(intadd_6_n1), .B(intadd_4_B_14_), .CI(intadd_4_n4), 
        .CO(intadd_4_n3), .S(intadd_4_SUM_14_) );
  fad1_hd intadd_4_U3 ( .A(intadd_19_SUM_0_), .B(intadd_4_B_15_), .CI(
        intadd_4_n3), .CO(intadd_4_n2), .S(intadd_4_SUM_15_) );
  fad1_hd intadd_6_U12 ( .A(intadd_6_A_0_), .B(intadd_6_B_0_), .CI(intadd_6_CI), .CO(intadd_6_n11), .S(intadd_4_A_3_) );
  fad1_hd intadd_6_U11 ( .A(intadd_6_A_1_), .B(intadd_6_B_1_), .CI(
        intadd_6_n11), .CO(intadd_6_n10), .S(intadd_4_A_4_) );
  fad1_hd intadd_6_U10 ( .A(intadd_6_A_2_), .B(intadd_6_B_2_), .CI(
        intadd_6_n10), .CO(intadd_6_n9), .S(intadd_4_A_5_) );
  fad1_hd intadd_6_U9 ( .A(intadd_6_A_3_), .B(intadd_5_SUM_0_), .CI(
        intadd_6_n9), .CO(intadd_6_n8), .S(intadd_4_A_6_) );
  fad1_hd intadd_6_U8 ( .A(intadd_5_SUM_1_), .B(intadd_6_B_4_), .CI(
        intadd_6_n8), .CO(intadd_6_n7), .S(intadd_4_A_7_) );
  fad1_hd intadd_6_U7 ( .A(intadd_6_A_5_), .B(intadd_5_SUM_2_), .CI(
        intadd_6_n7), .CO(intadd_6_n6), .S(intadd_4_A_8_) );
  fad1_hd intadd_6_U6 ( .A(intadd_6_A_6_), .B(intadd_5_SUM_3_), .CI(
        intadd_6_n6), .CO(intadd_6_n5), .S(intadd_4_A_9_) );
  fad1_hd intadd_6_U5 ( .A(intadd_6_A_7_), .B(intadd_5_SUM_4_), .CI(
        intadd_6_n5), .CO(intadd_6_n4), .S(intadd_4_A_10_) );
  fad1_hd intadd_6_U4 ( .A(intadd_6_A_8_), .B(intadd_5_SUM_5_), .CI(
        intadd_6_n4), .CO(intadd_6_n3), .S(intadd_4_A_11_) );
  fad1_hd intadd_6_U3 ( .A(intadd_5_SUM_6_), .B(intadd_6_B_9_), .CI(
        intadd_6_n3), .CO(intadd_6_n2), .S(intadd_4_A_12_) );
  fad1_hd intadd_6_U2 ( .A(intadd_6_A_10_), .B(intadd_5_SUM_7_), .CI(
        intadd_6_n2), .CO(intadd_6_n1), .S(intadd_4_B_13_) );
  fd1qd1_hd b_m_reg_1_ ( .D(n307), .CK(i_CLK), .Q(b_m[1]) );
  fad1_hd intadd_10_U2 ( .A(intadd_10_A_5_), .B(intadd_10_B_5_), .CI(
        intadd_10_n2), .CO(intadd_10_n1), .S(intadd_10_SUM_5_) );
  fad1_hd intadd_17_U2 ( .A(intadd_17_A_2_), .B(intadd_17_B_2_), .CI(
        intadd_17_n2), .CO(intadd_17_n1), .S(intadd_17_SUM_2_) );
  fad1_hd intadd_4_U2 ( .A(intadd_19_SUM_1_), .B(intadd_4_B_16_), .CI(
        intadd_4_n2), .CO(intadd_4_n1), .S(intadd_4_SUM_16_) );
  fad1_hd intadd_15_U2 ( .A(intadd_10_SUM_3_), .B(intadd_15_B_2_), .CI(
        intadd_15_n2), .CO(intadd_15_n1), .S(intadd_15_SUM_2_) );
  fad1_hd intadd_11_U2 ( .A(intadd_11_A_4_), .B(intadd_11_B_4_), .CI(
        intadd_11_n2), .CO(intadd_11_n1), .S(intadd_11_SUM_4_) );
  fad1_hd intadd_16_U2 ( .A(intadd_9_SUM_7_), .B(intadd_16_B_2_), .CI(
        intadd_16_n2), .CO(intadd_16_n1), .S(intadd_16_SUM_2_) );
  fad1_hd intadd_8_U2 ( .A(intadd_8_A_8_), .B(intadd_8_B_8_), .CI(intadd_8_n2), 
        .CO(intadd_8_n1), .S(intadd_8_SUM_8_) );
  fad1_hd intadd_7_U2 ( .A(intadd_7_A_10_), .B(intadd_7_B_10_), .CI(
        intadd_7_n2), .CO(intadd_7_n1), .S(intadd_7_SUM_10_) );
  fad1_hd intadd_14_U4 ( .A(intadd_14_A_0_), .B(intadd_14_B_0_), .CI(
        intadd_14_CI), .CO(intadd_14_n3), .S(intadd_14_SUM_0_) );
  fad1_hd intadd_13_U2 ( .A(intadd_13_A_2_), .B(intadd_13_B_2_), .CI(
        intadd_13_n2), .CO(intadd_13_n1), .S(intadd_13_SUM_2_) );
  fad1_hd intadd_3_U15 ( .A(intadd_3_B_5_), .B(intadd_3_B_4_), .CI(
        intadd_3_n15), .CO(intadd_3_n14), .S(intadd_3_SUM_4_) );
  fad1_hd intadd_3_U16 ( .A(intadd_3_B_4_), .B(intadd_3_B_3_), .CI(
        intadd_3_n16), .CO(intadd_3_n15), .S(intadd_3_SUM_3_) );
  fad1_hd intadd_3_U18 ( .A(intadd_3_B_2_), .B(intadd_3_B_1_), .CI(
        intadd_3_n18), .CO(intadd_3_n17), .S(intadd_3_SUM_1_) );
  fad1_hd intadd_3_U17 ( .A(intadd_3_B_3_), .B(intadd_3_B_2_), .CI(
        intadd_3_n17), .CO(intadd_3_n16), .S(intadd_3_SUM_2_) );
  fad1_hd intadd_3_U19 ( .A(intadd_3_B_1_), .B(intadd_3_B_0_), .CI(intadd_3_CI), .CO(intadd_3_n18), .S(intadd_3_SUM_0_) );
  fad2_hd intadd_0_U14 ( .A(intadd_0_A_24_), .B(intadd_0_B_24_), .CI(
        intadd_0_n14), .CO(intadd_0_n13), .S(N210) );
  fad2_hd intadd_0_U18 ( .A(intadd_0_A_20_), .B(intadd_0_B_20_), .CI(
        intadd_0_n18), .CO(intadd_0_n17), .S(N206) );
  fad1_hd intadd_3_U14 ( .A(intadd_3_B_6_), .B(intadd_3_B_5_), .CI(
        intadd_3_n14), .CO(intadd_3_n13), .S(intadd_3_SUM_5_) );
  fd1qd1_hd sticky_reg ( .D(n283), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd o_Z_STB_reg ( .D(n358), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n350), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd z_reg_30_ ( .D(n230), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n310), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n355), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd round_bit_reg ( .D(n284), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd a_m_reg_13_ ( .D(n336), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n331), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n328), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd z_reg_31_ ( .D(n229), .CK(i_CLK), .Q(z[31]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n308), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd z_reg_21_ ( .D(n239), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n240), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n241), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n242), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_25_ ( .D(n235), .CK(i_CLK), .Q(z[25]) );
  fd1qd1_hd z_reg_22_ ( .D(n238), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n337), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n349), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n335), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n340), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n343), .CK(i_CLK), .Q(a_m[6]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n333), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n341), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n330), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n345), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n329), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n332), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n354), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n347), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n342), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n339), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n346), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n348), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n334), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n338), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n344), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd z_reg_15_ ( .D(n245), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n246), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_11_ ( .D(n249), .CK(i_CLK), .Q(z[11]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n15), .CK(i_CLK), .Q(b[22]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n500), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n15), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n12), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n499), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n9), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n9), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n3), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n475), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n146), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n5), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n501), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n11), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd z_s_reg ( .D(b_s), .E(n490), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd product_reg_2_ ( .D(N176), .E(n490), .CK(i_CLK), .Q(product[2])
         );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n8), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n8), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n7), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n2), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n475), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n3), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n9), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n3), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n11), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n13), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n15), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n13), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n13), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n2), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n2), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n8), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n7), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n3), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n3), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n2), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n9), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n7), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n7), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n2), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n8), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n9), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n9), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n3), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n475), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n8), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n8), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n7), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n2), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1624), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n12), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n146), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n5), .CK(i_CLK), .Q(b[28]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n12), .CK(i_CLK), .Q(b[26]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n4), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n499), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n4), .CK(i_CLK), .Q(b[23]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n13), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n4), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n5), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n501), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n499), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n5), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n501), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n11), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n1), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n13), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n146), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n500), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n13), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n502), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n499), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n15), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n502), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n499), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n501), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n11), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n15), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n5), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n12), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n502), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n4), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n500), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n12), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n502), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n12), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n5), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n500), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n15), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n11), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd guard_reg ( .D(n104), .E(n105), .CK(i_CLK), .Q(net908) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n500), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n4), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n146), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n4), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n502), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd product_reg_3_ ( .D(N177), .E(n487), .CK(i_CLK), .Q(product[3])
         );
  fd1eqd1_hd product_reg_4_ ( .D(N178), .E(n490), .CK(i_CLK), .Q(product[4])
         );
  fd1eqd1_hd product_reg_5_ ( .D(N179), .E(n489), .CK(i_CLK), .Q(product[5])
         );
  fd1eqd1_hd product_reg_6_ ( .D(N180), .E(n491), .CK(i_CLK), .Q(product[6])
         );
  fd1eqd1_hd product_reg_7_ ( .D(N181), .E(n492), .CK(i_CLK), .Q(product[7])
         );
  fd1eqd1_hd product_reg_8_ ( .D(N182), .E(n488), .CK(i_CLK), .Q(product[8])
         );
  fd1eqd1_hd product_reg_9_ ( .D(N183), .E(n488), .CK(i_CLK), .Q(product[9])
         );
  fd1eqd1_hd product_reg_10_ ( .D(N184), .E(n495), .CK(i_CLK), .Q(product[10])
         );
  fd1eqd1_hd z_e_reg_8_ ( .D(N474), .E(n6), .CK(i_CLK), .Q(z_e[8]) );
  fd1eqd1_hd z_e_reg_7_ ( .D(N473), .E(n6), .CK(i_CLK), .Q(z_e[7]) );
  fd1eqd1_hd z_e_reg_6_ ( .D(N472), .E(n6), .CK(i_CLK), .Q(z_e[6]) );
  fd1eqd1_hd z_e_reg_5_ ( .D(N471), .E(n6), .CK(i_CLK), .Q(z_e[5]) );
  fd1eqd1_hd z_e_reg_4_ ( .D(N470), .E(n6), .CK(i_CLK), .Q(z_e[4]) );
  fd1eqd1_hd z_e_reg_3_ ( .D(N469), .E(n3276), .CK(i_CLK), .Q(z_e[3]) );
  fd1eqd1_hd z_e_reg_2_ ( .D(N468), .E(n3276), .CK(i_CLK), .Q(z_e[2]) );
  fd1eqd1_hd z_e_reg_1_ ( .D(N467), .E(n3276), .CK(i_CLK), .Q(z_e[1]) );
  fd1eqd1_hd z_e_reg_0_ ( .D(n3277), .E(n3276), .CK(i_CLK), .Q(z_e[0]) );
  fd1eqd1_hd product_reg_11_ ( .D(N185), .E(n493), .CK(i_CLK), .Q(product[11])
         );
  fd1eqd1_hd z_e_reg_9_ ( .D(N475), .E(n3276), .CK(i_CLK), .Q(z_e[9]) );
  fd1eqd1_hd product_reg_12_ ( .D(N186), .E(n487), .CK(i_CLK), .Q(product[12])
         );
  fd1eqd1_hd product_reg_13_ ( .D(N187), .E(n489), .CK(i_CLK), .Q(product[13])
         );
  fd1eqd1_hd product_reg_14_ ( .D(N188), .E(n494), .CK(i_CLK), .Q(product[14])
         );
  fd1eqd1_hd product_reg_15_ ( .D(N189), .E(n492), .CK(i_CLK), .Q(product[15])
         );
  fd1eqd1_hd product_reg_16_ ( .D(N190), .E(n494), .CK(i_CLK), .Q(product[16])
         );
  fd1eqd1_hd product_reg_17_ ( .D(N191), .E(n490), .CK(i_CLK), .Q(product[17])
         );
  fd1eqd1_hd product_reg_18_ ( .D(N192), .E(n489), .CK(i_CLK), .Q(product[18])
         );
  fd1eqd1_hd product_reg_19_ ( .D(N193), .E(n492), .CK(i_CLK), .Q(product[19])
         );
  fd1eqd1_hd product_reg_20_ ( .D(N194), .E(n493), .CK(i_CLK), .Q(product[20])
         );
  fd1eqd1_hd product_reg_21_ ( .D(N195), .E(n487), .CK(i_CLK), .Q(product[21])
         );
  fd1eqd1_hd product_reg_22_ ( .D(N196), .E(n488), .CK(i_CLK), .Q(product[22])
         );
  fd1eqd1_hd product_reg_23_ ( .D(N197), .E(n491), .CK(i_CLK), .Q(product[23])
         );
  fd1eqd1_hd product_reg_24_ ( .D(N198), .E(n494), .CK(i_CLK), .Q(product[24])
         );
  fd1eqd1_hd product_reg_25_ ( .D(N199), .E(n493), .CK(i_CLK), .Q(product[25])
         );
  fd1eqd1_hd product_reg_26_ ( .D(N200), .E(n489), .CK(i_CLK), .Q(product[26])
         );
  fd1eqd1_hd product_reg_27_ ( .D(N201), .E(n490), .CK(i_CLK), .Q(product[27])
         );
  fd1eqd1_hd product_reg_28_ ( .D(N202), .E(n490), .CK(i_CLK), .Q(product[28])
         );
  fd1eqd1_hd product_reg_29_ ( .D(N203), .E(n491), .CK(i_CLK), .Q(product[29])
         );
  fd1eqd1_hd product_reg_30_ ( .D(N204), .E(n487), .CK(i_CLK), .Q(product[30])
         );
  fd1eqd1_hd product_reg_31_ ( .D(N205), .E(n489), .CK(i_CLK), .Q(product[31])
         );
  fd1eqd1_hd product_reg_32_ ( .D(N206), .E(n494), .CK(i_CLK), .Q(product[32])
         );
  fd1eqd1_hd product_reg_33_ ( .D(N207), .E(n494), .CK(i_CLK), .Q(product[33])
         );
  fd1eqd1_hd product_reg_34_ ( .D(N208), .E(n491), .CK(i_CLK), .Q(product[34])
         );
  fd1eqd1_hd product_reg_35_ ( .D(N209), .E(n488), .CK(i_CLK), .Q(product[35])
         );
  fd1eqd1_hd product_reg_36_ ( .D(N210), .E(n487), .CK(i_CLK), .Q(product[36])
         );
  fd1eqd1_hd product_reg_37_ ( .D(N211), .E(n494), .CK(i_CLK), .Q(product[37])
         );
  fd1eqd1_hd product_reg_38_ ( .D(N212), .E(n492), .CK(i_CLK), .Q(product[38])
         );
  fd1eqd1_hd product_reg_39_ ( .D(N213), .E(n492), .CK(i_CLK), .Q(product[39])
         );
  fd1eqd1_hd product_reg_40_ ( .D(N214), .E(n488), .CK(i_CLK), .Q(product[40])
         );
  fd1eqd1_hd product_reg_41_ ( .D(N215), .E(n492), .CK(i_CLK), .Q(product[41])
         );
  fd1eqd1_hd product_reg_42_ ( .D(N216), .E(n493), .CK(i_CLK), .Q(product[42])
         );
  fd1eqd1_hd product_reg_43_ ( .D(N217), .E(n493), .CK(i_CLK), .Q(product[43])
         );
  fd1eqd1_hd product_reg_44_ ( .D(N218), .E(n489), .CK(i_CLK), .Q(product[44])
         );
  fd1eqd1_hd product_reg_45_ ( .D(N219), .E(n488), .CK(i_CLK), .Q(product[45])
         );
  fd1eqd1_hd product_reg_46_ ( .D(N220), .E(n491), .CK(i_CLK), .Q(product[46])
         );
  fd1eqd1_hd product_reg_47_ ( .D(N221), .E(n493), .CK(i_CLK), .Q(product[47])
         );
  fd1eqd1_hd product_reg_48_ ( .D(N222), .E(n491), .CK(i_CLK), .Q(product[48])
         );
  fd1eqd1_hd product_reg_49_ ( .D(N223), .E(n487), .CK(i_CLK), .Q(product[49])
         );
  fad1_hd intadd_3_U2 ( .A(intadd_3_A_17_), .B(intadd_3_B_17_), .CI(
        intadd_3_n2), .CO(intadd_3_n1), .S(intadd_3_SUM_17_) );
  fad1_hd intadd_3_U5 ( .A(intadd_3_B_15_), .B(b_m[17]), .CI(intadd_3_n5), 
        .CO(intadd_3_n4), .S(intadd_3_SUM_14_) );
  fad1_hd intadd_3_U8 ( .A(intadd_3_B_12_), .B(intadd_3_B_11_), .CI(
        intadd_3_n8), .CO(intadd_3_n7), .S(intadd_3_SUM_11_) );
  fad1_hd intadd_3_U12 ( .A(intadd_3_B_8_), .B(intadd_3_B_7_), .CI(
        intadd_3_n12), .CO(intadd_3_n11), .S(intadd_3_SUM_7_) );
  fad1_hd intadd_3_U9 ( .A(intadd_3_B_11_), .B(intadd_3_B_10_), .CI(
        intadd_3_n9), .CO(intadd_3_n8), .S(intadd_3_SUM_10_) );
  fad1_hd intadd_3_U10 ( .A(intadd_3_B_10_), .B(intadd_3_B_9_), .CI(
        intadd_3_n10), .CO(intadd_3_n9), .S(intadd_3_SUM_9_) );
  fad1_hd intadd_3_U11 ( .A(intadd_3_B_9_), .B(intadd_3_B_8_), .CI(
        intadd_3_n11), .CO(intadd_3_n10), .S(intadd_3_SUM_8_) );
  fad1_hd intadd_3_U13 ( .A(intadd_3_B_7_), .B(intadd_3_B_6_), .CI(
        intadd_3_n13), .CO(intadd_3_n12), .S(intadd_3_SUM_6_) );
  fad1_hd intadd_3_U4 ( .A(intadd_3_B_16_), .B(intadd_3_B_15_), .CI(
        intadd_3_n4), .CO(intadd_3_n3), .S(intadd_3_SUM_15_) );
  fad1_hd intadd_3_U3 ( .A(intadd_3_B_17_), .B(intadd_3_B_16_), .CI(
        intadd_3_n3), .CO(intadd_3_n2), .S(intadd_3_SUM_16_) );
  fad1_hd intadd_3_U7 ( .A(intadd_3_B_13_), .B(intadd_3_B_12_), .CI(
        intadd_3_n7), .CO(intadd_3_n6), .S(intadd_3_SUM_12_) );
  fad1_hd intadd_3_U6 ( .A(b_m[17]), .B(intadd_3_B_13_), .CI(intadd_3_n6), 
        .CO(intadd_3_n5), .S(intadd_3_SUM_13_) );
  fad1_hd intadd_0_U17 ( .A(intadd_0_A_21_), .B(intadd_0_B_21_), .CI(
        intadd_0_n17), .CO(intadd_0_n16), .S(N207) );
  fad1_hd intadd_0_U13 ( .A(intadd_8_SUM_8_), .B(intadd_0_B_25_), .CI(
        intadd_0_n13), .CO(intadd_0_n12), .S(N211) );
  fad1_hd intadd_0_U7 ( .A(intadd_0_A_31_), .B(intadd_0_B_31_), .CI(
        intadd_0_n7), .CO(intadd_0_n6), .S(N217) );
  fad4_hd intadd_0_U15 ( .A(intadd_0_A_23_), .B(intadd_7_n1), .CI(intadd_0_n15), .CO(intadd_0_n14), .S(N209) );
  fad4_hd intadd_0_U9 ( .A(intadd_0_A_29_), .B(intadd_11_n1), .CI(intadd_0_n9), 
        .CO(intadd_0_n8), .S(N215) );
  fad1_hd intadd_0_U6 ( .A(intadd_13_SUM_2_), .B(intadd_0_B_32_), .CI(
        intadd_0_n6), .CO(intadd_0_n5), .S(N218) );
  fad1_hd intadd_0_U8 ( .A(intadd_0_A_30_), .B(intadd_0_B_30_), .CI(
        intadd_0_n8), .CO(intadd_0_n7), .S(N216) );
  fad1_hd intadd_0_U5 ( .A(intadd_0_A_33_), .B(intadd_13_n1), .CI(intadd_0_n5), 
        .CO(intadd_0_n4), .S(N219) );
  fad2_hd intadd_2_U17 ( .A(intadd_2_A_3_), .B(intadd_2_B_3_), .CI(
        intadd_2_n17), .CO(intadd_2_n16), .S(intadd_1_A_6_) );
  fad2_hd intadd_2_U7 ( .A(intadd_2_A_13_), .B(intadd_2_B_13_), .CI(
        intadd_2_n7), .CO(intadd_2_n6), .S(intadd_1_A_16_) );
  fad2_hd intadd_0_U16 ( .A(intadd_7_SUM_10_), .B(intadd_0_B_22_), .CI(
        intadd_0_n16), .CO(intadd_0_n15), .S(N208) );
  fad2_hd intadd_0_U19 ( .A(intadd_0_A_19_), .B(intadd_0_B_19_), .CI(
        intadd_0_n19), .CO(intadd_0_n18), .S(N205) );
  fad2_hd intadd_0_U20 ( .A(intadd_0_A_18_), .B(intadd_0_B_18_), .CI(
        intadd_0_n20), .CO(intadd_0_n19), .S(N204) );
  fad2_hd intadd_2_U18 ( .A(intadd_2_A_2_), .B(intadd_2_B_2_), .CI(
        intadd_2_n18), .CO(intadd_2_n17), .S(intadd_1_B_5_) );
  fad2_hd U367 ( .A(intadd_11_SUM_4_), .B(intadd_0_B_28_), .CI(intadd_0_n10), 
        .CO(intadd_0_n9), .S(N214) );
  fad2_hd U368 ( .A(intadd_2_A_17_), .B(intadd_2_B_17_), .CI(intadd_2_n3), 
        .CO(intadd_2_n2), .S(intadd_1_A_20_) );
  ivd1_hd U369 ( .A(intadd_3_n1), .Y(n822) );
  ivd1_hd U370 ( .A(n86), .Y(n1391) );
  ivd1_hd U371 ( .A(a_m[8]), .Y(n609) );
  fad1_hd U372 ( .A(intadd_2_A_18_), .B(intadd_2_B_18_), .CI(intadd_2_n2), 
        .CO(intadd_2_n1), .S(intadd_1_B_21_) );
  fad1_hd U373 ( .A(intadd_2_A_12_), .B(intadd_2_B_12_), .CI(intadd_2_n8), 
        .CO(intadd_2_n7), .S(intadd_1_B_15_) );
  fad1_hd U374 ( .A(intadd_2_A_4_), .B(intadd_2_B_4_), .CI(intadd_2_n16), .CO(
        intadd_2_n15), .S(intadd_1_A_7_) );
  ivd1_hd U375 ( .A(a_m[5]), .Y(n85) );
  fad1_hd U376 ( .A(intadd_0_A_34_), .B(intadd_0_B_34_), .CI(intadd_0_n4), 
        .CO(intadd_0_n3), .S(N220) );
  clknd2d1_hd U377 ( .A(n744), .B(n745), .Y(n757) );
  clknd2d1_hd U378 ( .A(n701), .B(n700), .Y(n711) );
  ivd1_hd U379 ( .A(n92), .Y(n1369) );
  nid1_hd U380 ( .A(n399), .Y(n397) );
  clknd2d1_hd U381 ( .A(n666), .B(n667), .Y(n676) );
  nid1_hd U382 ( .A(n1391), .Y(n468) );
  nid1_hd U383 ( .A(n384), .Y(n386) );
  nid1_hd U384 ( .A(n850), .Y(n388) );
  nid1_hd U385 ( .A(n470), .Y(n472) );
  clknd2d1_hd U386 ( .A(n635), .B(n634), .Y(n636) );
  clknd2d1_hd U387 ( .A(n1069), .B(n1072), .Y(n1068) );
  clknd2d1_hd U388 ( .A(a_m[23]), .B(n119), .Y(n856) );
  clknd2d1_hd U389 ( .A(n814), .B(n815), .Y(n832) );
  clknd2d1_hd U390 ( .A(n205), .B(n778), .Y(n776) );
  clknd2d1_hd U391 ( .A(n203), .B(n775), .Y(n777) );
  clknd2d1_hd U392 ( .A(n619), .B(intadd_3_B_5_), .Y(n940) );
  clknd2d1_hd U393 ( .A(n619), .B(intadd_3_B_3_), .Y(intadd_9_B_2_) );
  nid1_hd U394 ( .A(n447), .Y(n445) );
  clknd2d1_hd U395 ( .A(n619), .B(intadd_3_B_2_), .Y(intadd_9_CI) );
  clknd2d1_hd U396 ( .A(n619), .B(n504), .Y(n886) );
  clknd2d1_hd U397 ( .A(n117), .B(n809), .Y(n813) );
  clknd2d1_hd U398 ( .A(n790), .B(n789), .Y(n808) );
  nid1_hd U399 ( .A(n428), .Y(n430) );
  nid1_hd U400 ( .A(n459), .Y(n461) );
  clknd2d1_hd U401 ( .A(a_m[23]), .B(n536), .Y(intadd_11_A_0_) );
  nid1_hd U402 ( .A(n1040), .Y(n438) );
  clknd2d1_hd U403 ( .A(n119), .B(n773), .Y(n775) );
  nid1_hd U404 ( .A(n420), .Y(n422) );
  clknd2d1_hd U405 ( .A(n111), .B(n718), .Y(n716) );
  clknd2d1_hd U406 ( .A(n110), .B(n715), .Y(n717) );
  clknd2d1_hd U407 ( .A(n620), .B(intadd_3_B_11_), .Y(n998) );
  nid1_hd U408 ( .A(n440), .Y(n442) );
  clknd2d1_hd U409 ( .A(n619), .B(intadd_3_B_9_), .Y(intadd_10_B_1_) );
  nid1_hd U410 ( .A(n1039), .Y(n433) );
  nid1_hd U411 ( .A(n438), .Y(n437) );
  nid1_hd U412 ( .A(n424), .Y(n425) );
  clknd2d1_hd U413 ( .A(n757), .B(n747), .Y(intadd_6_CI) );
  clknd2d1_hd U414 ( .A(n729), .B(n728), .Y(n740) );
  nid1_hd U415 ( .A(n966), .Y(n409) );
  nid1_hd U416 ( .A(n415), .Y(n414) );
  clknd2d1_hd U417 ( .A(n620), .B(n574), .Y(n1025) );
  nid1_hd U418 ( .A(n440), .Y(n441) );
  nid1_hd U419 ( .A(n1062), .Y(n440) );
  nid1_hd U420 ( .A(n447), .Y(n446) );
  nid1_hd U421 ( .A(n1039), .Y(n434) );
  nid1_hd U422 ( .A(n424), .Y(n426) );
  nid1_hd U423 ( .A(n416), .Y(n418) );
  nid1_hd U424 ( .A(n408), .Y(n410) );
  nid1_hd U425 ( .A(n1380), .Y(n465) );
  nid1_hd U426 ( .A(n416), .Y(n417) );
  nid1_hd U427 ( .A(n532), .Y(n534) );
  clknd2d1_hd U428 ( .A(n117), .B(n713), .Y(n715) );
  nid1_hd U429 ( .A(n400), .Y(n403) );
  clknd2d1_hd U430 ( .A(a_m[11]), .B(n691), .Y(n685) );
  clknd2d1_hd U431 ( .A(a_m[11]), .B(n688), .Y(n686) );
  nid1_hd U432 ( .A(n407), .Y(n405) );
  nid1_hd U433 ( .A(n620), .Y(n619) );
  clknd2d1_hd U434 ( .A(n620), .B(intadd_3_B_17_), .Y(n1044) );
  nid1_hd U435 ( .A(n440), .Y(n443) );
  nid1_hd U436 ( .A(n1064), .Y(n447) );
  clknd2d1_hd U437 ( .A(n620), .B(intadd_3_B_15_), .Y(intadd_14_B_1_) );
  clknd2d1_hd U438 ( .A(intadd_13_A_0_), .B(n1025), .Y(n1033) );
  clknd2d1_hd U439 ( .A(n785), .B(n773), .Y(n784) );
  nid1_hd U440 ( .A(n1040), .Y(n439) );
  nid1_hd U441 ( .A(n428), .Y(n431) );
  clknd2d1_hd U442 ( .A(n724), .B(n713), .Y(n723) );
  nid1_hd U443 ( .A(n1020), .Y(n428) );
  nid1_hd U444 ( .A(n967), .Y(n415) );
  clknd2d1_hd U445 ( .A(n696), .B(n683), .Y(n695) );
  nid1_hd U446 ( .A(n420), .Y(n423) );
  nid1_hd U447 ( .A(b_m[18]), .Y(n580) );
  nid1_hd U448 ( .A(n966), .Y(n408) );
  nid1_hd U449 ( .A(n935), .Y(n407) );
  nid1_hd U450 ( .A(n415), .Y(n413) );
  nid1_hd U451 ( .A(n465), .Y(n464) );
  nid1_hd U452 ( .A(n400), .Y(n402) );
  nr2bd1_hd U453 ( .AN(n673), .B(n674), .Y(n935) );
  ad3d1_hd U454 ( .A(n654), .B(n653), .C(n652), .Y(n906) );
  scg2d1_hd U455 ( .A(n1112), .B(n76), .C(n75), .D(n200), .Y(n1053) );
  nid1_hd U456 ( .A(n591), .Y(n590) );
  scg2d1_hd U457 ( .A(n1066), .B(intadd_3_n1), .C(n822), .D(n802), .Y(n1037)
         );
  nid1_hd U458 ( .A(n574), .Y(n577) );
  nid1_hd U459 ( .A(n906), .Y(n392) );
  nid1_hd U460 ( .A(n1391), .Y(n469) );
  nid1_hd U461 ( .A(n564), .Y(n562) );
  nid1_hd U462 ( .A(n907), .Y(n399) );
  clknd2d1_hd U463 ( .A(n119), .B(n683), .Y(n691) );
  nid1_hd U464 ( .A(n523), .Y(n525) );
  nid1_hd U465 ( .A(n519), .Y(n520) );
  nid1_hd U466 ( .A(n392), .Y(n393) );
  nid1_hd U467 ( .A(n399), .Y(n398) );
  nid1_hd U468 ( .A(n468), .Y(n467) );
  clknd2d1_hd U469 ( .A(n642), .B(a_m[5]), .Y(n645) );
  ivd1_hd U470 ( .A(a_m[11]), .Y(n1380) );
  nid1_hd U471 ( .A(n1369), .Y(n459) );
  nid1_hd U472 ( .A(b_m[5]), .Y(n519) );
  nid1_hd U473 ( .A(a_m[23]), .Y(n620) );
  nid1_hd U474 ( .A(n447), .Y(n444) );
  ad3d1_hd U475 ( .A(n829), .B(n828), .C(n827), .Y(n1062) );
  nid1_hd U476 ( .A(n432), .Y(n435) );
  nid1_hd U477 ( .A(n1039), .Y(n432) );
  nid1_hd U478 ( .A(n439), .Y(n436) );
  nid1_hd U479 ( .A(n1019), .Y(n424) );
  ivd1_hd U480 ( .A(n1053), .Y(n58) );
  clknd2d1_hd U481 ( .A(n755), .B(n753), .Y(n1012) );
  nid1_hd U482 ( .A(n1020), .Y(n429) );
  nid1_hd U483 ( .A(n1019), .Y(n427) );
  nid1_hd U484 ( .A(n992), .Y(n416) );
  nid1_hd U485 ( .A(n993), .Y(n421) );
  nid1_hd U486 ( .A(n992), .Y(n419) );
  clknd2d1_hd U487 ( .A(intadd_3_A_17_), .B(intadd_3_n1), .Y(n821) );
  nid1_hd U488 ( .A(n415), .Y(n412) );
  nid1_hd U489 ( .A(n966), .Y(n411) );
  nid1_hd U490 ( .A(n466), .Y(n463) );
  clknd2d1_hd U491 ( .A(n674), .B(n672), .Y(n927) );
  nid1_hd U492 ( .A(n399), .Y(n396) );
  nid1_hd U493 ( .A(n392), .Y(n395) );
  nid1_hd U494 ( .A(n935), .Y(n404) );
  nid1_hd U495 ( .A(n934), .Y(n401) );
  ivd1_hd U496 ( .A(n1053), .Y(n57) );
  nid1_hd U497 ( .A(n588), .Y(n589) );
  nid1_hd U498 ( .A(n579), .Y(n581) );
  nid1_hd U499 ( .A(n574), .Y(n575) );
  nid1_hd U500 ( .A(n574), .Y(n576) );
  nid1_hd U501 ( .A(n1397), .Y(n470) );
  nid1_hd U502 ( .A(b_m[14]), .Y(n561) );
  nid1_hd U503 ( .A(n555), .Y(n553) );
  clknd2d1_hd U504 ( .A(n196), .B(n1399), .Y(n632) );
  nid1_hd U505 ( .A(n470), .Y(n473) );
  nid1_hd U506 ( .A(n391), .Y(n390) );
  nid1_hd U507 ( .A(n532), .Y(n533) );
  nid1_hd U508 ( .A(n523), .Y(n524) );
  clknd2d1_hd U509 ( .A(n676), .B(n669), .Y(intadd_2_CI) );
  nid1_hd U510 ( .A(n384), .Y(n387) );
  nid1_hd U511 ( .A(n1397), .Y(n474) );
  clknd2d1_hd U512 ( .A(n118), .B(n643), .Y(n642) );
  nid1_hd U513 ( .A(n388), .Y(n391) );
  nid1_hd U514 ( .A(n849), .Y(n385) );
  clknd2d1_hd U515 ( .A(n1401), .B(a_m[1]), .Y(n847) );
  clknd2d1_hd U516 ( .A(a_m[0]), .B(n623), .Y(n630) );
  nid1_hd U517 ( .A(n850), .Y(n389) );
  clknd2d1_hd U518 ( .A(state[2]), .B(n1116), .Y(n622) );
  nid1_hd U519 ( .A(n609), .Y(n607) );
  clknd2d1_hd U520 ( .A(n1408), .B(n1126), .Y(n1127) );
  clknd2d1_hd U521 ( .A(n1340), .B(n1128), .Y(n1125) );
  clknd2d1_hd U522 ( .A(n1267), .B(n105), .Y(n1256) );
  clknd2d1_hd U523 ( .A(n1294), .B(n1419), .Y(n1266) );
  nid1_hd U524 ( .A(b_m[8]), .Y(n532) );
  nid1_hd U525 ( .A(n514), .Y(n513) );
  ivd1_hd U526 ( .A(b_m[7]), .Y(n531) );
  nid1_hd U527 ( .A(n519), .Y(n522) );
  nid1_hd U528 ( .A(b_m[6]), .Y(n523) );
  nid1_hd U529 ( .A(b_m[14]), .Y(n564) );
  nid1_hd U530 ( .A(b_m[12]), .Y(n552) );
  nid1_hd U531 ( .A(n552), .Y(n555) );
  nid1_hd U532 ( .A(b_m[17]), .Y(n574) );
  nid1_hd U533 ( .A(b_m[18]), .Y(n579) );
  nid1_hd U534 ( .A(n588), .Y(n591) );
  ivd1_hd U535 ( .A(b_m[21]), .Y(n597) );
  clknd2d1_hd U536 ( .A(n1121), .B(n1087), .Y(n1138) );
  nid1_hd U537 ( .A(n484), .Y(n482) );
  nid1_hd U538 ( .A(n621), .Y(n616) );
  clknd2d1_hd U539 ( .A(n1628), .B(state[3]), .Y(n1124) );
  clknd2d1_hd U540 ( .A(state[3]), .B(n1111), .Y(n1115) );
  nid1_hd U541 ( .A(n616), .Y(n617) );
  clknd2d1_hd U542 ( .A(intadd_3_A_17_), .B(n107), .Y(n1074) );
  clknd2d1_hd U543 ( .A(n620), .B(n1066), .Y(n1069) );
  clknd2d1_hd U544 ( .A(a_m[23]), .B(n1067), .Y(n1070) );
  clknd2d1_hd U545 ( .A(n656), .B(n648), .Y(intadd_1_A_0_) );
  clknd2d1_hd U546 ( .A(n642), .B(n636), .Y(n641) );
  clknd2d1_hd U547 ( .A(n640), .B(n641), .Y(intadd_1_CI) );
  nid1_hd U548 ( .A(n497), .Y(n498) );
  clknd2d1_hd U549 ( .A(n197), .B(n627), .Y(n625) );
  clknd2d1_hd U550 ( .A(n197), .B(n629), .Y(n626) );
  clknd2d1_hd U551 ( .A(a_m[0]), .B(n118), .Y(n627) );
  nid1_hd U553 ( .A(n1397), .Y(n471) );
  ivd1_hd U554 ( .A(n91), .Y(n92) );
  nid1_hd U555 ( .A(a_m[20]), .Y(n203) );
  nid1_hd U556 ( .A(n1332), .Y(n485) );
  ivd1_hd U557 ( .A(n608), .Y(n604) );
  nid1_hd U558 ( .A(n607), .Y(n608) );
  nid1_hd U559 ( .A(n486), .Y(n476) );
  nid1_hd U560 ( .A(n484), .Y(n483) );
  nid1_hd U561 ( .A(n466), .Y(n462) );
  nid1_hd U562 ( .A(n486), .Y(n477) );
  clknd2d1_hd U563 ( .A(n1174), .B(n1173), .Y(n1177) );
  clknd2d1_hd U564 ( .A(n1126), .B(n1125), .Y(n1131) );
  clknd2d1_hd U565 ( .A(n1128), .B(n1127), .Y(n1129) );
  nid1_hd U566 ( .A(n459), .Y(n460) );
  clknd2d1_hd U567 ( .A(n380), .B(n162), .Y(n1377) );
  ivd1_hd U568 ( .A(n602), .Y(n598) );
  clknd2d1_hd U569 ( .A(state[1]), .B(n1114), .Y(n1292) );
  nid1_hd U570 ( .A(n1303), .Y(n455) );
  clknd2d1_hd U571 ( .A(n1276), .B(n1258), .Y(n1262) );
  clknd2d1_hd U572 ( .A(n199), .B(n1240), .Y(n1244) );
  clknd2d1_hd U573 ( .A(n1276), .B(n1196), .Y(n1200) );
  clknd2d1_hd U574 ( .A(n198), .B(n1223), .Y(n1227) );
  clknd2d1_hd U575 ( .A(n199), .B(n1232), .Y(n1238) );
  clknd2d1_hd U576 ( .A(n198), .B(n1205), .Y(n1220) );
  clknd2d1_hd U577 ( .A(n199), .B(n1269), .Y(n1275) );
  clknd2d1_hd U578 ( .A(n1276), .B(n1187), .Y(n1194) );
  clknd2d1_hd U579 ( .A(n198), .B(n1249), .Y(n1255) );
  nid1_hd U580 ( .A(n1303), .Y(n457) );
  nid1_hd U581 ( .A(n455), .Y(n456) );
  nid1_hd U582 ( .A(n455), .Y(n458) );
  ivd1_hd U583 ( .A(n586), .Y(intadd_3_B_16_) );
  nid1_hd U584 ( .A(b_m[20]), .Y(n588) );
  nid1_hd U585 ( .A(n532), .Y(n535) );
  ivd1_hd U586 ( .A(n530), .Y(intadd_3_B_4_) );
  nid1_hd U587 ( .A(n522), .Y(n521) );
  ivd1_hd U588 ( .A(n518), .Y(intadd_3_B_1_) );
  nid1_hd U589 ( .A(n564), .Y(intadd_3_B_11_) );
  nid1_hd U590 ( .A(n569), .Y(n568) );
  ivd1_hd U591 ( .A(n513), .Y(intadd_3_B_0_) );
  nid1_hd U592 ( .A(n603), .Y(n602) );
  ivd1_hd U593 ( .A(n596), .Y(intadd_3_A_17_) );
  nid1_hd U594 ( .A(n484), .Y(n481) );
  nid1_hd U595 ( .A(b_m[6]), .Y(intadd_3_B_3_) );
  nid1_hd U596 ( .A(n531), .Y(n530) );
  nid1_hd U597 ( .A(n522), .Y(intadd_3_B_2_) );
  nid1_hd U598 ( .A(n523), .Y(n526) );
  ivd1_hd U599 ( .A(n540), .Y(intadd_3_B_6_) );
  ivd1_hd U600 ( .A(n545), .Y(intadd_3_B_7_) );
  nid1_hd U601 ( .A(n551), .Y(n550) );
  nid1_hd U602 ( .A(b_m[18]), .Y(intadd_3_B_15_) );
  nid1_hd U603 ( .A(n587), .Y(n586) );
  clknd2d1_hd U604 ( .A(n1152), .B(n1149), .Y(n1148) );
  clknd2d1_hd U605 ( .A(n1167), .B(n1163), .Y(n1162) );
  clknd2d1_hd U606 ( .A(n1159), .B(n1156), .Y(n1155) );
  ivd1_hd U607 ( .A(n559), .Y(intadd_3_B_10_) );
  nid1_hd U608 ( .A(n564), .Y(n563) );
  ivd1_hd U609 ( .A(n508), .Y(n503) );
  nid1_hd U610 ( .A(b_m[8]), .Y(intadd_3_B_5_) );
  nid1_hd U611 ( .A(n541), .Y(n540) );
  nid1_hd U612 ( .A(n485), .Y(n478) );
  nid1_hd U613 ( .A(n552), .Y(n554) );
  ivd1_hd U614 ( .A(n550), .Y(intadd_3_B_8_) );
  nid1_hd U615 ( .A(n555), .Y(intadd_3_B_9_) );
  nid1_hd U616 ( .A(n560), .Y(n559) );
  nid1_hd U617 ( .A(n485), .Y(n479) );
  ivd1_hd U618 ( .A(n568), .Y(intadd_3_B_12_) );
  ivd1_hd U619 ( .A(n573), .Y(intadd_3_B_13_) );
  nid1_hd U620 ( .A(n574), .Y(n578) );
  nid1_hd U621 ( .A(n579), .Y(n582) );
  nid1_hd U622 ( .A(n485), .Y(n480) );
  nid1_hd U623 ( .A(n509), .Y(n508) );
  nid1_hd U624 ( .A(n591), .Y(intadd_3_B_17_) );
  nid1_hd U625 ( .A(n597), .Y(n596) );
  nid1_hd U626 ( .A(n1332), .Y(n486) );
  clknd2d1_hd U627 ( .A(n1114), .B(n73), .Y(n1409) );
  clknd2d1_hd U628 ( .A(n1116), .B(n1087), .Y(n1349) );
  clknd2d1_hd U629 ( .A(n1085), .B(n1084), .Y(n1141) );
  clknd2d1_hd U630 ( .A(z_e[7]), .B(z_e[8]), .Y(n1140) );
  clknd2d1_hd U631 ( .A(n74), .B(n1120), .Y(n1183) );
  nid1_hd U632 ( .A(n616), .Y(n618) );
  clknd2d1_hd U633 ( .A(state[1]), .B(n1120), .Y(n1143) );
  xo2d1_hd U634 ( .A(intadd_0_n1), .B(n1077), .Y(N223) );
  fad1_hd U635 ( .A(intadd_0_A_35_), .B(intadd_0_B_35_), .CI(intadd_0_n3), 
        .CO(intadd_0_n2), .S(N221) );
  fad1_hd U636 ( .A(intadd_0_A_27_), .B(intadd_0_B_27_), .CI(intadd_0_n11), 
        .CO(intadd_0_n10), .S(N213) );
  fad1_hd U637 ( .A(intadd_0_A_17_), .B(intadd_0_B_17_), .CI(intadd_0_n21), 
        .CO(intadd_0_n20), .S(N203) );
  ivd1_hd U638 ( .A(intadd_1_n1), .Y(intadd_0_A_17_) );
  clknd2d1_hd U639 ( .A(z_m[23]), .B(n1416), .Y(n1418) );
  clknd2d1_hd U640 ( .A(n1417), .B(n1292), .Y(n105) );
  nid1_hd U641 ( .A(n499), .Y(n502) );
  nid1_hd U642 ( .A(n1), .Y(n4) );
  nid1_hd U643 ( .A(n1), .Y(n13) );
  nid1_hd U644 ( .A(n1), .Y(n5) );
  nid1_hd U645 ( .A(n11), .Y(n499) );
  nid1_hd U646 ( .A(n1), .Y(n12) );
  nid1_hd U647 ( .A(n1), .Y(n15) );
  clknd2d1_hd U648 ( .A(n191), .B(n1166), .Y(n235) );
  clknd2d1_hd U649 ( .A(n454), .B(n1135), .Y(n1136) );
  clknd2d1_hd U650 ( .A(z_e[7]), .B(n1148), .Y(n1146) );
  clknd2d1_hd U651 ( .A(n1345), .B(n138), .Y(n311) );
  clknd2d1_hd U652 ( .A(n1360), .B(n148), .Y(n320) );
  clknd2d1_hd U653 ( .A(n1277), .B(n195), .Y(n1278) );
  clknd2d1_hd U654 ( .A(n1281), .B(n1280), .Y(n1279) );
  clknd2d1_hd U655 ( .A(n1302), .B(n1280), .Y(n1283) );
  clknd2d1_hd U656 ( .A(n1346), .B(n138), .Y(n317) );
  clknd2d1_hd U657 ( .A(n1361), .B(n148), .Y(n326) );
  clknd2d1_hd U658 ( .A(n191), .B(n1158), .Y(n233) );
  clknd2d1_hd U659 ( .A(n452), .B(z[23]), .Y(n1170) );
  clknd2d1_hd U660 ( .A(n452), .B(z[24]), .Y(n1168) );
  clknd2d1_hd U661 ( .A(n191), .B(n1151), .Y(n231) );
  clknd2d1_hd U662 ( .A(n452), .B(z[26]), .Y(n1160) );
  clknd2d1_hd U663 ( .A(n452), .B(z[28]), .Y(n1153) );
  clknd2d1_hd U664 ( .A(n1413), .B(n1412), .Y(n1410) );
  clknd2d1_hd U665 ( .A(n1353), .B(n1352), .Y(n1350) );
  clknd2d1_hd U666 ( .A(n1134), .B(n1362), .Y(n148) );
  clknd2d1_hd U667 ( .A(n1134), .B(n1347), .Y(n138) );
  nid1_hd U668 ( .A(n7), .Y(n475) );
  nid1_hd U669 ( .A(n501), .Y(n500) );
  clknd2d1_hd U670 ( .A(n1116), .B(n74), .Y(n1117) );
  nid1_hd U671 ( .A(n502), .Y(n501) );
  clknd2d1_hd U672 ( .A(n1121), .B(n1111), .Y(n155) );
  ivd1_hd U673 ( .A(n75), .Y(n76) );
  ivd1_hd U674 ( .A(n1063), .Y(n75) );
  nid1_hd U675 ( .A(n146), .Y(n1) );
  scg12d1_hd U676 ( .A(o_AB_ACK), .B(i_AB_STB), .C(n155), .Y(n146) );
  ivd1_hd U677 ( .A(n3278), .Y(n2) );
  ivd1_hd U678 ( .A(n3278), .Y(n3) );
  nid1_hd U679 ( .A(n3276), .Y(n6) );
  or3d1_hd U680 ( .A(n73), .B(n1124), .C(n1629), .Y(n3278) );
  ivd1_hd U681 ( .A(n3278), .Y(n7) );
  ivd1_hd U682 ( .A(n3278), .Y(n8) );
  ivd1_hd U683 ( .A(n3278), .Y(n9) );
  nid1_hd U684 ( .A(n146), .Y(n11) );
  fad1_hd U685 ( .A(intadd_0_A_36_), .B(intadd_0_B_36_), .CI(intadd_0_n2), 
        .CO(intadd_0_n1), .S(N222) );
  ivd1_hd U686 ( .A(n1046), .Y(n59) );
  fad1_hd U687 ( .A(n108), .B(n598), .CI(n845), .CO(n1063), .S(n1046) );
  ivd1_hd U688 ( .A(intadd_3_SUM_17_), .Y(n61) );
  ivd1_hd U689 ( .A(intadd_3_SUM_16_), .Y(n63) );
  ivd1_hd U690 ( .A(intadd_3_SUM_15_), .Y(n55) );
  nr2d1_hd U691 ( .A(n657), .B(n656), .Y(n662) );
  ad2d1_hd U692 ( .A(n828), .B(n809), .Y(n1064) );
  ivd1_hd U693 ( .A(b_m[13]), .Y(n560) );
  ivd1_hd U694 ( .A(b_m[9]), .Y(n541) );
  ivd1_hd U695 ( .A(b_m[11]), .Y(n551) );
  nid1_hd U696 ( .A(a_m[23]), .Y(n621) );
  xo2d1_hd U697 ( .A(n472), .B(n848), .Y(intadd_1_B_20_) );
  fad1_hd U698 ( .A(n949), .B(n948), .CI(n947), .CO(n950), .S(n938) );
  xo2d1_hd U699 ( .A(n472), .B(n823), .Y(intadd_1_A_19_) );
  xo2d1_hd U700 ( .A(n1391), .B(n863), .Y(intadd_2_B_18_) );
  ivd1_hd U701 ( .A(n59), .Y(n60) );
  xo2d1_hd U702 ( .A(n472), .B(n803), .Y(intadd_1_A_18_) );
  xo2d1_hd U703 ( .A(n474), .B(n795), .Y(intadd_1_A_17_) );
  xo2d1_hd U704 ( .A(n85), .B(n844), .Y(intadd_2_B_17_) );
  xo2d1_hd U705 ( .A(n472), .B(n794), .Y(intadd_1_B_16_) );
  ivd1_hd U706 ( .A(n1037), .Y(n66) );
  ivd1_hd U707 ( .A(n1037), .Y(n65) );
  ivd1_hd U708 ( .A(n61), .Y(n62) );
  ao22d1_hd U709 ( .A(n596), .B(n822), .C(n602), .D(n821), .Y(n845) );
  xo2d1_hd U710 ( .A(n464), .B(n881), .Y(n904) );
  ivd1_hd U711 ( .A(n63), .Y(n64) );
  ivd1_hd U712 ( .A(n55), .Y(n56) );
  xo2d1_hd U713 ( .A(n465), .B(n868), .Y(intadd_6_A_10_) );
  xo2d1_hd U714 ( .A(n465), .B(n862), .Y(intadd_4_B_12_) );
  xo2d1_hd U715 ( .A(n474), .B(n749), .Y(intadd_1_B_12_) );
  xo2d1_hd U716 ( .A(n469), .B(n781), .Y(intadd_2_B_12_) );
  ivd1_hd U717 ( .A(intadd_3_SUM_14_), .Y(n53) );
  xo2d1_hd U718 ( .A(n465), .B(n843), .Y(intadd_4_B_11_) );
  ivd1_hd U719 ( .A(intadd_3_SUM_13_), .Y(n51) );
  xo2d1_hd U720 ( .A(n465), .B(n835), .Y(intadd_4_B_10_) );
  ivd1_hd U721 ( .A(intadd_3_SUM_12_), .Y(n47) );
  ivd1_hd U722 ( .A(intadd_3_SUM_11_), .Y(n49) );
  xo2d1_hd U723 ( .A(DP_OP_116J2_127_7148_n3), .B(n1356), .Y(n1113) );
  or2d1_hd U724 ( .A(n773), .B(n786), .Y(n1027) );
  nr2bd1_hd U725 ( .AN(n754), .B(n755), .Y(n1020) );
  or2d1_hd U726 ( .A(n754), .B(n755), .Y(n1001) );
  ad2d1_hd U727 ( .A(n654), .B(n643), .Y(n907) );
  or2d1_hd U728 ( .A(n683), .B(n697), .Y(n945) );
  or2d1_hd U729 ( .A(n828), .B(n827), .Y(n1047) );
  or2d1_hd U730 ( .A(n713), .B(n725), .Y(n976) );
  nid1_hd U731 ( .A(n170), .Y(n1334) );
  ivd1_hd U732 ( .A(n109), .Y(n110) );
  ivd1_hd U733 ( .A(a_m[14]), .Y(n109) );
  ivd1_hd U734 ( .A(a_m[17]), .Y(n91) );
  ivd1_hd U735 ( .A(b_m[10]), .Y(n545) );
  ivd1_hd U736 ( .A(b_m[16]), .Y(n573) );
  ivd1_hd U737 ( .A(b_m[19]), .Y(n587) );
  ivd1_hd U738 ( .A(b_m[15]), .Y(n569) );
  ivd1_hd U739 ( .A(intadd_16_n1), .Y(intadd_0_B_27_) );
  xo2d1_hd U740 ( .A(n610), .B(n1055), .Y(n1060) );
  xo2d1_hd U741 ( .A(n1076), .B(n1075), .Y(n1077) );
  xo2d1_hd U742 ( .A(n85), .B(n879), .Y(n892) );
  xo2d1_hd U743 ( .A(n109), .B(n988), .Y(intadd_16_B_2_) );
  xo2d1_hd U744 ( .A(n463), .B(n958), .Y(intadd_17_B_2_) );
  xo2d1_hd U745 ( .A(n608), .B(n928), .Y(intadd_19_B_2_) );
  xo2d1_hd U746 ( .A(n91), .B(n1013), .Y(intadd_15_B_2_) );
  xo2d1_hd U747 ( .A(a_m[5]), .B(n909), .Y(n912) );
  xo2d1_hd U748 ( .A(n852), .B(n471), .Y(intadd_1_A_21_) );
  xo2d1_hd U749 ( .A(n1042), .B(n116), .Y(n1050) );
  xo2d1_hd U750 ( .A(n995), .B(n124), .Y(n1003) );
  xo2d1_hd U751 ( .A(n937), .B(n607), .Y(n947) );
  xo2d1_hd U752 ( .A(n969), .B(n462), .Y(n978) );
  xo2d1_hd U753 ( .A(n1022), .B(n460), .Y(n1029) );
  xo2d1_hd U754 ( .A(a_m[14]), .B(n977), .Y(intadd_8_B_8_) );
  xo2d1_hd U755 ( .A(n608), .B(n920), .Y(intadd_4_B_16_) );
  xo2d1_hd U756 ( .A(n115), .B(n1028), .Y(intadd_10_B_5_) );
  xo2d1_hd U757 ( .A(n92), .B(n1002), .Y(intadd_11_B_4_) );
  xo2d1_hd U758 ( .A(n86), .B(n866), .Y(intadd_0_A_16_) );
  xo2d1_hd U759 ( .A(n611), .B(n1049), .Y(intadd_14_B_2_) );
  xo2d1_hd U760 ( .A(n114), .B(n1014), .Y(n1030) );
  xo2d1_hd U761 ( .A(n610), .B(n1038), .Y(n1051) );
  xo2d1_hd U762 ( .A(n463), .B(n929), .Y(n949) );
  xo2d1_hd U763 ( .A(n91), .B(n989), .Y(n1005) );
  xo2d1_hd U764 ( .A(n604), .B(n910), .Y(n911) );
  xo2d1_hd U765 ( .A(n126), .B(n959), .Y(n980) );
  xo2d1_hd U766 ( .A(n110), .B(n956), .Y(intadd_8_B_6_) );
  xo2d1_hd U767 ( .A(n612), .B(n1034), .Y(intadd_14_CI) );
  xo2d1_hd U768 ( .A(n116), .B(n1010), .Y(intadd_10_B_3_) );
  xo2d1_hd U769 ( .A(n91), .B(n986), .Y(intadd_9_B_7_) );
  xo2d1_hd U770 ( .A(n609), .B(n877), .Y(n893) );
  xo2d1_hd U771 ( .A(n463), .B(n925), .Y(intadd_5_B_11_) );
  xo2d1_hd U772 ( .A(n608), .B(n867), .Y(intadd_4_A_13_) );
  xo2d1_hd U773 ( .A(n115), .B(n1000), .Y(intadd_15_B_1_) );
  xo2d1_hd U774 ( .A(n125), .B(n944), .Y(intadd_17_B_1_) );
  xo2d1_hd U775 ( .A(n91), .B(n975), .Y(intadd_16_B_1_) );
  xo2d1_hd U776 ( .A(n464), .B(n914), .Y(intadd_19_A_1_) );
  xo2d1_hd U777 ( .A(n621), .B(n1024), .Y(intadd_13_A_1_) );
  xo2d1_hd U778 ( .A(n85), .B(n836), .Y(intadd_2_B_16_) );
  xo2d1_hd U779 ( .A(n459), .B(n965), .Y(intadd_16_CI) );
  xo2d1_hd U780 ( .A(n469), .B(n820), .Y(intadd_2_B_15_) );
  xo2d1_hd U781 ( .A(n124), .B(n933), .Y(intadd_17_CI) );
  fad1_hd U782 ( .A(intadd_2_A_11_), .B(intadd_2_B_11_), .CI(intadd_2_n9), 
        .CO(intadd_2_n8), .S(intadd_1_B_14_) );
  xo2d1_hd U783 ( .A(n463), .B(n903), .Y(intadd_19_CI) );
  xo2d1_hd U784 ( .A(a_m[8]), .B(n853), .Y(intadd_0_A_15_) );
  xo2d1_hd U785 ( .A(n470), .B(n767), .Y(intadd_1_A_15_) );
  xo2d1_hd U786 ( .A(n621), .B(n1018), .Y(intadd_13_CI) );
  xo2d1_hd U787 ( .A(n114), .B(n991), .Y(intadd_15_B_0_) );
  xo2d1_hd U788 ( .A(n604), .B(n837), .Y(intadd_0_A_14_) );
  xo2d1_hd U789 ( .A(n467), .B(n801), .Y(intadd_2_B_14_) );
  xo2d1_hd U790 ( .A(n470), .B(n761), .Y(intadd_1_A_14_) );
  xo2d1_hd U791 ( .A(n611), .B(n1009), .Y(n1015) );
  xo2d1_hd U792 ( .A(a_m[14]), .B(n924), .Y(intadd_7_B_8_) );
  xo2d1_hd U793 ( .A(n91), .B(n955), .Y(intadd_18_B_2_) );
  xo2d1_hd U794 ( .A(n469), .B(n793), .Y(intadd_2_B_13_) );
  xo2d1_hd U795 ( .A(n611), .B(n997), .Y(intadd_10_A_2_) );
  xo2d1_hd U796 ( .A(a_m[17]), .B(n943), .Y(intadd_8_B_5_) );
  xo2d1_hd U797 ( .A(n470), .B(n750), .Y(intadd_1_A_13_) );
  xo2d1_hd U798 ( .A(a_m[8]), .B(n824), .Y(intadd_0_A_13_) );
  xo2d1_hd U799 ( .A(n116), .B(n974), .Y(intadd_9_B_6_) );
  xo2d1_hd U800 ( .A(n109), .B(n915), .Y(intadd_5_A_10_) );
  xo2d1_hd U801 ( .A(n1369), .B(n932), .Y(intadd_17_B_0_) );
  xo2d1_hd U802 ( .A(n126), .B(n895), .Y(intadd_19_A_0_) );
  xo2d1_hd U803 ( .A(n115), .B(n964), .Y(intadd_16_B_0_) );
  xo2d1_hd U804 ( .A(a_m[8]), .B(n804), .Y(intadd_0_A_12_) );
  xo2d1_hd U805 ( .A(n611), .B(n990), .Y(intadd_15_A_0_) );
  xo2d1_hd U806 ( .A(n125), .B(n880), .Y(n905) );
  xo2d1_hd U807 ( .A(n611), .B(n984), .Y(intadd_10_CI) );
  xo2d1_hd U808 ( .A(n470), .B(n736), .Y(intadd_1_B_11_) );
  xo2d1_hd U809 ( .A(n469), .B(n766), .Y(intadd_2_B_11_) );
  xo2d1_hd U810 ( .A(n114), .B(n954), .Y(intadd_9_B_4_) );
  xo2d1_hd U811 ( .A(n92), .B(n923), .Y(intadd_8_B_3_) );
  xo2d1_hd U812 ( .A(a_m[8]), .B(n796), .Y(intadd_0_A_11_) );
  xo2d1_hd U813 ( .A(n473), .B(n731), .Y(intadd_1_B_10_) );
  xo2d1_hd U814 ( .A(a_m[17]), .B(n918), .Y(intadd_7_B_7_) );
  xo2d1_hd U815 ( .A(n116), .B(n942), .Y(intadd_18_B_1_) );
  xo2d1_hd U816 ( .A(n124), .B(n869), .Y(intadd_5_A_7_) );
  xo2d1_hd U817 ( .A(a_m[8]), .B(n782), .Y(intadd_0_A_10_) );
  xo2d1_hd U818 ( .A(n469), .B(n760), .Y(intadd_2_B_10_) );
  xo2d1_hd U819 ( .A(n621), .B(n971), .Y(intadd_11_A_1_) );
  xo2d1_hd U820 ( .A(n621), .B(n963), .Y(intadd_11_CI) );
  xo2d1_hd U821 ( .A(n1380), .B(n819), .Y(intadd_4_B_9_) );
  xo2d1_hd U822 ( .A(n109), .B(n861), .Y(intadd_6_B_9_) );
  xo2d1_hd U823 ( .A(n115), .B(n931), .Y(intadd_18_CI) );
  xo2d1_hd U824 ( .A(n468), .B(n737), .Y(intadd_2_A_9_) );
  xo2d1_hd U825 ( .A(n606), .B(n768), .Y(intadd_0_A_9_) );
  xo2d1_hd U826 ( .A(n473), .B(n720), .Y(intadd_1_B_9_) );
  xo2d1_hd U827 ( .A(n1369), .B(n902), .Y(intadd_5_B_9_) );
  xo2d1_hd U828 ( .A(n1082), .B(n1627), .Y(N475) );
  xo2d1_hd U829 ( .A(n459), .B(n882), .Y(intadd_5_A_8_) );
  xo2d1_hd U830 ( .A(n611), .B(n953), .Y(n960) );
  xo2d1_hd U831 ( .A(n473), .B(n707), .Y(intadd_1_B_8_) );
  xo2d1_hd U832 ( .A(n468), .B(n732), .Y(intadd_2_A_8_) );
  xo2d1_hd U833 ( .A(n605), .B(n762), .Y(intadd_0_A_8_) );
  xo2d1_hd U834 ( .A(n126), .B(n838), .Y(intadd_6_A_8_) );
  xo2d1_hd U835 ( .A(n92), .B(n870), .Y(intadd_7_A_4_) );
  xo2d1_hd U836 ( .A(n473), .B(n703), .Y(intadd_1_B_7_) );
  xo2d1_hd U837 ( .A(n468), .B(n721), .Y(intadd_2_A_7_) );
  xo2d1_hd U838 ( .A(n605), .B(n751), .Y(intadd_0_A_7_) );
  xo2d1_hd U839 ( .A(n125), .B(n825), .Y(intadd_6_A_7_) );
  xo2d1_hd U840 ( .A(n612), .B(n939), .Y(intadd_9_A_3_) );
  xo2d1_hd U841 ( .A(DP_OP_125J2_130_6300_n2), .B(n1081), .Y(n1082) );
  xo2d1_hd U842 ( .A(n605), .B(n738), .Y(intadd_0_A_6_) );
  xo2d1_hd U843 ( .A(n467), .B(n708), .Y(intadd_2_A_6_) );
  xo2d1_hd U844 ( .A(n612), .B(n930), .Y(intadd_18_B_0_) );
  xo2d1_hd U845 ( .A(n473), .B(n693), .Y(intadd_1_B_6_) );
  xo2d1_hd U846 ( .A(n459), .B(n860), .Y(intadd_5_B_6_) );
  xo2d1_hd U847 ( .A(n124), .B(n805), .Y(intadd_6_A_6_) );
  xo2d1_hd U848 ( .A(n468), .B(n704), .Y(intadd_2_A_5_) );
  xo2d1_hd U849 ( .A(n605), .B(n733), .Y(intadd_0_A_5_) );
  xo2d1_hd U850 ( .A(n459), .B(n839), .Y(intadd_5_A_5_) );
  xo2d1_hd U851 ( .A(n109), .B(n797), .Y(intadd_6_A_5_) );
  xo2d1_hd U852 ( .A(n473), .B(n679), .Y(intadd_1_A_5_) );
  xo2d1_hd U853 ( .A(n114), .B(n888), .Y(n897) );
  xo2d1_hd U854 ( .A(n612), .B(n921), .Y(intadd_9_B_1_) );
  xo2d1_hd U855 ( .A(n464), .B(n765), .Y(intadd_4_B_5_) );
  xo2d1_hd U856 ( .A(n605), .B(n730), .Y(intadd_0_B_4_) );
  xo2d1_hd U857 ( .A(n474), .B(n678), .Y(intadd_1_B_4_) );
  xo2d1_hd U858 ( .A(n618), .B(n916), .Y(intadd_12_A_1_) );
  xo2d1_hd U859 ( .A(n461), .B(n826), .Y(intadd_5_A_4_) );
  xo2d1_hd U860 ( .A(n126), .B(n791), .Y(intadd_6_B_4_) );
  xo2d1_hd U861 ( .A(n465), .B(n759), .Y(intadd_4_B_4_) );
  xo2d1_hd U862 ( .A(n618), .B(n900), .Y(intadd_12_CI) );
  xo2d1_hd U863 ( .A(n464), .B(n748), .Y(intadd_4_B_3_) );
  xo2d1_hd U864 ( .A(n474), .B(n670), .Y(intadd_1_B_3_) );
  xo2d1_hd U865 ( .A(n461), .B(n806), .Y(intadd_5_A_3_) );
  xo2d1_hd U866 ( .A(n605), .B(n709), .Y(intadd_0_A_3_) );
  xo2d1_hd U867 ( .A(n464), .B(n735), .Y(intadd_4_B_2_) );
  xo2d1_hd U868 ( .A(n474), .B(n660), .Y(intadd_1_B_2_) );
  xo2d1_hd U869 ( .A(n618), .B(n889), .Y(intadd_8_CI) );
  xo2d1_hd U870 ( .A(n461), .B(n799), .Y(intadd_5_B_2_) );
  xo2d1_hd U871 ( .A(n606), .B(n706), .Y(intadd_0_B_2_) );
  nd2bd1_hd U872 ( .AN(n645), .B(n646), .Y(n656) );
  xo2d1_hd U873 ( .A(n126), .B(n752), .Y(intadd_6_A_1_) );
  xo2d1_hd U874 ( .A(n461), .B(n783), .Y(intadd_5_A_1_) );
  xo2d1_hd U875 ( .A(n467), .B(n671), .Y(intadd_2_A_1_) );
  xo2d1_hd U876 ( .A(n612), .B(n874), .Y(n887) );
  xo2d1_hd U877 ( .A(n474), .B(n658), .Y(intadd_1_B_1_) );
  or2d1_hd U878 ( .A(n677), .B(n676), .Y(n690) );
  xo2d1_hd U879 ( .A(n464), .B(n722), .Y(intadd_4_A_1_) );
  xo2d1_hd U880 ( .A(n126), .B(n741), .Y(intadd_6_B_0_) );
  xo2d1_hd U881 ( .A(n468), .B(n663), .Y(intadd_2_B_0_) );
  xo2d1_hd U882 ( .A(n618), .B(n858), .Y(n871) );
  xo2d1_hd U883 ( .A(n472), .B(n651), .Y(intadd_1_B_0_) );
  scg6d1_hd U884 ( .A(n1340), .B(n1338), .C(n112), .Y(n1362) );
  xo2d1_hd U885 ( .A(n463), .B(n712), .Y(intadd_4_B_0_) );
  xo2d1_hd U886 ( .A(n467), .B(n655), .Y(n657) );
  xo2d1_hd U887 ( .A(n461), .B(n756), .Y(n758) );
  xo2d1_hd U888 ( .A(n613), .B(n831), .Y(n833) );
  nid1_hd U889 ( .A(n1377), .Y(n1402) );
  xo2d1_hd U890 ( .A(n612), .B(n841), .Y(n855) );
  nid1_hd U891 ( .A(n407), .Y(n406) );
  nid1_hd U892 ( .A(n934), .Y(n400) );
  xo2d1_hd U893 ( .A(n604), .B(n941), .Y(intadd_9_B_3_) );
  xo2d1_hd U894 ( .A(n111), .B(n999), .Y(intadd_10_B_2_) );
  xo2d1_hd U895 ( .A(n463), .B(n973), .Y(intadd_11_B_1_) );
  or2d1_hd U896 ( .A(n809), .B(n829), .Y(n1048) );
  or2d1_hd U897 ( .A(n643), .B(n653), .Y(n865) );
  nid1_hd U898 ( .A(n203), .Y(n1364) );
  oa22ad1_hd U899 ( .A(a_m[21]), .B(a_m[22]), .C(a_m[22]), .D(a_m[21]), .Y(
        n829) );
  fad2_hd U900 ( .A(intadd_0_A_26_), .B(intadd_8_n1), .CI(intadd_0_n12), .CO(
        intadd_0_n11), .S(N212) );
  xo2d1_hd U901 ( .A(n1380), .B(n800), .Y(intadd_4_B_8_) );
  xo2d1_hd U902 ( .A(n1380), .B(n792), .Y(intadd_4_B_7_) );
  scg2d1_hd U903 ( .A(b_e[3]), .B(n83), .C(C82_DATA2_3), .D(n82), .Y(n324) );
  scg2d1_hd U904 ( .A(b_e[2]), .B(n84), .C(C82_DATA2_2), .D(n81), .Y(n325) );
  scg2d1_hd U905 ( .A(n82), .B(n1363), .C(b_e[0]), .D(n84), .Y(n327) );
  xo2d1_hd U906 ( .A(n1380), .B(n780), .Y(intadd_4_B_6_) );
  scg2d1_hd U907 ( .A(b_e[5]), .B(n83), .C(C82_DATA2_5), .D(n82), .Y(n322) );
  scg2d1_hd U908 ( .A(b_e[6]), .B(n84), .C(C82_DATA2_6), .D(n81), .Y(n321) );
  scg2d1_hd U909 ( .A(b_e[4]), .B(n84), .C(C82_DATA2_4), .D(n81), .Y(n323) );
  scg2d1_hd U910 ( .A(a_e[5]), .B(n79), .C(C81_DATA2_5), .D(n78), .Y(n313) );
  scg2d1_hd U911 ( .A(a_e[6]), .B(n80), .C(C81_DATA2_6), .D(n77), .Y(n312) );
  scg2d1_hd U912 ( .A(n78), .B(n1348), .C(a_e[0]), .D(n80), .Y(n318) );
  scg2d1_hd U913 ( .A(a_e[2]), .B(n80), .C(C81_DATA2_2), .D(n77), .Y(n316) );
  scg2d1_hd U914 ( .A(a_e[3]), .B(n79), .C(C81_DATA2_3), .D(n78), .Y(n315) );
  scg2d1_hd U915 ( .A(a_e[4]), .B(n80), .C(C81_DATA2_4), .D(n77), .Y(n314) );
  xo2d1_hd U916 ( .A(n1391), .B(n702), .Y(intadd_2_B_4_) );
  xo2d1_hd U917 ( .A(n125), .B(n769), .Y(intadd_6_A_3_) );
  scg9d1_hd U918 ( .A(n83), .B(n1409), .C(n378), .Y(n1411) );
  xo2d1_hd U919 ( .A(n1391), .B(n682), .Y(intadd_2_A_3_) );
  scg9d1_hd U920 ( .A(n641), .B(n640), .C(intadd_1_CI), .Y(N179) );
  xo2d1_hd U921 ( .A(n1391), .B(n681), .Y(intadd_2_B_2_) );
  scg2d1_hd U922 ( .A(n483), .B(a[0]), .C(n123), .D(a_m[0]), .Y(n349) );
  scg9d1_hd U923 ( .A(n79), .B(n1349), .C(n380), .Y(n1351) );
  xo2d1_hd U924 ( .A(n124), .B(n764), .Y(intadd_6_B_2_) );
  nid1_hd U925 ( .A(n198), .Y(n1276) );
  xo2d1_hd U926 ( .A(n606), .B(n694), .Y(intadd_0_A_1_) );
  scg9d1_hd U927 ( .A(n701), .B(n700), .C(n711), .Y(intadd_0_B_1_) );
  scg9d1_hd U928 ( .A(n635), .B(n634), .C(n636), .Y(N178) );
  xo2d1_hd U929 ( .A(n606), .B(n692), .Y(intadd_0_CI) );
  xo2d1_hd U930 ( .A(n116), .B(n798), .Y(n807) );
  scg8d1_hd U931 ( .A(n1369), .B(n746), .C(n745), .D(n744), .Y(n747) );
  scg8d1_hd U932 ( .A(n609), .B(n668), .C(n667), .D(n666), .Y(n669) );
  xo2d1_hd U933 ( .A(n1369), .B(n772), .Y(intadd_5_B_0_) );
  xo2d1_hd U934 ( .A(n110), .B(n734), .Y(n739) );
  xo2d1_hd U935 ( .A(n86), .B(n659), .Y(n661) );
  or2d1_hd U936 ( .A(n1627), .B(n96), .Y(n1302) );
  xo2d1_hd U937 ( .A(n609), .B(n680), .Y(n689) );
  scg6d1_hd U938 ( .A(n1408), .B(n1338), .C(n1377), .Y(n1347) );
  xo2d1_hd U939 ( .A(a_m[17]), .B(n763), .Y(n770) );
  xo2d1_hd U940 ( .A(n110), .B(n727), .Y(n728) );
  scg10d1_hd U941 ( .A(n1175), .B(n1136), .C(z[31]), .D(n454), .Y(n229) );
  xo2d1_hd U942 ( .A(n609), .B(n675), .Y(n677) );
  scg2d1_hd U943 ( .A(n481), .B(b[0]), .C(b_m[0]), .D(n87), .Y(n308) );
  nid1_hd U944 ( .A(n454), .Y(n453) );
  scg2d1_hd U945 ( .A(z_e[1]), .B(n90), .C(n496), .D(DP_OP_125J2_130_6300_n35), 
        .Y(DP_OP_125J2_130_6300_n25) );
  scg2d1_hd U946 ( .A(z_e[2]), .B(n89), .C(n496), .D(DP_OP_125J2_130_6300_n36), 
        .Y(DP_OP_125J2_130_6300_n26) );
  scg2d1_hd U947 ( .A(z_e[3]), .B(n90), .C(n496), .D(DP_OP_125J2_130_6300_n37), 
        .Y(DP_OP_125J2_130_6300_n27) );
  scg2d1_hd U948 ( .A(z_e[4]), .B(n89), .C(n496), .D(DP_OP_125J2_130_6300_n38), 
        .Y(DP_OP_125J2_130_6300_n28) );
  scg2d1_hd U949 ( .A(z_e[5]), .B(n90), .C(n495), .D(DP_OP_125J2_130_6300_n39), 
        .Y(DP_OP_125J2_130_6300_n29) );
  scg2d1_hd U950 ( .A(z_e[6]), .B(n89), .C(n495), .D(DP_OP_125J2_130_6300_n40), 
        .Y(DP_OP_125J2_130_6300_n30) );
  scg2d1_hd U951 ( .A(z_e[7]), .B(n90), .C(n495), .D(DP_OP_125J2_130_6300_n41), 
        .Y(DP_OP_125J2_130_6300_n31) );
  scg2d1_hd U952 ( .A(z_e[8]), .B(n89), .C(n495), .D(DP_OP_125J2_130_6300_n42), 
        .Y(DP_OP_125J2_130_6300_n32) );
  ad2d1_hd U953 ( .A(n101), .B(n614), .Y(n1405) );
  xn2d1_hd U954 ( .A(n638), .B(n513), .Y(n840) );
  scg2d1_hd U955 ( .A(n482), .B(a[29]), .C(n102), .D(a_e[6]), .Y(C1_Z_6) );
  scg2d1_hd U956 ( .A(n483), .B(a[24]), .C(n101), .D(a_e[1]), .Y(C1_Z_1) );
  scg2d1_hd U957 ( .A(n483), .B(a[25]), .C(n101), .D(a_e[2]), .Y(C1_Z_2) );
  scg2d1_hd U958 ( .A(n483), .B(a[26]), .C(n102), .D(a_e[3]), .Y(C1_Z_3) );
  scg2d1_hd U959 ( .A(n483), .B(a[27]), .C(n102), .D(a_e[4]), .Y(C1_Z_4) );
  scg2d1_hd U960 ( .A(n483), .B(a[28]), .C(n101), .D(a_e[5]), .Y(C1_Z_5) );
  or2d1_hd U961 ( .A(n1103), .B(n649), .Y(n810) );
  xn2d1_hd U962 ( .A(n503), .B(n631), .Y(n830) );
  scg2d1_hd U963 ( .A(n482), .B(b[29]), .C(b_e[6]), .D(n106), .Y(n1213) );
  scg2d1_hd U964 ( .A(n482), .B(b[24]), .C(b_e[1]), .D(n103), .Y(n1208) );
  scg2d1_hd U965 ( .A(n482), .B(b[25]), .C(b_e[2]), .D(n103), .Y(n1209) );
  scg2d1_hd U966 ( .A(n482), .B(b[26]), .C(b_e[3]), .D(n106), .Y(n1210) );
  scg2d1_hd U967 ( .A(n482), .B(b[27]), .C(b_e[4]), .D(n103), .Y(n1211) );
  scg2d1_hd U968 ( .A(n481), .B(b[28]), .C(b_e[5]), .D(n103), .Y(n1212) );
  xo2d1_hd U969 ( .A(n460), .B(n1026), .Y(intadd_13_B_1_) );
  scg6d1_hd U970 ( .A(n107), .B(n106), .C(n481), .Y(n1335) );
  nid1_hd U971 ( .A(n993), .Y(n420) );
  ad2d1_hd U972 ( .A(n1115), .B(n1627), .Y(n1123) );
  or2d1_hd U973 ( .A(n673), .B(n674), .Y(n919) );
  or2d1_hd U974 ( .A(n1417), .B(n1183), .Y(n1296) );
  nid1_hd U975 ( .A(n381), .Y(n497) );
  nid1_hd U976 ( .A(n1332), .Y(n484) );
  scg2d1_hd U977 ( .A(n3279), .B(z_m[0]), .C(round_bit), .D(n377), .Y(n1083)
         );
  nid1_hd U978 ( .A(n849), .Y(n384) );
  or2d1_hd U979 ( .A(state[1]), .B(n622), .Y(n381) );
  ad4d1_hd U980 ( .A(n1089), .B(a_e[9]), .C(a_e[0]), .D(a_e[8]), .Y(n1408) );
  ad4d1_hd U981 ( .A(b_e[8]), .B(b_e[9]), .C(n1101), .D(b_e[0]), .Y(n1340) );
  nid1_hd U982 ( .A(n1380), .Y(n466) );
  ivd1_hd U983 ( .A(b_m[0]), .Y(n383) );
  ad2d1_hd U984 ( .A(o_Z_STB), .B(i_Z_ACK), .Y(n177) );
  ivd1_hd U985 ( .A(b_m[1]), .Y(n382) );
  ivd1_hd U986 ( .A(b_m[3]), .Y(n514) );
  ivd1_hd U987 ( .A(b_m[2]), .Y(n509) );
  or4d1_hd U988 ( .A(n14), .B(b_e[6]), .C(b_e[1]), .D(b_e[3]), .Y(n1091) );
  or4d1_hd U989 ( .A(a_e[5]), .B(a_e[4]), .C(a_e[1]), .D(a_e[3]), .Y(n1088) );
  ivd1_hd U990 ( .A(b_m[4]), .Y(n518) );
  or4d1_hd U991 ( .A(product[3]), .B(product[10]), .C(product[11]), .D(
        product[6]), .Y(n1289) );
  ivd1_hd U992 ( .A(z_m[11]), .Y(n16) );
  ivd1_hd U993 ( .A(n16), .Y(n17) );
  ivd1_hd U994 ( .A(z_m[15]), .Y(n18) );
  ivd1_hd U995 ( .A(n18), .Y(n19) );
  ivd1_hd U996 ( .A(z_m[19]), .Y(n20) );
  ivd1_hd U997 ( .A(n20), .Y(n21) );
  ivd1_hd U998 ( .A(z_m[0]), .Y(n22) );
  ivd1_hd U999 ( .A(n22), .Y(n23) );
  ivd1_hd U1000 ( .A(intadd_3_SUM_0_), .Y(n24) );
  ivd1_hd U1001 ( .A(n24), .Y(n25) );
  ivd1_hd U1002 ( .A(intadd_3_SUM_2_), .Y(n26) );
  ivd1_hd U1003 ( .A(n26), .Y(n27) );
  ivd1_hd U1004 ( .A(intadd_3_SUM_1_), .Y(n28) );
  ivd1_hd U1005 ( .A(n28), .Y(n29) );
  ivd1_hd U1006 ( .A(intadd_3_SUM_3_), .Y(n30) );
  ivd1_hd U1007 ( .A(n30), .Y(n31) );
  ivd1_hd U1008 ( .A(intadd_3_SUM_4_), .Y(n32) );
  ivd1_hd U1009 ( .A(n32), .Y(n33) );
  ivd1_hd U1010 ( .A(intadd_3_SUM_6_), .Y(n34) );
  ivd1_hd U1011 ( .A(n34), .Y(n35) );
  ivd1_hd U1012 ( .A(intadd_3_SUM_5_), .Y(n37) );
  ivd1_hd U1013 ( .A(n37), .Y(n38) );
  ivd1_hd U1014 ( .A(intadd_3_SUM_7_), .Y(n39) );
  ivd1_hd U1015 ( .A(n39), .Y(n40) );
  ivd1_hd U1016 ( .A(intadd_3_SUM_8_), .Y(n41) );
  ivd1_hd U1017 ( .A(n41), .Y(n42) );
  ivd1_hd U1018 ( .A(intadd_3_SUM_9_), .Y(n43) );
  ivd1_hd U1019 ( .A(n43), .Y(n44) );
  ivd1_hd U1020 ( .A(intadd_3_SUM_10_), .Y(n45) );
  ivd1_hd U1021 ( .A(n45), .Y(n46) );
  ivd1_hd U1022 ( .A(n47), .Y(n48) );
  ivd1_hd U1023 ( .A(n49), .Y(n50) );
  ivd1_hd U1024 ( .A(n51), .Y(n52) );
  ivd1_hd U1025 ( .A(n53), .Y(n54) );
  ivd1_hd U1026 ( .A(n810), .Y(n67) );
  ivd1_hd U1027 ( .A(n810), .Y(n68) );
  ivd1_hd U1028 ( .A(n840), .Y(n69) );
  ivd1_hd U1029 ( .A(n840), .Y(n70) );
  ivd1_hd U1030 ( .A(n830), .Y(n71) );
  ivd1_hd U1031 ( .A(n830), .Y(n72) );
  ivd1_hd U1032 ( .A(state[1]), .Y(n73) );
  ivd1_hd U1033 ( .A(state[1]), .Y(n74) );
  ivd1_hd U1034 ( .A(n1351), .Y(n77) );
  ivd1_hd U1035 ( .A(n1351), .Y(n78) );
  ivd1_hd U1036 ( .A(n1347), .Y(n79) );
  ivd1_hd U1037 ( .A(n1347), .Y(n80) );
  ivd1_hd U1038 ( .A(n1411), .Y(n81) );
  ivd1_hd U1039 ( .A(n1411), .Y(n82) );
  ivd1_hd U1040 ( .A(n1362), .Y(n83) );
  ivd1_hd U1041 ( .A(n1362), .Y(n84) );
  ivd1_hd U1042 ( .A(n85), .Y(n86) );
  ivd1_hd U1043 ( .A(n1335), .Y(n87) );
  ivd1_hd U1044 ( .A(n1335), .Y(n88) );
  ivd1_hd U1045 ( .A(n1123), .Y(n89) );
  ivd1_hd U1046 ( .A(n1123), .Y(n90) );
  ivd1_hd U1047 ( .A(n1334), .Y(n93) );
  ivd1_hd U1048 ( .A(n1334), .Y(n94) );
  ivd1_hd U1049 ( .A(n1266), .Y(n95) );
  ivd1_hd U1050 ( .A(n1266), .Y(n96) );
  ivd1_hd U1051 ( .A(n1276), .Y(n97) );
  ivd1_hd U1052 ( .A(n1276), .Y(n98) );
  ivd1_hd U1053 ( .A(n1302), .Y(n99) );
  ivd1_hd U1054 ( .A(n1302), .Y(n100) );
  ivd1_hd U1055 ( .A(n1349), .Y(n101) );
  ivd1_hd U1056 ( .A(n1349), .Y(n102) );
  ivd1_hd U1057 ( .A(n1409), .Y(n103) );
  ivd1_hd U1058 ( .A(n1409), .Y(n106) );
  ivd1_hd U1059 ( .A(b_m[23]), .Y(n107) );
  ivd1_hd U1060 ( .A(n107), .Y(n108) );
  ivd1_hd U1061 ( .A(n109), .Y(n111) );
  ivd1_hd U1062 ( .A(n87), .Y(n112) );
  ivd1_hd U1063 ( .A(n88), .Y(n113) );
  ivd1_hd U1064 ( .A(n1364), .Y(n114) );
  ivd1_hd U1065 ( .A(n1364), .Y(n115) );
  ivd1_hd U1066 ( .A(n1364), .Y(n116) );
  ivd1_hd U1067 ( .A(n383), .Y(n117) );
  ivd1_hd U1068 ( .A(n383), .Y(n118) );
  ivd1_hd U1069 ( .A(n383), .Y(n119) );
  ivd1_hd U1070 ( .A(n1402), .Y(n120) );
  ivd1_hd U1071 ( .A(n1402), .Y(n121) );
  ivd1_hd U1072 ( .A(n1402), .Y(n122) );
  ivd1_hd U1073 ( .A(n1402), .Y(n123) );
  ivd1_hd U1074 ( .A(a_m[14]), .Y(n124) );
  ivd1_hd U1075 ( .A(a_m[14]), .Y(n125) );
  ivd1_hd U1076 ( .A(n110), .Y(n126) );
  ivd1_hd U1077 ( .A(n847), .Y(n127) );
  ivd1_hd U1078 ( .A(n847), .Y(n128) );
  ivd1_hd U1079 ( .A(n847), .Y(n129) );
  ivd1_hd U1080 ( .A(n847), .Y(n130) );
  ivd1_hd U1081 ( .A(n927), .Y(n131) );
  ivd1_hd U1082 ( .A(n927), .Y(n132) );
  ivd1_hd U1083 ( .A(n927), .Y(n133) );
  ivd1_hd U1084 ( .A(n927), .Y(n134) );
  ivd1_hd U1085 ( .A(n695), .Y(n135) );
  ivd1_hd U1086 ( .A(n695), .Y(n136) );
  ivd1_hd U1087 ( .A(n695), .Y(n137) );
  ivd1_hd U1088 ( .A(n695), .Y(n139) );
  ivd1_hd U1089 ( .A(n723), .Y(n140) );
  ivd1_hd U1090 ( .A(n723), .Y(n142) );
  ivd1_hd U1091 ( .A(n723), .Y(n143) );
  ivd1_hd U1092 ( .A(n723), .Y(n144) );
  ivd1_hd U1093 ( .A(n1012), .Y(n145) );
  ivd1_hd U1094 ( .A(n1012), .Y(n147) );
  ivd1_hd U1095 ( .A(n1012), .Y(n149) );
  ivd1_hd U1096 ( .A(n1012), .Y(n150) );
  ivd1_hd U1097 ( .A(n784), .Y(n152) );
  ivd1_hd U1098 ( .A(n784), .Y(n153) );
  ivd1_hd U1099 ( .A(n784), .Y(n154) );
  ivd1_hd U1100 ( .A(n784), .Y(n159) );
  ivd1_hd U1101 ( .A(n1405), .Y(n162) );
  ivd1_hd U1102 ( .A(n1405), .Y(n163) );
  ivd1_hd U1103 ( .A(n1405), .Y(n164) );
  ivd1_hd U1104 ( .A(n1405), .Y(n165) );
  ivd1_hd U1105 ( .A(n1048), .Y(n166) );
  ivd1_hd U1106 ( .A(n1048), .Y(n167) );
  ivd1_hd U1107 ( .A(n1048), .Y(n168) );
  ivd1_hd U1108 ( .A(n1048), .Y(n169) );
  ivd1_hd U1109 ( .A(n382), .Y(n170) );
  ivd1_hd U1110 ( .A(n382), .Y(n175) );
  ivd1_hd U1111 ( .A(n382), .Y(n176) );
  ivd1_hd U1112 ( .A(n865), .Y(n178) );
  ivd1_hd U1113 ( .A(n865), .Y(n180) );
  ivd1_hd U1114 ( .A(n865), .Y(n181) );
  ivd1_hd U1115 ( .A(n865), .Y(n182) );
  ivd1_hd U1116 ( .A(n1296), .Y(n183) );
  ivd1_hd U1117 ( .A(n1296), .Y(n184) );
  ivd1_hd U1118 ( .A(n1296), .Y(n185) );
  ivd1_hd U1119 ( .A(n1296), .Y(n186) );
  nid1_hd U1120 ( .A(z_m[7]), .Y(n187) );
  nid1_hd U1121 ( .A(z_m[3]), .Y(n188) );
  ivd1_hd U1122 ( .A(n1226), .Y(n189) );
  ivd1_hd U1123 ( .A(n1199), .Y(n190) );
  nid1_hd U1124 ( .A(n1171), .Y(n191) );
  scg10d1_hd U1125 ( .A(n1139), .B(n1138), .C(n1173), .D(n1143), .Y(n1171) );
  ivd1_hd U1126 ( .A(b_m[0]), .Y(n192) );
  ivd1_hd U1127 ( .A(n117), .Y(n812) );
  ivd1_hd U1128 ( .A(n466), .Y(n193) );
  xo2d1_hd U1129 ( .A(n193), .B(n946), .Y(intadd_7_B_10_) );
  xo2d1_hd U1130 ( .A(n193), .B(n705), .Y(n710) );
  xo2d1_hd U1131 ( .A(a_m[11]), .B(n699), .Y(n700) );
  nid1_hd U1132 ( .A(n99), .Y(n1300) );
  ivd1_hd U1133 ( .A(n1300), .Y(n194) );
  ivd1_hd U1134 ( .A(n1300), .Y(n195) );
  nid1_hd U1135 ( .A(a_m[2]), .Y(n196) );
  nid1_hd U1136 ( .A(a_m[2]), .Y(n197) );
  xo2d1_hd U1137 ( .A(n197), .B(n639), .Y(n640) );
  xo2d1_hd U1138 ( .A(n196), .B(n633), .Y(n634) );
  or2d1_hd U1139 ( .A(n1267), .B(n95), .Y(n1307) );
  ivd1_hd U1140 ( .A(n1307), .Y(n198) );
  ivd1_hd U1141 ( .A(n1307), .Y(n199) );
  nid1_hd U1142 ( .A(b_m[23]), .Y(n1112) );
  ivd1_hd U1143 ( .A(n1112), .Y(n200) );
  ivd1_hd U1144 ( .A(n1112), .Y(n201) );
  ivd1_hd U1145 ( .A(n1112), .Y(n202) );
  nid1_hd U1146 ( .A(a_m[20]), .Y(n204) );
  nid1_hd U1147 ( .A(a_m[20]), .Y(n205) );
  xo2d1_hd U1148 ( .A(n205), .B(n1045), .Y(intadd_14_A_2_) );
  xo2d1_hd U1149 ( .A(n204), .B(n1036), .Y(intadd_13_B_2_) );
  xo2d1_hd U1150 ( .A(a_m[20]), .B(n985), .Y(intadd_11_B_2_) );
  xo2d1_hd U1151 ( .A(n205), .B(n922), .Y(intadd_12_B_2_) );
  xo2d1_hd U1152 ( .A(n204), .B(n917), .Y(intadd_8_B_2_) );
  xo2d1_hd U1153 ( .A(n203), .B(n901), .Y(intadd_7_B_6_) );
  xo2d1_hd U1154 ( .A(n1364), .B(n876), .Y(n883) );
  xo2d1_hd U1155 ( .A(n205), .B(n859), .Y(intadd_7_B_3_) );
  xo2d1_hd U1156 ( .A(n204), .B(n842), .Y(intadd_7_B_2_) );
  xo2d1_hd U1157 ( .A(n203), .B(n834), .Y(intadd_7_B_1_) );
  xo2d1_hd U1158 ( .A(n204), .B(n818), .Y(intadd_7_CI) );
  xo2d1_hd U1159 ( .A(n204), .B(n788), .Y(n789) );
  ivd1_hd U1160 ( .A(n1177), .Y(n206) );
  ivd1_hd U1161 ( .A(n1177), .Y(n207) );
  ivd1_hd U1162 ( .A(n1177), .Y(n208) );
  ivd1_hd U1163 ( .A(n1177), .Y(n209) );
  scg2d1_hd U1164 ( .A(n23), .B(n207), .C(n450), .D(z[0]), .Y(n260) );
  scg2d1_hd U1165 ( .A(z_m[1]), .B(n206), .C(n448), .D(z[1]), .Y(n259) );
  scg2d1_hd U1166 ( .A(z_m[2]), .B(n209), .C(n448), .D(z[2]), .Y(n258) );
  scg2d1_hd U1167 ( .A(n188), .B(n208), .C(n448), .D(z[3]), .Y(n257) );
  scg2d1_hd U1168 ( .A(z_m[4]), .B(n207), .C(n448), .D(z[4]), .Y(n256) );
  scg2d1_hd U1169 ( .A(z_m[5]), .B(n206), .C(n448), .D(z[5]), .Y(n255) );
  scg2d1_hd U1170 ( .A(z_m[6]), .B(n209), .C(n448), .D(z[6]), .Y(n254) );
  scg2d1_hd U1171 ( .A(n187), .B(n208), .C(n449), .D(z[7]), .Y(n253) );
  scg2d1_hd U1172 ( .A(z_m[8]), .B(n207), .C(n449), .D(z[8]), .Y(n252) );
  scg2d1_hd U1173 ( .A(z_m[9]), .B(n206), .C(n449), .D(z[9]), .Y(n251) );
  scg2d1_hd U1174 ( .A(z_m[10]), .B(n209), .C(n449), .D(z[10]), .Y(n250) );
  scg2d1_hd U1175 ( .A(z_m[11]), .B(n208), .C(n449), .D(z[11]), .Y(n249) );
  scg2d1_hd U1176 ( .A(z_m[12]), .B(n207), .C(n449), .D(z[12]), .Y(n248) );
  scg2d1_hd U1177 ( .A(n189), .B(n206), .C(n450), .D(z[13]), .Y(n247) );
  scg2d1_hd U1178 ( .A(z_m[14]), .B(n209), .C(n450), .D(z[14]), .Y(n246) );
  scg2d1_hd U1179 ( .A(z_m[15]), .B(n208), .C(n450), .D(z[15]), .Y(n245) );
  scg2d1_hd U1180 ( .A(z_m[16]), .B(n207), .C(n450), .D(z[16]), .Y(n244) );
  scg2d1_hd U1181 ( .A(n190), .B(n206), .C(n450), .D(z[17]), .Y(n243) );
  scg2d1_hd U1182 ( .A(z_m[18]), .B(n209), .C(n451), .D(z[18]), .Y(n242) );
  scg2d1_hd U1183 ( .A(z_m[19]), .B(n208), .C(n451), .D(z[19]), .Y(n241) );
  scg2d1_hd U1184 ( .A(z_m[20]), .B(n207), .C(n451), .D(z[20]), .Y(n240) );
  scg2d1_hd U1185 ( .A(z_m[21]), .B(n206), .C(n451), .D(z[21]), .Y(n239) );
  or2d1_hd U1186 ( .A(n88), .B(n1409), .Y(n1336) );
  ivd1_hd U1187 ( .A(n1336), .Y(n210) );
  ivd1_hd U1188 ( .A(n1336), .Y(n211) );
  ivd1_hd U1189 ( .A(n1336), .Y(n212) );
  ivd1_hd U1190 ( .A(n1336), .Y(n213) );
  ivd1_hd U1191 ( .A(n630), .Y(n214) );
  ivd1_hd U1192 ( .A(n630), .Y(n215) );
  ivd1_hd U1193 ( .A(n630), .Y(n216) );
  ivd1_hd U1194 ( .A(n630), .Y(n217) );
  or2d1_hd U1195 ( .A(n654), .B(n652), .Y(n864) );
  ivd1_hd U1196 ( .A(n864), .Y(n218) );
  ivd1_hd U1197 ( .A(n864), .Y(n219) );
  ivd1_hd U1198 ( .A(n864), .Y(n220) );
  ivd1_hd U1199 ( .A(n864), .Y(n221) );
  ivd1_hd U1200 ( .A(n919), .Y(n222) );
  ivd1_hd U1201 ( .A(n919), .Y(n223) );
  ivd1_hd U1202 ( .A(n919), .Y(n224) );
  ivd1_hd U1203 ( .A(n919), .Y(n225) );
  ivd1_hd U1204 ( .A(n1001), .Y(n226) );
  ivd1_hd U1205 ( .A(n1001), .Y(n227) );
  ivd1_hd U1206 ( .A(n1001), .Y(n228) );
  ivd1_hd U1207 ( .A(n1001), .Y(n359) );
  ivd1_hd U1208 ( .A(n1047), .Y(n360) );
  ivd1_hd U1209 ( .A(n1047), .Y(n361) );
  ivd1_hd U1210 ( .A(n1047), .Y(n362) );
  ivd1_hd U1211 ( .A(n1047), .Y(n363) );
  ivd1_hd U1212 ( .A(n945), .Y(n364) );
  ivd1_hd U1213 ( .A(n945), .Y(n365) );
  ivd1_hd U1214 ( .A(n945), .Y(n366) );
  ivd1_hd U1215 ( .A(n945), .Y(n367) );
  ivd1_hd U1216 ( .A(n976), .Y(n368) );
  ivd1_hd U1217 ( .A(n976), .Y(n369) );
  ivd1_hd U1218 ( .A(n976), .Y(n370) );
  ivd1_hd U1219 ( .A(n976), .Y(n371) );
  ivd1_hd U1220 ( .A(n1027), .Y(n372) );
  ivd1_hd U1221 ( .A(n1027), .Y(n373) );
  ivd1_hd U1222 ( .A(n1027), .Y(n374) );
  ivd1_hd U1223 ( .A(n1027), .Y(n375) );
  or2d1_hd U1224 ( .A(n73), .B(n622), .Y(n1627) );
  ivd1_hd U1225 ( .A(n1627), .Y(n376) );
  ivd1_hd U1226 ( .A(n1627), .Y(n377) );
  ad2d1_hd U1227 ( .A(n1111), .B(n1116), .Y(n1624) );
  ivd1_hd U1228 ( .A(n1624), .Y(n378) );
  ivd1_hd U1229 ( .A(n1624), .Y(n379) );
  ivd1_hd U1230 ( .A(n1624), .Y(n380) );
  ivd1_hd U1231 ( .A(n378), .Y(n1332) );
  oa211d1_hd U1232 ( .A(n1419), .B(n1418), .C(n1417), .D(n498), .Y(n3276) );
  scg12d1_hd U1233 ( .A(n755), .B(n754), .C(n753), .Y(n1019) );
  ivd1_hd U1234 ( .A(n787), .Y(n773) );
  scg12d1_hd U1235 ( .A(n787), .B(n786), .C(n785), .Y(n1039) );
  scg4d1_hd U1236 ( .A(n592), .B(n360), .C(b_m[19]), .D(n440), .E(n166), .F(
        n588), .G(n447), .H(n62), .Y(n1034) );
  ivd1_hd U1237 ( .A(n1178), .Y(n454) );
  scg12d1_hd U1238 ( .A(n674), .B(n673), .C(n672), .Y(n934) );
  ivd1_hd U1239 ( .A(n1006), .Y(intadd_0_B_28_) );
  scg12d1_hd U1240 ( .A(n726), .B(n725), .C(n724), .Y(n992) );
  ivd1_hd U1241 ( .A(intadd_10_n1), .Y(intadd_0_B_32_) );
  ivd1_hd U1242 ( .A(n617), .Y(n612) );
  ivd1_hd U1243 ( .A(n617), .Y(n611) );
  ivd1_hd U1244 ( .A(n616), .Y(n614) );
  ivd1_hd U1245 ( .A(n809), .Y(n827) );
  ivd1_hd U1246 ( .A(n381), .Y(n489) );
  ivd1_hd U1247 ( .A(n381), .Y(n490) );
  ivd1_hd U1248 ( .A(n454), .Y(n451) );
  ivd1_hd U1249 ( .A(n453), .Y(n450) );
  ivd1_hd U1250 ( .A(n453), .Y(n449) );
  ivd1_hd U1251 ( .A(n453), .Y(n448) );
  ivd1_hd U1252 ( .A(n453), .Y(n452) );
  ivd1_hd U1253 ( .A(n1143), .Y(n1174) );
  ivd1_hd U1254 ( .A(n1292), .Y(n1303) );
  ivd1_hd U1255 ( .A(n105), .Y(n1294) );
  ivd1_hd U1256 ( .A(n1222), .Y(n1267) );
  ivd1_hd U1257 ( .A(n1138), .Y(n1134) );
  scg17d1_hd U1258 ( .A(n1179), .B(n22), .C(net908), .D(n1222), .Y(n1419) );
  ivd1_hd U1259 ( .A(n497), .Y(n495) );
  ivd1_hd U1260 ( .A(n950), .Y(intadd_0_B_22_) );
  ivd1_hd U1261 ( .A(n981), .Y(intadd_0_B_25_) );
  scg12d1_hd U1262 ( .A(n698), .B(n697), .C(n696), .Y(n966) );
  ivd1_hd U1263 ( .A(intadd_16_SUM_2_), .Y(intadd_0_A_26_) );
  ivd1_hd U1264 ( .A(n726), .Y(n713) );
  ivd1_hd U1265 ( .A(intadd_15_SUM_2_), .Y(intadd_0_A_29_) );
  ivd1_hd U1266 ( .A(n1031), .Y(intadd_0_B_31_) );
  ivd1_hd U1267 ( .A(n1043), .Y(intadd_0_A_33_) );
  ivd1_hd U1268 ( .A(n1061), .Y(intadd_0_A_36_) );
  ivd1_hd U1269 ( .A(b_m[22]), .Y(n603) );
  ivd1_hd U1270 ( .A(n617), .Y(n610) );
  ivd1_hd U1271 ( .A(n497), .Y(n494) );
  ivd1_hd U1272 ( .A(n498), .Y(n492) );
  ivd1_hd U1273 ( .A(n498), .Y(n493) );
  ivd1_hd U1274 ( .A(n498), .Y(n491) );
  ivd1_hd U1275 ( .A(n498), .Y(n487) );
  ivd1_hd U1276 ( .A(n498), .Y(n488) );
  ivd1_hd U1277 ( .A(n1165), .Y(n1172) );
  ao21d1_hd U1278 ( .A(n1134), .B(n1122), .C(n1174), .Y(n1178) );
  nr2d1_hd U1279 ( .A(n1628), .B(n1118), .Y(n1114) );
  nr2d1_hd U1280 ( .A(n1122), .B(n1138), .Y(n1338) );
  nd3d1_hd U1281 ( .A(n1139), .B(n1127), .C(n1125), .Y(n1122) );
  ao21d1_hd U1282 ( .A(n377), .B(n1310), .C(n1290), .Y(n1417) );
  nr2d1_hd U1283 ( .A(n1629), .B(n1115), .Y(n1222) );
  ivd1_hd U1284 ( .A(n497), .Y(n496) );
  nr2d1_hd U1285 ( .A(state[3]), .B(n1629), .Y(n1116) );
  ivd1_hd U1286 ( .A(state[0]), .Y(n1629) );
  ivd1_hd U1287 ( .A(n894), .Y(intadd_0_A_18_) );
  ivd1_hd U1288 ( .A(intadd_4_SUM_16_), .Y(intadd_0_B_19_) );
  fad1_hd U1289 ( .A(n913), .B(n912), .CI(n911), .CO(intadd_0_A_19_), .S(
        intadd_0_B_18_) );
  ivd1_hd U1290 ( .A(intadd_17_SUM_2_), .Y(intadd_0_A_23_) );
  ivd1_hd U1291 ( .A(intadd_17_n1), .Y(intadd_0_B_24_) );
  ivd1_hd U1292 ( .A(n698), .Y(n683) );
  ivd1_hd U1293 ( .A(n970), .Y(intadd_0_A_24_) );
  ivd1_hd U1294 ( .A(n196), .Y(n1397) );
  ivd1_hd U1295 ( .A(n996), .Y(intadd_0_A_27_) );
  ivd1_hd U1296 ( .A(a_m[13]), .Y(n1376) );
  ivd1_hd U1297 ( .A(n607), .Y(n606) );
  ivd1_hd U1298 ( .A(n602), .Y(n599) );
  ivd1_hd U1299 ( .A(intadd_10_SUM_5_), .Y(intadd_0_A_31_) );
  ivd1_hd U1300 ( .A(n616), .Y(n613) );
  fad1_hd U1301 ( .A(n1051), .B(intadd_14_SUM_1_), .CI(n1050), .CO(n1052), .S(
        n1043) );
  ivd1_hd U1302 ( .A(a_m[19]), .Y(n1366) );
  ivd1_hd U1303 ( .A(a_m[18]), .Y(n1368) );
  ivd1_hd U1304 ( .A(intadd_14_n1), .Y(intadd_0_B_35_) );
  ivd1_hd U1305 ( .A(n602), .Y(n600) );
  ivd1_hd U1306 ( .A(n596), .Y(n592) );
  ivd1_hd U1307 ( .A(n1058), .Y(intadd_0_A_35_) );
  scg14d1_hd U1308 ( .A(n582), .B(n88), .C(n1315), .Y(n290) );
  scg14d1_hd U1309 ( .A(n535), .B(n87), .C(n1325), .Y(n300) );
  scg14d1_hd U1310 ( .A(n563), .B(n88), .C(n1319), .Y(n294) );
  scg14d1_hd U1311 ( .A(n554), .B(n87), .C(n1321), .Y(n296) );
  scg14d1_hd U1312 ( .A(n521), .B(n88), .C(n1328), .Y(n303) );
  scg14d1_hd U1313 ( .A(n526), .B(n88), .C(n1327), .Y(n302) );
  scg14d1_hd U1314 ( .A(n578), .B(n87), .C(n1316), .Y(n291) );
  scg14d1_hd U1315 ( .A(n588), .B(n87), .C(n1313), .Y(n288) );
  scg17d1_hd U1316 ( .A(z_m[4]), .B(n100), .C(n1265), .D(n1264), .Y(n278) );
  scg17d1_hd U1317 ( .A(z_m[8]), .B(n99), .C(n1247), .D(n1246), .Y(n274) );
  scg17d1_hd U1318 ( .A(z_m[12]), .B(n100), .C(n1230), .D(n1229), .Y(n270) );
  scg17d1_hd U1319 ( .A(z_m[16]), .B(n99), .C(n1203), .D(n1202), .Y(n266) );
  oa21d1_hd U1320 ( .A(z_e[7]), .B(z_e[8]), .C(n1137), .Y(n1173) );
  ivd1_hd U1321 ( .A(z_e[9]), .Y(n1137) );
  scg17d1_hd U1322 ( .A(z_m[20]), .B(n100), .C(n1185), .D(n1184), .Y(n262) );
  ivd1_hd U1323 ( .A(n1121), .Y(n1118) );
  nr2d1_hd U1324 ( .A(state[3]), .B(state[0]), .Y(n1121) );
  ivd1_hd U1325 ( .A(state[2]), .Y(n1628) );
  ivd1_hd U1326 ( .A(z_m[23]), .Y(n1310) );
  scg12d1_hd U1327 ( .A(n1240), .B(z_m[10]), .C(n1243), .Y(n1232) );
  scg12d1_hd U1328 ( .A(n1258), .B(z_m[6]), .C(n1261), .Y(n1249) );
  scg12d1_hd U1329 ( .A(z_m[1]), .B(z_m[2]), .C(n22), .Y(n1269) );
  ivd1_hd U1330 ( .A(z_m[22]), .Y(n1306) );
  nr2d1_hd U1331 ( .A(state[1]), .B(state[2]), .Y(n1111) );
  fad1_hd U1332 ( .A(n893), .B(n892), .CI(intadd_4_SUM_14_), .CO(n894), .S(
        n891) );
  nr2d1_hd U1333 ( .A(n626), .B(n625), .Y(n635) );
  nr2d1_hd U1334 ( .A(n623), .B(n1401), .Y(n850) );
  ivd1_hd U1335 ( .A(a_m[0]), .Y(n1401) );
  ivd1_hd U1336 ( .A(a_m[1]), .Y(n1399) );
  ivd1_hd U1337 ( .A(n607), .Y(n605) );
  ivd1_hd U1338 ( .A(a_m[3]), .Y(n1395) );
  ivd1_hd U1339 ( .A(a_m[4]), .Y(n1393) );
  ivd1_hd U1340 ( .A(a_m[6]), .Y(n1389) );
  ivd1_hd U1341 ( .A(n508), .Y(n505) );
  fad1_hd U1342 ( .A(n980), .B(n979), .CI(n978), .CO(n981), .S(n970) );
  ivd1_hd U1343 ( .A(a_m[10]), .Y(n1382) );
  ivd1_hd U1344 ( .A(a_m[9]), .Y(n1384) );
  ivd1_hd U1345 ( .A(n508), .Y(n504) );
  fad1_hd U1346 ( .A(n1005), .B(n1004), .CI(n1003), .CO(n1006), .S(n996) );
  ivd1_hd U1347 ( .A(a_m[12]), .Y(n1378) );
  ivd1_hd U1348 ( .A(n586), .Y(n583) );
  ivd1_hd U1349 ( .A(a_m[15]), .Y(n1373) );
  ivd1_hd U1350 ( .A(a_m[16]), .Y(n1371) );
  ivd1_hd U1351 ( .A(n540), .Y(n536) );
  ivd1_hd U1352 ( .A(a_m[21]), .Y(n1404) );
  nr2d1_hd U1353 ( .A(state[2]), .B(n74), .Y(n1087) );
  nr2d1_hd U1354 ( .A(n1124), .B(state[0]), .Y(n1120) );
  nr2d1_hd U1355 ( .A(n36), .B(n1183), .Y(n1290) );
  nr2d1_hd U1356 ( .A(n614), .B(n597), .Y(n1073) );
  fad1_hd U1357 ( .A(intadd_1_A_21_), .B(intadd_1_B_21_), .CI(intadd_1_n3), 
        .CO(intadd_1_n2), .S(intadd_1_SUM_21_) );
  fad1_hd U1358 ( .A(intadd_2_A_6_), .B(intadd_2_B_6_), .CI(intadd_2_n14), 
        .CO(intadd_2_n13), .S(intadd_1_A_9_) );
  ivd1_hd U1359 ( .A(n518), .Y(n517) );
  ivd1_hd U1360 ( .A(n530), .Y(n529) );
  ivd1_hd U1361 ( .A(n545), .Y(n544) );
  ivd1_hd U1362 ( .A(n559), .Y(n558) );
  ivd1_hd U1363 ( .A(n568), .Y(n567) );
  nid2_hd U1364 ( .A(n392), .Y(n394) );
  ivd1_hd U1365 ( .A(n597), .Y(n595) );
  ivd1_hd U1366 ( .A(n643), .Y(n652) );
  ivd1_hd U1367 ( .A(n518), .Y(n516) );
  ivd1_hd U1368 ( .A(n530), .Y(n528) );
  ivd1_hd U1369 ( .A(n545), .Y(n543) );
  ivd1_hd U1370 ( .A(n559), .Y(n557) );
  ivd1_hd U1371 ( .A(n568), .Y(n566) );
  ivd1_hd U1372 ( .A(n540), .Y(n537) );
  ivd1_hd U1373 ( .A(n508), .Y(n507) );
  ivd1_hd U1374 ( .A(n550), .Y(n546) );
  ivd1_hd U1375 ( .A(n513), .Y(n512) );
  ivd1_hd U1376 ( .A(n518), .Y(n515) );
  ivd1_hd U1377 ( .A(n513), .Y(n510) );
  ivd1_hd U1378 ( .A(n616), .Y(n615) );
  ivd1_hd U1379 ( .A(n509), .Y(n506) );
  ivd1_hd U1380 ( .A(n513), .Y(n511) );
  ivd1_hd U1381 ( .A(n530), .Y(n527) );
  ivd1_hd U1382 ( .A(n597), .Y(n594) );
  ivd1_hd U1383 ( .A(n545), .Y(n542) );
  ivd1_hd U1384 ( .A(n573), .Y(n571) );
  ivd1_hd U1385 ( .A(n540), .Y(n538) );
  ivd1_hd U1386 ( .A(n540), .Y(n539) );
  ivd1_hd U1387 ( .A(n550), .Y(n547) );
  ivd1_hd U1388 ( .A(n550), .Y(n549) );
  ivd1_hd U1389 ( .A(n573), .Y(n570) );
  ivd1_hd U1390 ( .A(n551), .Y(n548) );
  ivd1_hd U1391 ( .A(n559), .Y(n556) );
  ivd1_hd U1392 ( .A(n586), .Y(n584) );
  ivd1_hd U1393 ( .A(n573), .Y(n572) );
  ivd1_hd U1394 ( .A(n568), .Y(n565) );
  ivd1_hd U1395 ( .A(n597), .Y(n593) );
  ivd1_hd U1396 ( .A(n586), .Y(n585) );
  ivd1_hd U1397 ( .A(n602), .Y(n601) );
  ao22d1_hd U1398 ( .A(n496), .B(DP_OP_125J2_130_6300_n34), .C(z_e[0]), .D(n89), .Y(n3277) );
  ivd1_hd U1399 ( .A(n627), .Y(N176) );
  nr2d1_hd U1400 ( .A(n118), .B(n175), .Y(n1103) );
  nr2d1_hd U1401 ( .A(n812), .B(n93), .Y(n649) );
  oa22d1_hd U1402 ( .A(n472), .B(n1399), .C(a_m[1]), .D(n197), .Y(n623) );
  oa22d1_hd U1403 ( .A(n812), .B(n847), .C(n93), .D(n630), .Y(n624) );
  ao21d1_hd U1404 ( .A(n68), .B(n389), .C(n624), .Y(n629) );
  nr3d1_hd U1405 ( .A(n629), .B(n627), .C(n471), .Y(n628) );
  ao211d1_hd U1406 ( .A(n629), .B(n471), .C(n635), .D(n628), .Y(N177) );
  nr2d1_hd U1407 ( .A(n119), .B(n93), .Y(n631) );
  nr2d1_hd U1408 ( .A(a_m[0]), .B(n632), .Y(n849) );
  scg4d1_hd U1409 ( .A(n505), .B(n214), .C(n175), .D(n127), .E(n850), .F(n72), 
        .G(n385), .H(n119), .Y(n633) );
  oa22d1_hd U1410 ( .A(n1395), .B(n197), .C(n471), .D(a_m[3]), .Y(n643) );
  nr2d1_hd U1411 ( .A(n503), .B(n94), .Y(n637) );
  ao22d1_hd U1412 ( .A(n118), .B(n637), .C(n503), .D(n93), .Y(n638) );
  scg4d1_hd U1413 ( .A(intadd_3_B_0_), .B(n216), .C(n170), .D(n385), .E(n391), 
        .F(n70), .G(n129), .H(n504), .Y(n639) );
  oa22d1_hd U1414 ( .A(n1393), .B(n1395), .C(a_m[3]), .D(a_m[4]), .Y(n653) );
  ao22d1_hd U1415 ( .A(a_m[4]), .B(n86), .C(n469), .D(n1393), .Y(n654) );
  ao22d1_hd U1416 ( .A(n170), .B(n218), .C(n68), .D(n396), .Y(n644) );
  oa21d1_hd U1417 ( .A(n812), .B(n865), .C(n644), .Y(n647) );
  nr2d1_hd U1418 ( .A(n467), .B(n647), .Y(n646) );
  scg17d1_hd U1419 ( .A(n467), .B(n647), .C(n646), .D(n645), .Y(n648) );
  nr2d1_hd U1420 ( .A(n503), .B(n649), .Y(n650) );
  oa22d1_hd U1421 ( .A(n513), .B(n650), .C(n94), .D(n508), .Y(intadd_3_CI) );
  scg4d1_hd U1422 ( .A(n515), .B(n215), .C(n506), .D(n386), .E(n388), .F(n25), 
        .G(intadd_3_B_0_), .H(n128), .Y(n651) );
  ivd1_hd U1423 ( .A(intadd_1_SUM_0_), .Y(N180) );
  scg4d1_hd U1424 ( .A(n505), .B(n219), .C(n176), .D(n180), .E(n395), .F(n117), 
        .G(n71), .H(n396), .Y(n655) );
  scg6d1_hd U1425 ( .A(n657), .B(n656), .C(n662), .Y(intadd_1_A_1_) );
  scg4d1_hd U1426 ( .A(n517), .B(n130), .C(n511), .D(n387), .E(n388), .F(n29), 
        .G(n217), .H(intadd_3_B_2_), .Y(n658) );
  ivd1_hd U1427 ( .A(intadd_1_SUM_1_), .Y(N181) );
  ao22d1_hd U1428 ( .A(a_m[6]), .B(n85), .C(a_m[5]), .D(n1389), .Y(n674) );
  nr2d1_hd U1429 ( .A(n812), .B(n674), .Y(n665) );
  scg4d1_hd U1430 ( .A(intadd_3_B_0_), .B(n220), .C(n1334), .D(n394), .E(n69), 
        .F(n398), .G(n504), .H(n181), .Y(n659) );
  xn3d1_hd U1431 ( .A(n665), .B(n661), .C(n662), .Y(intadd_1_A_2_) );
  scg4d1_hd U1432 ( .A(n517), .B(n384), .C(n522), .D(n127), .E(n523), .F(n214), 
        .G(n389), .H(n27), .Y(n660) );
  ivd1_hd U1433 ( .A(intadd_1_SUM_2_), .Y(N182) );
  oa21d1_hd U1434 ( .A(n665), .B(n662), .C(n661), .Y(intadd_2_A_0_) );
  scg4d1_hd U1435 ( .A(n517), .B(n221), .C(n507), .D(n394), .E(n182), .F(n512), 
        .G(n397), .H(n25), .Y(n663) );
  ivd1_hd U1436 ( .A(a_m[7]), .Y(n1387) );
  oa22d1_hd U1437 ( .A(n1387), .B(a_m[6]), .C(n1389), .D(a_m[7]), .Y(n672) );
  nr2d1_hd U1438 ( .A(a_m[7]), .B(n606), .Y(n1093) );
  ao21d1_hd U1439 ( .A(n604), .B(a_m[7]), .C(n1093), .Y(n673) );
  ao22d1_hd U1440 ( .A(n176), .B(n222), .C(n67), .D(n404), .Y(n664) );
  oa21d1_hd U1441 ( .A(n812), .B(n927), .C(n664), .Y(n668) );
  nr2d1_hd U1442 ( .A(n609), .B(n668), .Y(n666) );
  nr2d1_hd U1443 ( .A(n665), .B(n607), .Y(n667) );
  scg4d1_hd U1444 ( .A(n527), .B(n215), .C(n522), .D(n387), .E(n388), .F(n31), 
        .G(intadd_3_B_3_), .H(n128), .Y(n670) );
  ivd1_hd U1445 ( .A(intadd_1_SUM_3_), .Y(N183) );
  scg4d1_hd U1446 ( .A(n517), .B(n178), .C(n511), .D(n393), .E(n520), .F(n218), 
        .G(n397), .H(n29), .Y(n671) );
  scg4d1_hd U1447 ( .A(n505), .B(n223), .C(n175), .D(n131), .E(n406), .F(n72), 
        .G(n401), .H(n119), .Y(n675) );
  scg14d1_hd U1448 ( .A(n677), .B(n676), .C(n690), .Y(intadd_2_B_1_) );
  scg4d1_hd U1449 ( .A(n529), .B(n129), .C(n524), .D(n387), .E(n388), .F(n33), 
        .G(n216), .H(intadd_3_B_5_), .Y(n678) );
  ivd1_hd U1450 ( .A(intadd_1_SUM_4_), .Y(N184) );
  scg4d1_hd U1451 ( .A(n529), .B(n387), .C(n533), .D(n130), .E(n538), .F(n217), 
        .G(n390), .H(n38), .Y(n679) );
  oa22d1_hd U1452 ( .A(n608), .B(n1384), .C(a_m[9]), .D(n604), .Y(n698) );
  scg4d1_hd U1453 ( .A(n510), .B(n224), .C(n170), .D(n402), .E(n132), .F(
        b_m[2]), .G(n405), .H(n70), .Y(n680) );
  xo3d1_hd U1454 ( .A(n690), .B(n691), .C(n689), .Y(intadd_2_A_2_) );
  scg4d1_hd U1455 ( .A(n516), .B(n394), .C(n519), .D(n180), .E(n525), .F(n219), 
        .G(n397), .H(n27), .Y(n681) );
  ivd1_hd U1456 ( .A(intadd_1_SUM_5_), .Y(N185) );
  scg4d1_hd U1457 ( .A(n529), .B(n220), .C(n522), .D(n393), .E(n181), .F(n526), 
        .G(n397), .H(n31), .Y(n682) );
  oa22d1_hd U1458 ( .A(n462), .B(n1382), .C(a_m[10]), .D(a_m[11]), .Y(n696) );
  nr2d1_hd U1459 ( .A(n698), .B(n696), .Y(n967) );
  oa22d1_hd U1460 ( .A(n1384), .B(n1382), .C(a_m[10]), .D(a_m[9]), .Y(n697) );
  oa22d1_hd U1461 ( .A(n812), .B(n945), .C(n94), .D(n695), .Y(n684) );
  ao21d1_hd U1462 ( .A(n67), .B(n412), .C(n684), .Y(n688) );
  nr2d1_hd U1463 ( .A(n686), .B(n685), .Y(n701) );
  nr3d1_hd U1464 ( .A(n688), .B(n691), .C(n462), .Y(n687) );
  ao211d1_hd U1465 ( .A(n688), .B(n462), .C(n701), .D(n687), .Y(intadd_0_A_0_)
         );
  ao21d1_hd U1466 ( .A(n691), .B(n690), .C(n689), .Y(intadd_0_B_0_) );
  scg4d1_hd U1467 ( .A(n516), .B(n225), .C(n507), .D(n403), .E(n133), .F(n512), 
        .G(n405), .H(n25), .Y(n692) );
  ivd1_hd U1468 ( .A(intadd_0_SUM_0_), .Y(intadd_2_B_3_) );
  scg4d1_hd U1469 ( .A(n537), .B(n127), .C(n542), .D(n214), .E(n849), .F(n535), 
        .G(n390), .H(n35), .Y(n693) );
  ivd1_hd U1470 ( .A(intadd_1_SUM_6_), .Y(N186) );
  scg4d1_hd U1471 ( .A(n516), .B(n134), .C(n512), .D(n403), .E(n521), .F(n222), 
        .G(n405), .H(n29), .Y(n694) );
  scg4d1_hd U1472 ( .A(n506), .B(n135), .C(n176), .D(n365), .E(n411), .F(n117), 
        .G(n71), .H(n412), .Y(n699) );
  ivd1_hd U1473 ( .A(intadd_0_SUM_1_), .Y(intadd_2_A_4_) );
  scg4d1_hd U1474 ( .A(n529), .B(n182), .C(n524), .D(n393), .E(n535), .F(n221), 
        .G(n397), .H(n33), .Y(n702) );
  scg4d1_hd U1475 ( .A(n546), .B(n215), .C(n544), .D(n128), .E(n384), .F(n539), 
        .G(n390), .H(n40), .Y(n703) );
  ivd1_hd U1476 ( .A(intadd_1_SUM_7_), .Y(N187) );
  scg4d1_hd U1477 ( .A(n528), .B(n394), .C(n533), .D(n178), .E(n538), .F(n218), 
        .G(n397), .H(n38), .Y(n704) );
  scg4d1_hd U1478 ( .A(n510), .B(n136), .C(n176), .D(n410), .E(n69), .F(n414), 
        .G(n504), .H(n366), .Y(n705) );
  oa22d1_hd U1479 ( .A(n1378), .B(n462), .C(a_m[11]), .D(a_m[12]), .Y(n726) );
  xo3d1_hd U1480 ( .A(n710), .B(n715), .C(n711), .Y(intadd_0_A_2_) );
  scg4d1_hd U1481 ( .A(n516), .B(n400), .C(n519), .D(n131), .E(n407), .F(n27), 
        .G(n524), .H(n223), .Y(n706) );
  ivd1_hd U1482 ( .A(intadd_0_SUM_2_), .Y(intadd_2_B_5_) );
  scg4d1_hd U1483 ( .A(intadd_3_B_9_), .B(n216), .C(n544), .D(n386), .E(n388), 
        .F(n42), .G(n546), .H(n129), .Y(n707) );
  ivd1_hd U1484 ( .A(intadd_1_SUM_8_), .Y(N188) );
  scg4d1_hd U1485 ( .A(n537), .B(n180), .C(n544), .D(n219), .E(n535), .F(n395), 
        .G(n399), .H(n35), .Y(n708) );
  scg4d1_hd U1486 ( .A(n528), .B(n224), .C(b_m[5]), .D(n403), .E(n132), .F(
        n526), .G(n405), .H(n31), .Y(n709) );
  scg14d1_hd U1487 ( .A(n715), .B(n711), .C(n710), .Y(intadd_4_A_0_) );
  scg4d1_hd U1488 ( .A(n516), .B(n137), .C(n507), .D(n410), .E(n367), .F(n512), 
        .G(n414), .H(intadd_3_SUM_0_), .Y(n712) );
  oa22d1_hd U1489 ( .A(n1376), .B(n124), .C(n111), .D(a_m[13]), .Y(n724) );
  nr2d1_hd U1490 ( .A(n726), .B(n724), .Y(n993) );
  oa22d1_hd U1491 ( .A(n1378), .B(n1376), .C(a_m[13]), .D(a_m[12]), .Y(n725)
         );
  oa22d1_hd U1492 ( .A(n192), .B(n976), .C(n94), .D(n723), .Y(n714) );
  ao21d1_hd U1493 ( .A(n67), .B(n421), .C(n714), .Y(n718) );
  nr2d1_hd U1494 ( .A(n716), .B(n717), .Y(n729) );
  oa211d1_hd U1495 ( .A(n111), .B(n718), .C(n717), .D(n716), .Y(n719) );
  nd2bd1_hd U1496 ( .AN(n729), .B(n719), .Y(intadd_4_CI) );
  ivd1_hd U1497 ( .A(intadd_4_SUM_0_), .Y(intadd_0_B_3_) );
  ivd1_hd U1498 ( .A(intadd_0_SUM_3_), .Y(intadd_2_B_6_) );
  scg4d1_hd U1499 ( .A(n553), .B(n130), .C(n556), .D(n217), .E(n384), .F(n549), 
        .G(n390), .H(n44), .Y(n720) );
  ivd1_hd U1500 ( .A(intadd_1_SUM_9_), .Y(N189) );
  scg4d1_hd U1501 ( .A(n547), .B(n220), .C(n544), .D(n181), .E(n395), .F(n539), 
        .G(n399), .H(n40), .Y(n721) );
  scg4d1_hd U1502 ( .A(n516), .B(n364), .C(n512), .D(n409), .E(n521), .F(n139), 
        .G(n415), .H(intadd_3_SUM_1_), .Y(n722) );
  scg4d1_hd U1503 ( .A(n505), .B(n140), .C(b_m[1]), .D(n369), .E(n419), .F(
        b_m[0]), .G(n71), .H(n421), .Y(n727) );
  oa21d1_hd U1504 ( .A(n729), .B(n728), .C(n740), .Y(intadd_4_B_1_) );
  ivd1_hd U1505 ( .A(intadd_4_SUM_1_), .Y(intadd_0_A_4_) );
  scg4d1_hd U1506 ( .A(n528), .B(n133), .C(n524), .D(n403), .E(n535), .F(n225), 
        .G(n405), .H(n33), .Y(n730) );
  ivd1_hd U1507 ( .A(intadd_0_SUM_4_), .Y(intadd_2_B_7_) );
  scg4d1_hd U1508 ( .A(n554), .B(n387), .C(n558), .D(n127), .E(n561), .F(n214), 
        .G(n390), .H(n46), .Y(n731) );
  ivd1_hd U1509 ( .A(intadd_1_SUM_10_), .Y(N190) );
  scg4d1_hd U1510 ( .A(n554), .B(n221), .C(n543), .D(n393), .E(n182), .F(n549), 
        .G(n907), .H(n42), .Y(n732) );
  scg4d1_hd U1511 ( .A(n528), .B(n403), .C(n533), .D(n134), .E(n407), .F(n38), 
        .G(n536), .H(n222), .Y(n733) );
  ao22d1_hd U1512 ( .A(a_m[15]), .B(n125), .C(n111), .D(n1373), .Y(n755) );
  nr2d1_hd U1513 ( .A(n192), .B(n755), .Y(n743) );
  scg4d1_hd U1514 ( .A(n510), .B(n142), .C(n175), .D(n418), .E(n69), .F(n423), 
        .G(n505), .H(n370), .Y(n734) );
  xo3d1_hd U1515 ( .A(n743), .B(n739), .C(n740), .Y(intadd_4_A_2_) );
  scg4d1_hd U1516 ( .A(n517), .B(n410), .C(n522), .D(n365), .E(n525), .F(n135), 
        .G(n414), .H(intadd_3_SUM_2_), .Y(n735) );
  ivd1_hd U1517 ( .A(intadd_4_SUM_2_), .Y(intadd_0_B_5_) );
  ivd1_hd U1518 ( .A(intadd_0_SUM_5_), .Y(intadd_2_B_8_) );
  scg4d1_hd U1519 ( .A(n565), .B(n215), .C(n558), .D(n386), .E(n391), .F(n50), 
        .G(intadd_3_B_11_), .H(n128), .Y(n736) );
  ivd1_hd U1520 ( .A(intadd_1_SUM_11_), .Y(N191) );
  scg4d1_hd U1521 ( .A(n554), .B(n178), .C(n558), .D(n218), .E(n547), .F(n395), 
        .G(n907), .H(n44), .Y(n737) );
  scg4d1_hd U1522 ( .A(n537), .B(n131), .C(n543), .D(n223), .E(n534), .F(n400), 
        .G(n935), .H(n35), .Y(n738) );
  scg16d1_hd U1523 ( .A(n740), .B(n743), .C(n739), .Y(intadd_6_A_0_) );
  scg4d1_hd U1524 ( .A(n517), .B(n143), .C(n507), .D(n418), .E(n371), .F(
        b_m[3]), .G(n422), .H(n25), .Y(n741) );
  oa22d1_hd U1525 ( .A(n1371), .B(a_m[15]), .C(n1373), .D(a_m[16]), .Y(n753)
         );
  ao22d1_hd U1526 ( .A(a_m[17]), .B(a_m[16]), .C(n1371), .D(n460), .Y(n754) );
  ao22d1_hd U1527 ( .A(b_m[1]), .B(n226), .C(n68), .D(n429), .Y(n742) );
  oa21d1_hd U1528 ( .A(n192), .B(n1012), .C(n742), .Y(n746) );
  nr2d1_hd U1529 ( .A(n1369), .B(n746), .Y(n744) );
  nr2d1_hd U1530 ( .A(n743), .B(n461), .Y(n745) );
  scg4d1_hd U1531 ( .A(n528), .B(n136), .C(b_m[5]), .D(n409), .E(n366), .F(
        n526), .G(n414), .H(intadd_3_SUM_3_), .Y(n748) );
  ivd1_hd U1532 ( .A(intadd_4_SUM_3_), .Y(intadd_0_B_6_) );
  ivd1_hd U1533 ( .A(intadd_0_SUM_6_), .Y(intadd_2_B_9_) );
  scg4d1_hd U1534 ( .A(n567), .B(n129), .C(b_m[14]), .D(n386), .E(n391), .F(
        n48), .G(n216), .H(intadd_3_B_13_), .Y(n749) );
  ivd1_hd U1535 ( .A(intadd_1_SUM_12_), .Y(N192) );
  scg4d1_hd U1536 ( .A(n567), .B(n387), .C(intadd_3_B_13_), .D(n130), .E(n576), 
        .F(n217), .G(n390), .H(n52), .Y(n750) );
  scg4d1_hd U1537 ( .A(n546), .B(n224), .C(n543), .D(n132), .E(n405), .F(n40), 
        .G(n401), .H(n536), .Y(n751) );
  scg4d1_hd U1538 ( .A(b_m[4]), .B(n368), .C(n511), .D(n417), .E(n521), .F(
        n144), .G(n422), .H(n29), .Y(n752) );
  scg4d1_hd U1539 ( .A(n506), .B(n227), .C(n176), .D(n145), .E(n427), .F(n118), 
        .G(n72), .H(n429), .Y(n756) );
  nr2d1_hd U1540 ( .A(n758), .B(n757), .Y(n771) );
  scg6d1_hd U1541 ( .A(n758), .B(n757), .C(n771), .Y(intadd_6_B_1_) );
  scg4d1_hd U1542 ( .A(n528), .B(n367), .C(n523), .D(n409), .E(n535), .F(n137), 
        .G(n967), .H(intadd_3_SUM_4_), .Y(n759) );
  ivd1_hd U1543 ( .A(intadd_4_SUM_4_), .Y(intadd_0_B_7_) );
  ivd1_hd U1544 ( .A(intadd_0_SUM_7_), .Y(intadd_2_A_10_) );
  scg4d1_hd U1545 ( .A(n554), .B(n394), .C(n558), .D(n180), .E(n562), .F(n219), 
        .G(n907), .H(n46), .Y(n760) );
  ivd1_hd U1546 ( .A(intadd_1_SUM_13_), .Y(N193) );
  scg4d1_hd U1547 ( .A(intadd_3_B_15_), .B(n214), .C(n571), .D(n386), .E(n391), 
        .F(n54), .G(n574), .H(n127), .Y(n761) );
  scg4d1_hd U1548 ( .A(n554), .B(n225), .C(n543), .D(n402), .E(n133), .F(n549), 
        .G(n935), .H(n42), .Y(n762) );
  scg4d1_hd U1549 ( .A(n510), .B(n228), .C(n170), .D(n426), .E(n70), .F(n431), 
        .G(n505), .H(n147), .Y(n763) );
  oa22d1_hd U1550 ( .A(n460), .B(n1368), .C(a_m[18]), .D(n92), .Y(n787) );
  xo3d1_hd U1551 ( .A(n771), .B(n770), .C(n775), .Y(intadd_6_A_2_) );
  scg4d1_hd U1552 ( .A(b_m[4]), .B(n418), .C(b_m[5]), .D(n369), .E(n525), .F(
        n140), .G(n422), .H(n27), .Y(n764) );
  scg4d1_hd U1553 ( .A(n529), .B(n410), .C(n533), .D(n364), .E(n538), .F(n139), 
        .G(n967), .H(intadd_3_SUM_5_), .Y(n765) );
  ivd1_hd U1554 ( .A(intadd_4_SUM_5_), .Y(intadd_0_B_8_) );
  ivd1_hd U1555 ( .A(intadd_0_SUM_8_), .Y(intadd_2_A_11_) );
  scg4d1_hd U1556 ( .A(n567), .B(n220), .C(n557), .D(n393), .E(n181), .F(n563), 
        .G(n398), .H(n50), .Y(n766) );
  ivd1_hd U1557 ( .A(intadd_1_SUM_14_), .Y(N194) );
  scg4d1_hd U1558 ( .A(n581), .B(n128), .C(n575), .D(n386), .E(n391), .F(n56), 
        .G(n215), .H(intadd_3_B_16_), .Y(n767) );
  scg4d1_hd U1559 ( .A(n553), .B(n134), .C(n557), .D(n222), .E(n547), .F(n934), 
        .G(n935), .H(n44), .Y(n768) );
  scg4d1_hd U1560 ( .A(n529), .B(n142), .C(b_m[5]), .D(n417), .E(n370), .F(
        n525), .G(n422), .H(n31), .Y(n769) );
  scg16d1_hd U1561 ( .A(n775), .B(n771), .C(n770), .Y(intadd_5_A_0_) );
  scg4d1_hd U1562 ( .A(b_m[4]), .B(n359), .C(n507), .D(n426), .E(n149), .F(
        b_m[3]), .G(n430), .H(intadd_3_SUM_0_), .Y(n772) );
  oa22d1_hd U1563 ( .A(n114), .B(n1366), .C(a_m[19]), .D(n204), .Y(n785) );
  nr2d1_hd U1564 ( .A(n787), .B(n785), .Y(n1040) );
  oa22d1_hd U1565 ( .A(n1368), .B(n1366), .C(a_m[19]), .D(a_m[18]), .Y(n786)
         );
  oa22d1_hd U1566 ( .A(n192), .B(n1027), .C(n93), .D(n784), .Y(n774) );
  ao21d1_hd U1567 ( .A(n67), .B(n436), .C(n774), .Y(n778) );
  nr2d1_hd U1568 ( .A(n776), .B(n777), .Y(n790) );
  oa211d1_hd U1569 ( .A(n205), .B(n778), .C(n777), .D(n776), .Y(n779) );
  nd2bd1_hd U1570 ( .AN(n790), .B(n779), .Y(intadd_5_CI) );
  scg4d1_hd U1571 ( .A(n537), .B(n365), .C(n543), .D(n135), .E(n534), .F(n411), 
        .G(n415), .H(intadd_3_SUM_6_), .Y(n780) );
  ivd1_hd U1572 ( .A(intadd_4_SUM_6_), .Y(intadd_0_B_9_) );
  ivd1_hd U1573 ( .A(intadd_0_SUM_9_), .Y(intadd_2_A_12_) );
  scg4d1_hd U1574 ( .A(n567), .B(n182), .C(b_m[14]), .D(n392), .E(n572), .F(
        n221), .G(n398), .H(n48), .Y(n781) );
  ivd1_hd U1575 ( .A(intadd_1_SUM_15_), .Y(N195) );
  scg4d1_hd U1576 ( .A(n553), .B(n403), .C(n557), .D(n131), .E(n407), .F(n46), 
        .G(b_m[14]), .H(n223), .Y(n782) );
  scg4d1_hd U1577 ( .A(n515), .B(n150), .C(n511), .D(n425), .E(n521), .F(n226), 
        .G(n430), .H(intadd_3_SUM_1_), .Y(n783) );
  scg4d1_hd U1578 ( .A(n506), .B(n152), .C(n175), .D(n373), .E(n435), .F(
        b_m[0]), .G(n71), .H(n436), .Y(n788) );
  oa21d1_hd U1579 ( .A(n790), .B(n789), .C(n808), .Y(intadd_5_B_1_) );
  scg4d1_hd U1580 ( .A(b_m[7]), .B(n371), .C(n524), .D(n417), .E(n534), .F(
        n143), .G(n422), .H(n33), .Y(n791) );
  scg4d1_hd U1581 ( .A(n546), .B(n136), .C(n543), .D(n366), .E(n411), .F(n539), 
        .G(n415), .H(intadd_3_SUM_7_), .Y(n792) );
  ivd1_hd U1582 ( .A(intadd_4_SUM_7_), .Y(intadd_0_B_10_) );
  ivd1_hd U1583 ( .A(intadd_0_SUM_10_), .Y(intadd_2_A_13_) );
  scg4d1_hd U1584 ( .A(n566), .B(n394), .C(n571), .D(n178), .E(n577), .F(n218), 
        .G(n398), .H(n52), .Y(n793) );
  scg4d1_hd U1585 ( .A(n582), .B(n849), .C(intadd_3_B_16_), .D(n129), .E(n589), 
        .F(n216), .G(n389), .H(n64), .Y(n794) );
  ivd1_hd U1586 ( .A(intadd_1_SUM_16_), .Y(N196) );
  scg4d1_hd U1587 ( .A(n592), .B(n217), .C(n584), .D(n385), .E(n850), .F(n62), 
        .G(n588), .H(n130), .Y(n795) );
  scg4d1_hd U1588 ( .A(n566), .B(n224), .C(n557), .D(n402), .E(n132), .F(n563), 
        .G(n935), .H(n50), .Y(n796) );
  scg4d1_hd U1589 ( .A(b_m[7]), .B(n418), .C(n532), .D(n368), .E(n537), .F(
        n144), .G(n422), .H(n38), .Y(n797) );
  oa22d1_hd U1590 ( .A(n115), .B(a_m[21]), .C(n1404), .D(n205), .Y(n809) );
  scg4d1_hd U1591 ( .A(n510), .B(n153), .C(n176), .D(n434), .E(n69), .F(n437), 
        .G(n504), .H(n374), .Y(n798) );
  xo3d1_hd U1592 ( .A(n813), .B(n807), .C(n808), .Y(intadd_5_A_2_) );
  scg4d1_hd U1593 ( .A(n515), .B(n426), .C(n519), .D(n145), .E(n525), .F(n227), 
        .G(n430), .H(intadd_3_SUM_2_), .Y(n799) );
  scg4d1_hd U1594 ( .A(n553), .B(n137), .C(n544), .D(n409), .E(n367), .F(n548), 
        .G(n967), .H(intadd_3_SUM_8_), .Y(n800) );
  ivd1_hd U1595 ( .A(intadd_4_SUM_8_), .Y(intadd_0_B_11_) );
  ivd1_hd U1596 ( .A(intadd_0_SUM_11_), .Y(intadd_2_A_14_) );
  scg4d1_hd U1597 ( .A(n582), .B(n219), .C(n571), .D(n392), .E(n180), .F(n578), 
        .G(n398), .H(n54), .Y(n801) );
  ivd1_hd U1598 ( .A(intadd_1_SUM_17_), .Y(N197) );
  oa22d1_hd U1599 ( .A(n596), .B(n603), .C(n598), .D(intadd_3_A_17_), .Y(n802)
         );
  ivd1_hd U1600 ( .A(n802), .Y(n1066) );
  scg4d1_hd U1601 ( .A(n595), .B(n127), .C(n589), .D(n385), .E(n850), .F(n65), 
        .G(n214), .H(n599), .Y(n803) );
  scg4d1_hd U1602 ( .A(n566), .B(n133), .C(b_m[14]), .D(n402), .E(n572), .F(
        n225), .G(n406), .H(n48), .Y(n804) );
  scg4d1_hd U1603 ( .A(n537), .B(n369), .C(n544), .D(n140), .E(n534), .F(n419), 
        .G(n420), .H(n35), .Y(n805) );
  scg4d1_hd U1604 ( .A(b_m[7]), .B(n228), .C(n520), .D(n425), .E(n147), .F(
        n525), .G(n430), .H(intadd_3_SUM_3_), .Y(n806) );
  ao21d1_hd U1605 ( .A(n813), .B(n808), .C(n807), .Y(intadd_7_A_0_) );
  nr2d1_hd U1606 ( .A(n619), .B(a_m[22]), .Y(n1094) );
  ao21d1_hd U1607 ( .A(a_m[22]), .B(n616), .C(n1094), .Y(n828) );
  ao22d1_hd U1608 ( .A(b_m[1]), .B(n360), .C(n68), .D(n444), .Y(n811) );
  oa21d1_hd U1609 ( .A(n192), .B(n1048), .C(n811), .Y(n816) );
  nr2d1_hd U1610 ( .A(n615), .B(n816), .Y(n814) );
  nr2bd1_hd U1611 ( .AN(n813), .B(n610), .Y(n815) );
  ao211d1_hd U1612 ( .A(n610), .B(n816), .C(n815), .D(n814), .Y(n817) );
  nr2bd1_hd U1613 ( .AN(n832), .B(n817), .Y(intadd_7_B_0_) );
  scg4d1_hd U1614 ( .A(n515), .B(n154), .C(n507), .D(n434), .E(n375), .F(
        b_m[3]), .G(n437), .H(n25), .Y(n818) );
  ivd1_hd U1615 ( .A(intadd_7_SUM_0_), .Y(intadd_5_B_3_) );
  scg4d1_hd U1616 ( .A(n553), .B(n364), .C(n557), .D(n139), .E(n548), .F(n411), 
        .G(n967), .H(intadd_3_SUM_9_), .Y(n819) );
  ivd1_hd U1617 ( .A(intadd_4_SUM_9_), .Y(intadd_0_B_12_) );
  ivd1_hd U1618 ( .A(intadd_0_SUM_12_), .Y(intadd_2_A_15_) );
  scg4d1_hd U1619 ( .A(n582), .B(n181), .C(n575), .D(n393), .E(n585), .F(n220), 
        .G(n907), .H(n56), .Y(n820) );
  ivd1_hd U1620 ( .A(intadd_1_SUM_18_), .Y(N198) );
  scg4d1_hd U1621 ( .A(n595), .B(n849), .C(n600), .D(n128), .E(b_m[23]), .F(
        n215), .G(n389), .H(n60), .Y(n823) );
  scg4d1_hd U1622 ( .A(n566), .B(n400), .C(n570), .D(n134), .E(n407), .F(n52), 
        .G(n575), .H(n222), .Y(n824) );
  scg4d1_hd U1623 ( .A(n546), .B(n142), .C(b_m[10]), .D(n370), .E(n419), .F(
        b_m[9]), .G(n420), .H(n40), .Y(n825) );
  scg4d1_hd U1624 ( .A(n527), .B(n149), .C(b_m[6]), .D(n425), .E(n534), .F(
        n359), .G(n430), .H(intadd_3_SUM_4_), .Y(n826) );
  scg4d1_hd U1625 ( .A(n506), .B(n361), .C(n170), .D(n167), .E(n443), .F(n118), 
        .G(n72), .H(n444), .Y(n831) );
  nr2d1_hd U1626 ( .A(n833), .B(n832), .Y(n854) );
  ao21d1_hd U1627 ( .A(n833), .B(n832), .C(n854), .Y(intadd_7_A_1_) );
  scg4d1_hd U1628 ( .A(b_m[4]), .B(n372), .C(n511), .D(n433), .E(n521), .F(
        n159), .G(n438), .H(n29), .Y(n834) );
  ivd1_hd U1629 ( .A(intadd_7_SUM_1_), .Y(intadd_5_B_4_) );
  scg4d1_hd U1630 ( .A(n553), .B(n410), .C(n557), .D(n365), .E(n562), .F(n135), 
        .G(n414), .H(intadd_3_SUM_10_), .Y(n835) );
  ivd1_hd U1631 ( .A(intadd_4_SUM_10_), .Y(intadd_0_B_13_) );
  ivd1_hd U1632 ( .A(intadd_0_SUM_13_), .Y(intadd_2_A_16_) );
  scg4d1_hd U1633 ( .A(n582), .B(n395), .C(n584), .D(n182), .E(n590), .F(n221), 
        .G(n398), .H(n64), .Y(n836) );
  ivd1_hd U1634 ( .A(intadd_1_SUM_19_), .Y(N199) );
  scg4d1_hd U1635 ( .A(n582), .B(n223), .C(n570), .D(n402), .E(n131), .F(n578), 
        .G(n404), .H(n54), .Y(n837) );
  scg4d1_hd U1636 ( .A(b_m[12]), .B(n143), .C(b_m[10]), .D(n417), .E(n371), 
        .F(n548), .G(n993), .H(n42), .Y(n838) );
  scg4d1_hd U1637 ( .A(n527), .B(n426), .C(n533), .D(n150), .E(n538), .F(n226), 
        .G(n430), .H(intadd_3_SUM_5_), .Y(n839) );
  scg4d1_hd U1638 ( .A(n510), .B(n362), .C(n175), .D(n442), .E(n70), .F(n446), 
        .G(n504), .H(n168), .Y(n841) );
  xo3d1_hd U1639 ( .A(n855), .B(n854), .C(n856), .Y(intadd_7_A_2_) );
  scg4d1_hd U1640 ( .A(n515), .B(n434), .C(n520), .D(n373), .E(n523), .F(n152), 
        .G(n437), .H(n27), .Y(n842) );
  ivd1_hd U1641 ( .A(intadd_7_SUM_2_), .Y(intadd_5_B_5_) );
  scg4d1_hd U1642 ( .A(n566), .B(n136), .C(n558), .D(n409), .E(n366), .F(n563), 
        .G(n413), .H(intadd_3_SUM_11_), .Y(n843) );
  ivd1_hd U1643 ( .A(intadd_4_SUM_11_), .Y(intadd_0_B_14_) );
  ivd1_hd U1644 ( .A(intadd_0_SUM_14_), .Y(intadd_2_A_17_) );
  scg4d1_hd U1645 ( .A(n595), .B(n218), .C(n584), .D(n392), .E(n178), .F(n590), 
        .G(n399), .H(n62), .Y(n844) );
  ao22d1_hd U1646 ( .A(n601), .B(n385), .C(n389), .D(n57), .Y(n846) );
  oa21d1_hd U1647 ( .A(n201), .B(n847), .C(n846), .Y(n848) );
  ivd1_hd U1648 ( .A(intadd_1_SUM_20_), .Y(N200) );
  ao21d1_hd U1649 ( .A(n76), .B(n389), .C(n385), .Y(n851) );
  nr2d1_hd U1650 ( .A(n202), .B(n851), .Y(n852) );
  scg4d1_hd U1651 ( .A(n581), .B(n133), .C(n575), .D(n402), .E(n585), .F(n225), 
        .G(n406), .H(n56), .Y(n853) );
  ivd1_hd U1652 ( .A(n854), .Y(n857) );
  ao21d1_hd U1653 ( .A(n857), .B(n856), .C(n855), .Y(n873) );
  nr2d1_hd U1654 ( .A(n614), .B(n94), .Y(n872) );
  scg4d1_hd U1655 ( .A(n515), .B(n360), .C(n506), .D(n442), .E(n166), .F(n512), 
        .G(n445), .H(intadd_3_SUM_0_), .Y(n858) );
  scg4d1_hd U1656 ( .A(n527), .B(n153), .C(n520), .D(n433), .E(n375), .F(n526), 
        .G(n437), .H(n31), .Y(n859) );
  ivd1_hd U1657 ( .A(intadd_7_SUM_3_), .Y(intadd_5_A_6_) );
  scg4d1_hd U1658 ( .A(n536), .B(n147), .C(b_m[10]), .D(n228), .E(b_m[8]), .F(
        n427), .G(n428), .H(intadd_3_SUM_6_), .Y(n860) );
  scg4d1_hd U1659 ( .A(b_m[12]), .B(n368), .C(n558), .D(n144), .E(n547), .F(
        n419), .G(n993), .H(n44), .Y(n861) );
  scg4d1_hd U1660 ( .A(n566), .B(n367), .C(n561), .D(n966), .E(n571), .F(n137), 
        .G(n413), .H(intadd_3_SUM_12_), .Y(n862) );
  ivd1_hd U1661 ( .A(intadd_4_SUM_12_), .Y(intadd_0_B_15_) );
  ivd1_hd U1662 ( .A(intadd_0_SUM_15_), .Y(intadd_2_A_18_) );
  scg4d1_hd U1663 ( .A(n595), .B(n180), .C(n588), .D(n906), .E(n601), .F(n219), 
        .G(n396), .H(n66), .Y(n863) );
  ivd1_hd U1664 ( .A(intadd_1_SUM_21_), .Y(N201) );
  scg4d1_hd U1665 ( .A(n595), .B(n395), .C(n599), .D(n181), .E(n108), .F(n220), 
        .G(n396), .H(n60), .Y(n866) );
  scg4d1_hd U1666 ( .A(n581), .B(n934), .C(n583), .D(n132), .E(n406), .F(
        intadd_3_SUM_16_), .G(intadd_3_B_17_), .H(n224), .Y(n867) );
  scg4d1_hd U1667 ( .A(n567), .B(n410), .C(n570), .D(n364), .E(n577), .F(n139), 
        .G(n413), .H(intadd_3_SUM_13_), .Y(n868) );
  scg4d1_hd U1668 ( .A(b_m[12]), .B(n418), .C(b_m[13]), .D(n369), .E(n562), 
        .F(n140), .G(n993), .H(n46), .Y(n869) );
  scg4d1_hd U1669 ( .A(n546), .B(n227), .C(n542), .D(n145), .E(n427), .F(n539), 
        .G(n428), .H(intadd_3_SUM_7_), .Y(n870) );
  fad1_hd U1670 ( .A(n873), .B(n872), .CI(n871), .CO(n885), .S(intadd_7_A_3_)
         );
  scg4d1_hd U1671 ( .A(intadd_3_B_1_), .B(n169), .C(n511), .D(n441), .E(n520), 
        .F(n363), .G(n445), .H(intadd_3_SUM_1_), .Y(n874) );
  ivd1_hd U1672 ( .A(n875), .Y(n884) );
  scg4d1_hd U1673 ( .A(b_m[7]), .B(n374), .C(b_m[6]), .D(n433), .E(n532), .F(
        n154), .G(n1040), .H(n33), .Y(n876) );
  ivd1_hd U1674 ( .A(intadd_7_SUM_4_), .Y(intadd_5_B_7_) );
  ivd1_hd U1675 ( .A(intadd_4_SUM_13_), .Y(intadd_0_B_16_) );
  ivd1_hd U1676 ( .A(intadd_0_SUM_16_), .Y(intadd_1_B_22_) );
  ivd1_hd U1677 ( .A(intadd_1_SUM_22_), .Y(N202) );
  scg4d1_hd U1678 ( .A(n595), .B(n222), .C(n583), .D(n401), .E(n134), .F(
        b_m[20]), .G(n404), .H(n62), .Y(n877) );
  ao22d1_hd U1679 ( .A(b_m[22]), .B(n906), .C(n396), .D(n58), .Y(n878) );
  oa21d1_hd U1680 ( .A(n202), .B(n865), .C(n878), .Y(n879) );
  scg4d1_hd U1681 ( .A(n567), .B(n142), .C(b_m[13]), .D(n417), .E(n370), .F(
        n562), .G(n423), .H(n50), .Y(n880) );
  scg4d1_hd U1682 ( .A(n581), .B(n135), .C(n570), .D(n408), .E(n365), .F(n578), 
        .G(n413), .H(intadd_3_SUM_14_), .Y(n881) );
  scg4d1_hd U1683 ( .A(b_m[12]), .B(n359), .C(n542), .D(n425), .E(n149), .F(
        n549), .G(n428), .H(intadd_3_SUM_8_), .Y(n882) );
  fad1_hd U1684 ( .A(n885), .B(n884), .CI(n883), .CO(intadd_7_A_5_), .S(
        intadd_7_B_4_) );
  fad1_hd U1685 ( .A(n471), .B(n887), .CI(n886), .CO(n898), .S(n875) );
  scg4d1_hd U1686 ( .A(n527), .B(n434), .C(n532), .D(n372), .E(n538), .F(n159), 
        .G(n1040), .H(n38), .Y(n888) );
  nr2d1_hd U1687 ( .A(n613), .B(n514), .Y(intadd_8_B_0_) );
  scg4d1_hd U1688 ( .A(intadd_3_B_1_), .B(n442), .C(n520), .D(n167), .E(b_m[6]), .F(n361), .G(n445), .H(intadd_3_SUM_2_), .Y(n889) );
  ivd1_hd U1689 ( .A(intadd_8_SUM_0_), .Y(n896) );
  ivd1_hd U1690 ( .A(n890), .Y(intadd_7_B_5_) );
  ivd1_hd U1691 ( .A(intadd_7_SUM_5_), .Y(intadd_5_B_8_) );
  ivd1_hd U1692 ( .A(n891), .Y(intadd_0_B_17_) );
  scg4d1_hd U1693 ( .A(b_m[15]), .B(n371), .C(n564), .D(n992), .E(n571), .F(
        n143), .G(n423), .H(n48), .Y(n895) );
  fad1_hd U1694 ( .A(n898), .B(n897), .CI(n896), .CO(n899), .S(n890) );
  ivd1_hd U1695 ( .A(n899), .Y(intadd_8_A_1_) );
  nr2d1_hd U1696 ( .A(n613), .B(n518), .Y(intadd_12_B_0_) );
  scg4d1_hd U1697 ( .A(n527), .B(n362), .C(n519), .D(n441), .E(n168), .F(n526), 
        .G(n445), .H(intadd_3_SUM_3_), .Y(n900) );
  scg4d1_hd U1698 ( .A(n536), .B(n373), .C(n542), .D(n152), .E(b_m[8]), .F(
        n435), .G(n438), .H(n35), .Y(n901) );
  ivd1_hd U1699 ( .A(intadd_7_SUM_6_), .Y(intadd_5_A_9_) );
  scg4d1_hd U1700 ( .A(n552), .B(n150), .C(b_m[13]), .D(n226), .E(n548), .F(
        n427), .G(n1020), .H(intadd_3_SUM_9_), .Y(n902) );
  scg4d1_hd U1701 ( .A(n581), .B(n366), .C(n576), .D(n409), .E(n584), .F(n136), 
        .G(n414), .H(intadd_3_SUM_15_), .Y(n903) );
  fad1_hd U1702 ( .A(n905), .B(n904), .CI(intadd_5_SUM_8_), .CO(intadd_4_B_15_), .S(intadd_4_B_14_) );
  ivd1_hd U1703 ( .A(intadd_4_SUM_15_), .Y(n913) );
  ao21d1_hd U1704 ( .A(n396), .B(n76), .C(n906), .Y(n908) );
  nr2d1_hd U1705 ( .A(n200), .B(n908), .Y(n909) );
  scg4d1_hd U1706 ( .A(n594), .B(n131), .C(n591), .D(n401), .E(n601), .F(n223), 
        .G(n404), .H(n65), .Y(n910) );
  scg4d1_hd U1707 ( .A(n581), .B(n411), .C(n583), .D(n364), .E(n589), .F(n139), 
        .G(n413), .H(n64), .Y(n914) );
  scg4d1_hd U1708 ( .A(b_m[15]), .B(n418), .C(n570), .D(n369), .E(n577), .F(
        n140), .G(n423), .H(n52), .Y(n915) );
  scg4d1_hd U1709 ( .A(intadd_3_B_4_), .B(n166), .C(n524), .D(n441), .E(n534), 
        .F(n360), .G(n445), .H(intadd_3_SUM_4_), .Y(n916) );
  ivd1_hd U1710 ( .A(intadd_9_SUM_0_), .Y(intadd_12_B_1_) );
  scg4d1_hd U1711 ( .A(n547), .B(n153), .C(b_m[10]), .D(n374), .E(n435), .F(
        n539), .G(n438), .H(n40), .Y(n917) );
  scg4d1_hd U1712 ( .A(n552), .B(n426), .C(n556), .D(n145), .E(n562), .F(n227), 
        .G(n1020), .H(intadd_3_SUM_10_), .Y(n918) );
  ivd1_hd U1713 ( .A(intadd_7_SUM_7_), .Y(intadd_5_B_10_) );
  scg4d1_hd U1714 ( .A(n594), .B(n934), .C(n599), .D(n132), .E(n406), .F(n60), 
        .G(b_m[23]), .H(n224), .Y(n920) );
  ivd1_hd U1715 ( .A(intadd_9_B_2_), .Y(intadd_9_A_1_) );
  scg4d1_hd U1716 ( .A(intadd_3_B_4_), .B(n442), .C(n533), .D(n169), .E(n538), 
        .F(n363), .G(n445), .H(intadd_3_SUM_5_), .Y(n921) );
  ivd1_hd U1717 ( .A(intadd_9_SUM_1_), .Y(intadd_12_A_2_) );
  scg4d1_hd U1718 ( .A(n552), .B(n154), .C(n542), .D(n433), .E(n375), .F(n549), 
        .G(n438), .H(n42), .Y(n922) );
  scg4d1_hd U1719 ( .A(b_m[15]), .B(n228), .C(n556), .D(n425), .E(n147), .F(
        n562), .G(n431), .H(intadd_3_SUM_11_), .Y(n923) );
  scg4d1_hd U1720 ( .A(n580), .B(n144), .C(n572), .D(n416), .E(n368), .F(n577), 
        .G(n423), .H(n54), .Y(n924) );
  ivd1_hd U1721 ( .A(intadd_7_SUM_8_), .Y(intadd_5_A_11_) );
  scg4d1_hd U1722 ( .A(n594), .B(n137), .C(n583), .D(n408), .E(n367), .F(n590), 
        .G(n413), .H(intadd_3_SUM_17_), .Y(n925) );
  ao22d1_hd U1723 ( .A(b_m[22]), .B(n401), .C(n404), .D(n57), .Y(n926) );
  oa21d1_hd U1724 ( .A(n201), .B(n927), .C(n926), .Y(n928) );
  ivd1_hd U1725 ( .A(intadd_19_SUM_2_), .Y(intadd_0_A_20_) );
  ivd1_hd U1726 ( .A(intadd_4_n1), .Y(intadd_0_B_20_) );
  scg4d1_hd U1727 ( .A(n594), .B(n365), .C(n591), .D(n408), .E(n600), .F(n135), 
        .G(n412), .H(n66), .Y(n929) );
  ivd1_hd U1728 ( .A(intadd_5_n1), .Y(intadd_7_A_9_) );
  nr2d1_hd U1729 ( .A(n613), .B(n531), .Y(intadd_9_A_2_) );
  scg4d1_hd U1730 ( .A(n536), .B(n167), .C(n542), .D(n361), .E(b_m[8]), .F(
        n443), .G(n447), .H(intadd_3_SUM_6_), .Y(n930) );
  scg4d1_hd U1731 ( .A(n555), .B(n372), .C(n556), .D(n159), .E(n548), .F(n435), 
        .G(n438), .H(n44), .Y(n931) );
  ivd1_hd U1732 ( .A(intadd_18_SUM_0_), .Y(intadd_8_B_4_) );
  ivd1_hd U1733 ( .A(intadd_8_SUM_4_), .Y(intadd_17_A_0_) );
  scg4d1_hd U1734 ( .A(n565), .B(n149), .C(n561), .D(n1019), .E(n572), .F(n359), .G(n431), .H(intadd_3_SUM_12_), .Y(n932) );
  scg4d1_hd U1735 ( .A(n580), .B(n370), .C(n575), .D(n417), .E(n584), .F(n142), 
        .G(n993), .H(n56), .Y(n933) );
  ivd1_hd U1736 ( .A(intadd_17_SUM_0_), .Y(intadd_7_B_9_) );
  ivd1_hd U1737 ( .A(intadd_7_SUM_9_), .Y(n948) );
  ao21d1_hd U1738 ( .A(n1063), .B(n404), .C(n401), .Y(n936) );
  nr2d1_hd U1739 ( .A(n201), .B(n936), .Y(n937) );
  ivd1_hd U1740 ( .A(n938), .Y(intadd_0_A_21_) );
  ivd1_hd U1741 ( .A(intadd_19_n1), .Y(intadd_0_B_21_) );
  scg4d1_hd U1742 ( .A(n547), .B(n362), .C(intadd_3_B_7_), .D(n168), .E(n443), 
        .F(n539), .G(n447), .H(intadd_3_SUM_7_), .Y(n939) );
  nr2bd1_hd U1743 ( .AN(n940), .B(intadd_9_A_2_), .Y(n952) );
  nr2d1_hd U1744 ( .A(n531), .B(n940), .Y(n951) );
  nr2d1_hd U1745 ( .A(n952), .B(n951), .Y(n941) );
  scg4d1_hd U1746 ( .A(n555), .B(n434), .C(b_m[13]), .D(n373), .E(n561), .F(
        n152), .G(n437), .H(n46), .Y(n942) );
  ivd1_hd U1747 ( .A(intadd_18_SUM_1_), .Y(intadd_8_A_5_) );
  scg4d1_hd U1748 ( .A(n565), .B(n426), .C(n572), .D(n150), .E(n577), .F(n226), 
        .G(n431), .H(intadd_3_SUM_13_), .Y(n943) );
  ivd1_hd U1749 ( .A(intadd_8_SUM_5_), .Y(intadd_17_A_1_) );
  scg4d1_hd U1750 ( .A(n580), .B(n419), .C(n583), .D(n371), .E(n589), .F(n143), 
        .G(n423), .H(intadd_3_SUM_16_), .Y(n944) );
  ivd1_hd U1751 ( .A(intadd_17_SUM_1_), .Y(intadd_7_A_10_) );
  scg4d1_hd U1752 ( .A(n594), .B(n411), .C(n600), .D(n366), .E(b_m[23]), .F(
        n136), .G(n412), .H(n1046), .Y(n946) );
  ivd1_hd U1753 ( .A(intadd_11_A_0_), .Y(n962) );
  scg20d1_hd U1754 ( .A(n606), .B(n952), .C(n951), .Y(n961) );
  scg4d1_hd U1755 ( .A(n552), .B(n363), .C(intadd_3_B_7_), .D(n441), .E(n169), 
        .F(n549), .G(n1064), .H(intadd_3_SUM_8_), .Y(n953) );
  scg4d1_hd U1756 ( .A(n565), .B(n153), .C(n556), .D(n433), .E(n374), .F(n563), 
        .G(n439), .H(n50), .Y(n954) );
  scg4d1_hd U1757 ( .A(n580), .B(n227), .C(b_m[16]), .D(n424), .E(n145), .F(
        n577), .G(n431), .H(intadd_3_SUM_14_), .Y(n955) );
  ivd1_hd U1758 ( .A(intadd_18_SUM_2_), .Y(intadd_8_A_6_) );
  scg4d1_hd U1759 ( .A(n594), .B(n144), .C(n585), .D(n416), .E(n368), .F(
        b_m[20]), .G(n420), .H(intadd_3_SUM_17_), .Y(n956) );
  ivd1_hd U1760 ( .A(intadd_8_SUM_6_), .Y(intadd_17_A_2_) );
  ao22d1_hd U1761 ( .A(b_m[22]), .B(n408), .C(n412), .D(n58), .Y(n957) );
  oa21d1_hd U1762 ( .A(n202), .B(n945), .C(n957), .Y(n958) );
  scg4d1_hd U1763 ( .A(n593), .B(n369), .C(n591), .D(n416), .E(n600), .F(n140), 
        .G(n421), .H(n65), .Y(n959) );
  ivd1_hd U1764 ( .A(intadd_18_n1), .Y(intadd_8_A_7_) );
  fad1_hd U1765 ( .A(n962), .B(n961), .CI(n960), .CO(intadd_9_A_5_), .S(
        intadd_9_A_4_) );
  nr2d1_hd U1766 ( .A(n613), .B(n545), .Y(intadd_11_B_0_) );
  scg4d1_hd U1767 ( .A(n555), .B(n166), .C(n556), .D(n360), .E(n548), .F(n443), 
        .G(n1064), .H(intadd_3_SUM_9_), .Y(n963) );
  ivd1_hd U1768 ( .A(intadd_11_SUM_0_), .Y(intadd_9_B_5_) );
  scg4d1_hd U1769 ( .A(b_m[15]), .B(n375), .C(n561), .D(n432), .E(n571), .F(
        n154), .G(n439), .H(n48), .Y(n964) );
  scg4d1_hd U1770 ( .A(n580), .B(n147), .C(n576), .D(n425), .E(n585), .F(n228), 
        .G(n1020), .H(intadd_3_SUM_15_), .Y(n965) );
  ivd1_hd U1771 ( .A(intadd_16_SUM_0_), .Y(intadd_8_B_7_) );
  ivd1_hd U1772 ( .A(intadd_8_SUM_7_), .Y(n979) );
  ao21d1_hd U1773 ( .A(n412), .B(n76), .C(n408), .Y(n968) );
  nr2d1_hd U1774 ( .A(n200), .B(n968), .Y(n969) );
  scg4d1_hd U1775 ( .A(n555), .B(n442), .C(intadd_3_B_10_), .D(n167), .E(n561), 
        .F(n362), .G(n1064), .H(intadd_3_SUM_10_), .Y(n971) );
  nr2d1_hd U1776 ( .A(intadd_3_B_8_), .B(intadd_3_B_6_), .Y(n972) );
  ao211d1_hd U1777 ( .A(intadd_3_B_8_), .B(intadd_3_B_6_), .C(n610), .D(n972), 
        .Y(n973) );
  ivd1_hd U1778 ( .A(intadd_11_SUM_1_), .Y(intadd_9_A_6_) );
  scg4d1_hd U1779 ( .A(n565), .B(n434), .C(n570), .D(n373), .E(n576), .F(n152), 
        .G(n439), .H(n52), .Y(n974) );
  scg4d1_hd U1780 ( .A(n579), .B(n427), .C(b_m[19]), .D(n150), .E(n590), .F(
        n226), .G(n428), .H(n64), .Y(n975) );
  ivd1_hd U1781 ( .A(intadd_16_SUM_1_), .Y(intadd_8_A_8_) );
  scg4d1_hd U1782 ( .A(n593), .B(n419), .C(n599), .D(n370), .E(n108), .F(n142), 
        .G(n421), .H(n60), .Y(n977) );
  ivd1_hd U1783 ( .A(intadd_10_B_1_), .Y(intadd_10_A_0_) );
  nr2d1_hd U1784 ( .A(n193), .B(intadd_11_A_0_), .Y(n983) );
  ao211d1_hd U1785 ( .A(n193), .B(n541), .C(n610), .D(n551), .Y(n982) );
  nr2d1_hd U1786 ( .A(n983), .B(n982), .Y(intadd_10_B_0_) );
  scg4d1_hd U1787 ( .A(n565), .B(n361), .C(intadd_3_B_10_), .D(n441), .E(n168), 
        .F(n563), .G(n446), .H(intadd_3_SUM_11_), .Y(n984) );
  ivd1_hd U1788 ( .A(intadd_10_SUM_0_), .Y(intadd_11_A_2_) );
  scg4d1_hd U1789 ( .A(n579), .B(n159), .C(b_m[16]), .D(n432), .E(n372), .F(
        n578), .G(n439), .H(n54), .Y(n985) );
  ivd1_hd U1790 ( .A(intadd_11_SUM_2_), .Y(intadd_9_A_7_) );
  scg4d1_hd U1791 ( .A(n593), .B(n359), .C(n585), .D(n424), .E(n149), .F(
        b_m[20]), .G(n431), .H(n62), .Y(n986) );
  ao22d1_hd U1792 ( .A(b_m[22]), .B(n416), .C(n421), .D(n57), .Y(n987) );
  oa21d1_hd U1793 ( .A(n201), .B(n976), .C(n987), .Y(n988) );
  scg4d1_hd U1794 ( .A(n593), .B(n145), .C(n591), .D(n424), .E(n601), .F(n227), 
        .G(n429), .H(n66), .Y(n989) );
  ivd1_hd U1795 ( .A(intadd_9_n1), .Y(intadd_11_A_3_) );
  scg4d1_hd U1796 ( .A(intadd_3_B_12_), .B(n169), .C(n564), .D(n440), .E(n572), 
        .F(n363), .G(n446), .H(intadd_3_SUM_12_), .Y(n990) );
  scg4d1_hd U1797 ( .A(n579), .B(n374), .C(n576), .D(n433), .E(n584), .F(n153), 
        .G(n437), .H(n56), .Y(n991) );
  nr2d1_hd U1798 ( .A(n613), .B(n560), .Y(intadd_10_A_1_) );
  ivd1_hd U1799 ( .A(intadd_15_SUM_0_), .Y(intadd_11_B_3_) );
  ivd1_hd U1800 ( .A(intadd_11_SUM_3_), .Y(n1004) );
  ao21d1_hd U1801 ( .A(n421), .B(n1063), .C(n992), .Y(n994) );
  nr2d1_hd U1802 ( .A(n107), .B(n994), .Y(n995) );
  scg4d1_hd U1803 ( .A(intadd_3_B_12_), .B(n442), .C(b_m[16]), .D(n166), .E(
        n576), .F(n360), .G(n446), .H(intadd_3_SUM_13_), .Y(n997) );
  nr2bd1_hd U1804 ( .AN(n998), .B(intadd_10_A_1_), .Y(n1008) );
  nr2d1_hd U1805 ( .A(n560), .B(n998), .Y(n1007) );
  nr2d1_hd U1806 ( .A(n1008), .B(n1007), .Y(n999) );
  scg4d1_hd U1807 ( .A(n579), .B(n435), .C(n583), .D(n375), .E(n590), .F(n154), 
        .G(n439), .H(intadd_3_SUM_16_), .Y(n1000) );
  ivd1_hd U1808 ( .A(intadd_15_SUM_1_), .Y(intadd_11_A_4_) );
  scg4d1_hd U1809 ( .A(n593), .B(n427), .C(n599), .D(n147), .E(n1112), .F(n228), .G(n429), .H(n1046), .Y(n1002) );
  nr2d1_hd U1810 ( .A(n614), .B(n569), .Y(n1017) );
  scg20d1_hd U1811 ( .A(n110), .B(n1008), .C(n1007), .Y(n1016) );
  scg4d1_hd U1812 ( .A(n580), .B(n361), .C(b_m[16]), .D(n440), .E(n167), .F(
        n578), .G(n446), .H(intadd_3_SUM_14_), .Y(n1009) );
  scg4d1_hd U1813 ( .A(n592), .B(n159), .C(b_m[19]), .D(n432), .E(n372), .F(
        b_m[20]), .G(n1040), .H(intadd_3_SUM_17_), .Y(n1010) );
  ao22d1_hd U1814 ( .A(n598), .B(n424), .C(n429), .D(n58), .Y(n1011) );
  oa21d1_hd U1815 ( .A(n202), .B(n1012), .C(n1011), .Y(n1013) );
  scg4d1_hd U1816 ( .A(n592), .B(n373), .C(n589), .D(n432), .E(n601), .F(n152), 
        .G(n436), .H(n65), .Y(n1014) );
  fad1_hd U1817 ( .A(n1017), .B(n1016), .CI(n1015), .CO(intadd_10_A_4_), .S(
        intadd_10_A_3_) );
  ivd1_hd U1818 ( .A(n1017), .Y(intadd_13_A_0_) );
  nr2d1_hd U1819 ( .A(n614), .B(n573), .Y(intadd_13_B_0_) );
  scg4d1_hd U1820 ( .A(b_m[18]), .B(n168), .C(n575), .D(n441), .E(n585), .F(
        n362), .G(n1064), .H(intadd_3_SUM_15_), .Y(n1018) );
  ivd1_hd U1821 ( .A(intadd_13_SUM_0_), .Y(intadd_10_B_4_) );
  ao21d1_hd U1822 ( .A(n429), .B(n76), .C(n1019), .Y(n1021) );
  nr2d1_hd U1823 ( .A(n200), .B(n1021), .Y(n1022) );
  ivd1_hd U1824 ( .A(n1023), .Y(intadd_0_A_30_) );
  ivd1_hd U1825 ( .A(intadd_15_n1), .Y(intadd_0_B_30_) );
  scg4d1_hd U1826 ( .A(b_m[18]), .B(n443), .C(b_m[19]), .D(n169), .E(n590), 
        .F(n363), .G(n446), .H(n64), .Y(n1024) );
  nr2d1_hd U1827 ( .A(n569), .B(n1025), .Y(n1032) );
  nr2bd1_hd U1828 ( .AN(n1033), .B(n1032), .Y(n1026) );
  ivd1_hd U1829 ( .A(intadd_13_SUM_1_), .Y(intadd_10_A_5_) );
  scg4d1_hd U1830 ( .A(n593), .B(n435), .C(n600), .D(n374), .E(b_m[23]), .F(
        n153), .G(n436), .H(n60), .Y(n1028) );
  fad1_hd U1831 ( .A(n1030), .B(intadd_10_SUM_4_), .CI(n1029), .CO(n1031), .S(
        n1023) );
  ivd1_hd U1832 ( .A(intadd_14_B_1_), .Y(intadd_14_A_0_) );
  ao21d1_hd U1833 ( .A(n460), .B(n1033), .C(n1032), .Y(intadd_14_B_0_) );
  ivd1_hd U1834 ( .A(intadd_14_SUM_0_), .Y(intadd_13_A_2_) );
  ao22d1_hd U1835 ( .A(b_m[22]), .B(n1039), .C(n436), .D(n57), .Y(n1035) );
  oa21d1_hd U1836 ( .A(n200), .B(n1027), .C(n1035), .Y(n1036) );
  scg4d1_hd U1837 ( .A(n592), .B(n167), .C(n589), .D(n1062), .E(n601), .F(n361), .G(n444), .H(n66), .Y(n1038) );
  nr2d1_hd U1838 ( .A(n614), .B(n587), .Y(intadd_14_A_1_) );
  ao21d1_hd U1839 ( .A(n436), .B(n1063), .C(n432), .Y(n1041) );
  nr2d1_hd U1840 ( .A(n202), .B(n1041), .Y(n1042) );
  nr2bd1_hd U1841 ( .AN(n1044), .B(intadd_14_A_1_), .Y(n1057) );
  nr2d1_hd U1842 ( .A(n587), .B(n1044), .Y(n1056) );
  nr2d1_hd U1843 ( .A(n1057), .B(n1056), .Y(n1045) );
  scg4d1_hd U1844 ( .A(n592), .B(n443), .C(n600), .D(n168), .E(n108), .F(n362), 
        .G(n444), .H(n1046), .Y(n1049) );
  ivd1_hd U1845 ( .A(intadd_14_SUM_2_), .Y(intadd_0_A_34_) );
  ivd1_hd U1846 ( .A(n1052), .Y(intadd_0_B_34_) );
  ao22d1_hd U1847 ( .A(n598), .B(n1062), .C(n444), .D(n58), .Y(n1054) );
  oa21d1_hd U1848 ( .A(n200), .B(n1048), .C(n1054), .Y(n1055) );
  scg20d1_hd U1849 ( .A(a_m[20]), .B(n1057), .C(n1056), .Y(n1059) );
  fad1_hd U1850 ( .A(n1060), .B(n1073), .CI(n1059), .CO(n1061), .S(n1058) );
  ao21d1_hd U1851 ( .A(n444), .B(n76), .C(n1062), .Y(n1065) );
  nr2d1_hd U1852 ( .A(n201), .B(n1065), .Y(n1067) );
  oa21d1_hd U1853 ( .A(n617), .B(n1067), .C(n1070), .Y(n1072) );
  scg16d1_hd U1854 ( .A(n1070), .B(n1069), .C(n1068), .Y(intadd_0_B_36_) );
  oa211d1_hd U1855 ( .A(n597), .B(n1070), .C(n617), .D(n599), .Y(n1071) );
  oa21d1_hd U1856 ( .A(n1073), .B(n1072), .C(n1071), .Y(n1076) );
  oa211d1_hd U1857 ( .A(intadd_3_A_17_), .B(n202), .C(n617), .D(n1074), .Y(
        n1075) );
  ivd1_hd U1858 ( .A(b_e[9]), .Y(n1415) );
  ivd1_hd U1859 ( .A(a_e[9]), .Y(n1355) );
  ao22d1_hd U1860 ( .A(a_e[9]), .B(b_e[9]), .C(n1415), .D(n1355), .Y(n1079) );
  nr2d1_hd U1861 ( .A(DP_OP_125J2_130_6300_n12), .B(n1079), .Y(n1078) );
  ao211d1_hd U1862 ( .A(DP_OP_125J2_130_6300_n12), .B(n1079), .C(n497), .D(
        n1078), .Y(n1080) );
  ao21d1_hd U1863 ( .A(z_e[9]), .B(n90), .C(n1080), .Y(n1081) );
  ivd1_hd U1864 ( .A(n1183), .Y(n3279) );
  ao21d1_hd U1865 ( .A(n456), .B(product[25]), .C(n1083), .Y(n104) );
  nr2d1_hd U1866 ( .A(z_e[4]), .B(z_e[3]), .Y(n1085) );
  nr2d1_hd U1867 ( .A(z_e[6]), .B(z_e[5]), .Y(n1084) );
  nr3d1_hd U1868 ( .A(z_e[2]), .B(z_e[1]), .C(n1141), .Y(n1086) );
  oa21d1_hd U1869 ( .A(n1086), .B(n1140), .C(z_e[9]), .Y(n36) );
  ao22d1_hd U1870 ( .A(n481), .B(a[23]), .C(n102), .D(a_e[0]), .Y(n1348) );
  ivd1_hd U1871 ( .A(n1348), .Y(n1206) );
  ao22d1_hd U1872 ( .A(n481), .B(b[23]), .C(b_e[0]), .D(n106), .Y(n1363) );
  ivd1_hd U1873 ( .A(n1363), .Y(n1207) );
  nr4d1_hd U1874 ( .A(a_e[2]), .B(n10), .C(a_e[6]), .D(n1088), .Y(n1089) );
  ivd1_hd U1875 ( .A(n1089), .Y(n1090) );
  nr4d1_hd U1876 ( .A(a_e[0]), .B(a_e[9]), .C(a_e[8]), .D(n1090), .Y(n1132) );
  nr4d1_hd U1877 ( .A(n1091), .B(b_e[2]), .C(b_e[5]), .D(b_e[4]), .Y(n1101) );
  ivd1_hd U1878 ( .A(n1101), .Y(n1092) );
  nr4d1_hd U1879 ( .A(b_e[8]), .B(b_e[9]), .C(b_e[0]), .D(n1092), .Y(n1130) );
  nr2d1_hd U1880 ( .A(n1132), .B(n1130), .Y(n1139) );
  nd4d1_hd U1881 ( .A(n1094), .B(n1093), .C(n1366), .D(n1376), .Y(n1100) );
  nr4d1_hd U1882 ( .A(a_m[4]), .B(a_m[3]), .C(a_m[2]), .D(a_m[0]), .Y(n1098)
         );
  nr4d1_hd U1883 ( .A(a_m[1]), .B(a_m[12]), .C(a_m[17]), .D(n203), .Y(n1097)
         );
  nr4d1_hd U1884 ( .A(a_m[6]), .B(n111), .C(a_m[10]), .D(n86), .Y(n1096) );
  nr4d1_hd U1885 ( .A(a_m[16]), .B(a_m[15]), .C(n193), .D(a_m[9]), .Y(n1095)
         );
  nd4d1_hd U1886 ( .A(n1098), .B(n1097), .C(n1096), .D(n1095), .Y(n1099) );
  nr4d1_hd U1887 ( .A(a_m[18]), .B(a_m[21]), .C(n1100), .D(n1099), .Y(n1126)
         );
  nr2d1_hd U1888 ( .A(intadd_3_B_0_), .B(n503), .Y(n1102) );
  nd4d1_hd U1889 ( .A(n1103), .B(n1102), .C(n596), .D(n201), .Y(n1109) );
  nr4d1_hd U1890 ( .A(intadd_3_B_9_), .B(intadd_3_B_8_), .C(intadd_3_B_4_), 
        .D(intadd_3_B_6_), .Y(n1107) );
  nr4d1_hd U1891 ( .A(intadd_3_B_5_), .B(intadd_3_B_1_), .C(intadd_3_B_3_), 
        .D(intadd_3_B_2_), .Y(n1106) );
  nr4d1_hd U1892 ( .A(intadd_3_B_13_), .B(intadd_3_B_11_), .C(intadd_3_B_10_), 
        .D(intadd_3_B_7_), .Y(n1105) );
  nr4d1_hd U1893 ( .A(intadd_3_B_17_), .B(intadd_3_B_16_), .C(intadd_3_B_12_), 
        .D(b_m[17]), .Y(n1104) );
  nd4d1_hd U1894 ( .A(n1107), .B(n1106), .C(n1105), .D(n1104), .Y(n1108) );
  nr4d1_hd U1895 ( .A(n598), .B(intadd_3_B_15_), .C(n1109), .D(n1108), .Y(
        n1128) );
  nr2d1_hd U1896 ( .A(n1349), .B(n10), .Y(n1343) );
  ivd1_hd U1897 ( .A(n1343), .Y(n1341) );
  ivd1_hd U1898 ( .A(DP_OP_113J2_124_6892_n3), .Y(n1342) );
  ao22d1_hd U1899 ( .A(DP_OP_113J2_124_6892_n3), .B(n1341), .C(n1343), .D(
        n1342), .Y(n1110) );
  ao22d1_hd U1900 ( .A(n79), .B(a_e[7]), .C(n78), .D(n1110), .Y(n141) );
  ao22d1_hd U1901 ( .A(n480), .B(b[30]), .C(n103), .D(b_e[7]), .Y(n1356) );
  ao22d1_hd U1902 ( .A(n83), .B(b_e[7]), .C(n82), .D(n1113), .Y(n151) );
  nr3d1_hd U1903 ( .A(n1114), .B(n101), .C(n495), .Y(n156) );
  oa211d1_hd U1904 ( .A(n1118), .B(n73), .C(n1117), .D(n1143), .Y(n1119) );
  nr2d1_hd U1905 ( .A(n1222), .B(n1119), .Y(n160) );
  nr2d1_hd U1906 ( .A(n1121), .B(n1120), .Y(n161) );
  nr2d1_hd U1907 ( .A(n454), .B(n89), .Y(n171) );
  ao22d1_hd U1908 ( .A(z_m[23]), .B(n376), .C(n475), .D(n177), .Y(n172) );
  ao22d1_hd U1909 ( .A(n101), .B(n618), .C(n1112), .D(n106), .Y(n173) );
  nr2d1_hd U1910 ( .A(n475), .B(o_Z_STB), .Y(n179) );
  ao22d1_hd U1911 ( .A(n1132), .B(n1131), .C(n1130), .D(n1129), .Y(n1133) );
  nr2d1_hd U1912 ( .A(n1133), .B(n1138), .Y(n1175) );
  ao22d1_hd U1913 ( .A(n1134), .B(b_s), .C(n1174), .D(z_s), .Y(n1135) );
  nr2d1_hd U1914 ( .A(z_e[1]), .B(z_e[0]), .Y(n1167) );
  ivd1_hd U1915 ( .A(z_e[2]), .Y(n1163) );
  nr2d1_hd U1916 ( .A(z_e[3]), .B(n1162), .Y(n1159) );
  ivd1_hd U1917 ( .A(z_e[4]), .Y(n1156) );
  nr2d1_hd U1918 ( .A(z_e[5]), .B(n1155), .Y(n1152) );
  ivd1_hd U1919 ( .A(z_e[6]), .Y(n1149) );
  nr2d1_hd U1920 ( .A(z_m[23]), .B(z_e[0]), .Y(n1145) );
  ivd1_hd U1921 ( .A(z_e[1]), .Y(n1142) );
  nr4d1_hd U1922 ( .A(z_e[2]), .B(n1142), .C(n1141), .D(n1140), .Y(n1144) );
  ao21d1_hd U1923 ( .A(n1145), .B(n1144), .C(n1143), .Y(n1165) );
  oa211d1_hd U1924 ( .A(z_e[7]), .B(n1148), .C(n1165), .D(n1146), .Y(n1147) );
  scg15d1_hd U1925 ( .A(n1178), .B(z[30]), .C(n1171), .D(n1147), .Y(n230) );
  oa21d1_hd U1926 ( .A(n1152), .B(n1149), .C(n1148), .Y(n1150) );
  ao22d1_hd U1927 ( .A(n452), .B(z[29]), .C(n1165), .D(n1150), .Y(n1151) );
  ao21d1_hd U1928 ( .A(z_e[5]), .B(n1155), .C(n1152), .Y(n1154) );
  oa211d1_hd U1929 ( .A(n1154), .B(n1172), .C(n1171), .D(n1153), .Y(n232) );
  oa21d1_hd U1930 ( .A(n1159), .B(n1156), .C(n1155), .Y(n1157) );
  ao22d1_hd U1931 ( .A(n452), .B(z[27]), .C(n1165), .D(n1157), .Y(n1158) );
  ao21d1_hd U1932 ( .A(z_e[3]), .B(n1162), .C(n1159), .Y(n1161) );
  oa211d1_hd U1933 ( .A(n1161), .B(n1172), .C(n1171), .D(n1160), .Y(n234) );
  oa21d1_hd U1934 ( .A(n1167), .B(n1163), .C(n1162), .Y(n1164) );
  ao22d1_hd U1935 ( .A(n451), .B(z[25]), .C(n1165), .D(n1164), .Y(n1166) );
  ao21d1_hd U1936 ( .A(z_e[0]), .B(z_e[1]), .C(n1167), .Y(n1169) );
  oa211d1_hd U1937 ( .A(n1169), .B(n1172), .C(n1171), .D(n1168), .Y(n236) );
  oa211d1_hd U1938 ( .A(z_e[0]), .B(n1172), .C(n1171), .D(n1170), .Y(n237) );
  ao21d1_hd U1939 ( .A(n451), .B(z[22]), .C(n1175), .Y(n1176) );
  oa21d1_hd U1940 ( .A(n1306), .B(n1177), .C(n1176), .Y(n238) );
  nr2d1_hd U1941 ( .A(sticky), .B(round_bit), .Y(n1179) );
  nd3d1_hd U1942 ( .A(n1269), .B(z_m[4]), .C(z_m[3]), .Y(n1257) );
  ivd1_hd U1943 ( .A(n1257), .Y(n1258) );
  ivd1_hd U1944 ( .A(z_m[5]), .Y(n1261) );
  nd3d1_hd U1945 ( .A(n1249), .B(z_m[8]), .C(z_m[7]), .Y(n1239) );
  ivd1_hd U1946 ( .A(n1239), .Y(n1240) );
  ivd1_hd U1947 ( .A(z_m[9]), .Y(n1243) );
  nd3d1_hd U1948 ( .A(n1232), .B(z_m[12]), .C(n17), .Y(n1221) );
  ivd1_hd U1949 ( .A(n1221), .Y(n1223) );
  nd3d1_hd U1950 ( .A(n1223), .B(z_m[14]), .C(z_m[13]), .Y(n1204) );
  ivd1_hd U1951 ( .A(n1204), .Y(n1205) );
  nd3d1_hd U1952 ( .A(n1205), .B(z_m[16]), .C(n19), .Y(n1195) );
  ivd1_hd U1953 ( .A(n1195), .Y(n1196) );
  nd3d1_hd U1954 ( .A(n1196), .B(z_m[18]), .C(z_m[17]), .Y(n1186) );
  ivd1_hd U1955 ( .A(n1186), .Y(n1187) );
  nd3d1_hd U1956 ( .A(n1187), .B(z_m[20]), .C(n21), .Y(n1304) );
  ao21d1_hd U1957 ( .A(n199), .B(n1304), .C(n95), .Y(n1182) );
  oa21d1_hd U1958 ( .A(z_m[21]), .B(n98), .C(n1182), .Y(n1301) );
  nd2bd1_hd U1959 ( .AN(n1304), .B(n199), .Y(n1181) );
  oa21d1_hd U1960 ( .A(z_m[22]), .B(n1181), .C(n194), .Y(n1180) );
  scg4d1_hd U1961 ( .A(n1301), .B(z_m[22]), .C(n1180), .D(z_m[21]), .E(z_m[23]), .F(n1290), .G(n458), .H(product[48]), .Y(n261) );
  ivd1_hd U1962 ( .A(z_m[21]), .Y(n1305) );
  ao22d1_hd U1963 ( .A(z_m[21]), .B(n1182), .C(n1181), .D(n1305), .Y(n1185) );
  ao22d1_hd U1964 ( .A(n456), .B(product[47]), .C(z_m[22]), .D(n185), .Y(n1184) );
  oa21d1_hd U1965 ( .A(n96), .B(n1186), .C(n1256), .Y(n1190) );
  oa21d1_hd U1966 ( .A(n21), .B(n97), .C(n1190), .Y(n1189) );
  oa21d1_hd U1967 ( .A(z_m[20]), .B(n1194), .C(n194), .Y(n1188) );
  scg4d1_hd U1968 ( .A(n1189), .B(z_m[20]), .C(n1188), .D(z_m[19]), .E(z_m[21]), .F(n185), .G(n1303), .H(product[46]), .Y(n263) );
  ao22d1_hd U1969 ( .A(n456), .B(product[45]), .C(z_m[20]), .D(n184), .Y(n1193) );
  ivd1_hd U1970 ( .A(n1190), .Y(n1191) );
  ao22d1_hd U1971 ( .A(z_m[18]), .B(n99), .C(n21), .D(n1191), .Y(n1192) );
  oa211d1_hd U1972 ( .A(n21), .B(n1194), .C(n1193), .D(n1192), .Y(n264) );
  ao21d1_hd U1973 ( .A(n1222), .B(n1195), .C(n95), .Y(n1201) );
  oa21d1_hd U1974 ( .A(z_m[17]), .B(n98), .C(n1201), .Y(n1198) );
  oa21d1_hd U1975 ( .A(z_m[18]), .B(n1200), .C(n195), .Y(n1197) );
  scg4d1_hd U1976 ( .A(n1198), .B(z_m[18]), .C(n1197), .D(n190), .E(n21), .F(
        n183), .G(n1303), .H(product[44]), .Y(n265) );
  ivd1_hd U1977 ( .A(z_m[17]), .Y(n1199) );
  ao22d1_hd U1978 ( .A(z_m[17]), .B(n1201), .C(n1200), .D(n1199), .Y(n1203) );
  ao22d1_hd U1979 ( .A(n457), .B(product[43]), .C(z_m[18]), .D(n184), .Y(n1202) );
  oa21d1_hd U1980 ( .A(n95), .B(n1204), .C(n1256), .Y(n1216) );
  oa21d1_hd U1981 ( .A(n19), .B(n98), .C(n1216), .Y(n1215) );
  oa21d1_hd U1982 ( .A(z_m[16]), .B(n1220), .C(n195), .Y(n1214) );
  scg4d1_hd U1983 ( .A(n1215), .B(z_m[16]), .C(n1214), .D(z_m[15]), .E(n190), 
        .F(n184), .G(n455), .H(product[42]), .Y(n267) );
  ao22d1_hd U1984 ( .A(n457), .B(product[41]), .C(z_m[16]), .D(n183), .Y(n1219) );
  ivd1_hd U1985 ( .A(n1216), .Y(n1217) );
  ao22d1_hd U1986 ( .A(z_m[14]), .B(n100), .C(n19), .D(n1217), .Y(n1218) );
  oa211d1_hd U1987 ( .A(n19), .B(n1220), .C(n1219), .D(n1218), .Y(n268) );
  ao21d1_hd U1988 ( .A(n1222), .B(n1221), .C(n96), .Y(n1228) );
  oa21d1_hd U1989 ( .A(z_m[13]), .B(n97), .C(n1228), .Y(n1225) );
  oa21d1_hd U1990 ( .A(z_m[14]), .B(n1227), .C(n194), .Y(n1224) );
  scg4d1_hd U1991 ( .A(n1225), .B(z_m[14]), .C(n1224), .D(n189), .E(n19), .F(
        n186), .G(n455), .H(product[40]), .Y(n269) );
  ivd1_hd U1992 ( .A(z_m[13]), .Y(n1226) );
  ao22d1_hd U1993 ( .A(z_m[13]), .B(n1228), .C(n1227), .D(n1226), .Y(n1230) );
  ao22d1_hd U1994 ( .A(n456), .B(product[39]), .C(z_m[14]), .D(n183), .Y(n1229) );
  oa21d1_hd U1995 ( .A(n1267), .B(n1232), .C(n1266), .Y(n1235) );
  ivd1_hd U1996 ( .A(n1235), .Y(n1231) );
  oa21d1_hd U1997 ( .A(n17), .B(n97), .C(n1231), .Y(n1234) );
  oa21d1_hd U1998 ( .A(z_m[12]), .B(n1238), .C(n195), .Y(n1233) );
  scg4d1_hd U1999 ( .A(n1234), .B(z_m[12]), .C(n1233), .D(z_m[11]), .E(n189), 
        .F(n183), .G(n455), .H(product[38]), .Y(n271) );
  ao22d1_hd U2000 ( .A(n457), .B(product[37]), .C(z_m[12]), .D(n185), .Y(n1237) );
  ao22d1_hd U2001 ( .A(z_m[10]), .B(n99), .C(n17), .D(n1235), .Y(n1236) );
  oa211d1_hd U2002 ( .A(n17), .B(n1238), .C(n1237), .D(n1236), .Y(n272) );
  oa21d1_hd U2003 ( .A(n96), .B(n1239), .C(n1256), .Y(n1245) );
  oa21d1_hd U2004 ( .A(z_m[9]), .B(n98), .C(n1245), .Y(n1242) );
  oa21d1_hd U2005 ( .A(z_m[10]), .B(n1244), .C(n195), .Y(n1241) );
  scg4d1_hd U2006 ( .A(n1242), .B(z_m[10]), .C(n1241), .D(z_m[9]), .E(n17), 
        .F(n183), .G(n1303), .H(product[36]), .Y(n273) );
  ao22d1_hd U2007 ( .A(z_m[9]), .B(n1245), .C(n1244), .D(n1243), .Y(n1247) );
  ao22d1_hd U2008 ( .A(n458), .B(product[35]), .C(z_m[10]), .D(n186), .Y(n1246) );
  oa21d1_hd U2009 ( .A(n1267), .B(n1249), .C(n1266), .Y(n1252) );
  ivd1_hd U2010 ( .A(n1252), .Y(n1248) );
  oa21d1_hd U2011 ( .A(z_m[7]), .B(n97), .C(n1248), .Y(n1251) );
  oa21d1_hd U2012 ( .A(z_m[8]), .B(n1255), .C(n194), .Y(n1250) );
  scg4d1_hd U2013 ( .A(n1251), .B(z_m[8]), .C(n1250), .D(z_m[7]), .E(z_m[9]), 
        .F(n186), .G(n455), .H(product[34]), .Y(n275) );
  ao22d1_hd U2014 ( .A(n457), .B(product[33]), .C(z_m[8]), .D(n186), .Y(n1254)
         );
  ao22d1_hd U2015 ( .A(z_m[6]), .B(n99), .C(z_m[7]), .D(n1252), .Y(n1253) );
  oa211d1_hd U2016 ( .A(n187), .B(n1255), .C(n1254), .D(n1253), .Y(n276) );
  oa21d1_hd U2017 ( .A(n95), .B(n1257), .C(n1256), .Y(n1263) );
  oa21d1_hd U2018 ( .A(z_m[5]), .B(n98), .C(n1263), .Y(n1260) );
  oa21d1_hd U2019 ( .A(z_m[6]), .B(n1262), .C(n194), .Y(n1259) );
  scg4d1_hd U2020 ( .A(n1260), .B(z_m[6]), .C(n1259), .D(z_m[5]), .E(n187), 
        .F(n185), .G(n1303), .H(product[32]), .Y(n277) );
  ao22d1_hd U2021 ( .A(z_m[5]), .B(n1263), .C(n1262), .D(n1261), .Y(n1265) );
  ao22d1_hd U2022 ( .A(n458), .B(product[31]), .C(z_m[6]), .D(n185), .Y(n1264)
         );
  oa21d1_hd U2023 ( .A(n1267), .B(n1269), .C(n1266), .Y(n1272) );
  ivd1_hd U2024 ( .A(n1272), .Y(n1268) );
  oa21d1_hd U2025 ( .A(z_m[3]), .B(n97), .C(n1268), .Y(n1271) );
  oa21d1_hd U2026 ( .A(z_m[4]), .B(n1275), .C(n195), .Y(n1270) );
  scg4d1_hd U2027 ( .A(n1271), .B(z_m[4]), .C(n1270), .D(z_m[3]), .E(z_m[5]), 
        .F(n184), .G(n458), .H(product[30]), .Y(n279) );
  ao22d1_hd U2028 ( .A(n457), .B(product[29]), .C(z_m[4]), .D(n184), .Y(n1274)
         );
  ao22d1_hd U2029 ( .A(z_m[2]), .B(n100), .C(z_m[3]), .D(n1272), .Y(n1273) );
  oa211d1_hd U2030 ( .A(n188), .B(n1275), .C(n1274), .D(n1273), .Y(n280) );
  nr2d1_hd U2031 ( .A(n23), .B(n97), .Y(n1297) );
  nr2d1_hd U2032 ( .A(n96), .B(n1297), .Y(n1281) );
  nd2bd1_hd U2033 ( .AN(z_m[1]), .B(n198), .Y(n1280) );
  nd3bd1_hd U2034 ( .AN(z_m[2]), .B(n199), .C(n23), .Y(n1277) );
  scg4d1_hd U2035 ( .A(n1279), .B(z_m[2]), .C(n1278), .D(z_m[1]), .E(n188), 
        .F(n184), .G(n458), .H(product[28]), .Y(n281) );
  ivd1_hd U2036 ( .A(n1281), .Y(n1282) );
  scg4d1_hd U2037 ( .A(n1283), .B(n23), .C(n1282), .D(z_m[1]), .E(z_m[2]), .F(
        n186), .G(n458), .H(product[27]), .Y(n282) );
  nr4d1_hd U2038 ( .A(product[14]), .B(product[12]), .C(product[19]), .D(
        product[17]), .Y(n1287) );
  nr4d1_hd U2039 ( .A(product[15]), .B(product[8]), .C(product[20]), .D(
        product[4]), .Y(n1286) );
  nr4d1_hd U2040 ( .A(product[21]), .B(product[2]), .C(product[13]), .D(
        product[16]), .Y(n1285) );
  nr4d1_hd U2041 ( .A(product[23]), .B(product[5]), .C(product[22]), .D(
        product[18]), .Y(n1284) );
  nd4d1_hd U2042 ( .A(n1287), .B(n1286), .C(n1285), .D(n1284), .Y(n1288) );
  nr4d1_hd U2043 ( .A(product[9]), .B(product[7]), .C(n1289), .D(n1288), .Y(
        n1293) );
  ao22d1_hd U2044 ( .A(round_bit), .B(n1290), .C(sticky), .D(n1292), .Y(n1291)
         );
  oa21d1_hd U2045 ( .A(n1293), .B(n1292), .C(n1291), .Y(n283) );
  ao22d1_hd U2046 ( .A(n456), .B(product[24]), .C(round_bit), .D(n1294), .Y(
        n1295) );
  scg16d1_hd U2047 ( .A(n185), .B(net908), .C(n1295), .Y(n284) );
  ao22d1_hd U2048 ( .A(n456), .B(product[26]), .C(z_m[1]), .D(n183), .Y(n1299)
         );
  ao21d1_hd U2049 ( .A(n95), .B(z_m[0]), .C(n1297), .Y(n1298) );
  oa211d1_hd U2050 ( .A(net908), .B(n194), .C(n1299), .D(n1298), .Y(n285) );
  ao21d1_hd U2051 ( .A(n1276), .B(n1306), .C(n1301), .Y(n1311) );
  ao22d1_hd U2052 ( .A(n457), .B(product[49]), .C(z_m[22]), .D(n100), .Y(n1309) );
  nr3d1_hd U2053 ( .A(n1306), .B(n1305), .C(n1304), .Y(n1416) );
  nd3d1_hd U2054 ( .A(n198), .B(n1416), .C(n1310), .Y(n1308) );
  oa211d1_hd U2055 ( .A(n1311), .B(n1310), .C(n1309), .D(n1308), .Y(n286) );
  ao22d1_hd U2056 ( .A(n481), .B(b[22]), .C(intadd_3_A_17_), .D(n210), .Y(
        n1312) );
  oa21d1_hd U2057 ( .A(n602), .B(n113), .C(n1312), .Y(n287) );
  ao22d1_hd U2058 ( .A(n480), .B(b[20]), .C(intadd_3_B_16_), .D(n212), .Y(
        n1313) );
  ao22d1_hd U2059 ( .A(n480), .B(b[19]), .C(intadd_3_B_15_), .D(n211), .Y(
        n1314) );
  oa21d1_hd U2060 ( .A(n586), .B(n113), .C(n1314), .Y(n289) );
  ao22d1_hd U2061 ( .A(n480), .B(b[18]), .C(b_m[17]), .D(n211), .Y(n1315) );
  ao22d1_hd U2062 ( .A(n480), .B(b[17]), .C(intadd_3_B_13_), .D(n210), .Y(
        n1316) );
  ao22d1_hd U2063 ( .A(n480), .B(b[16]), .C(intadd_3_B_12_), .D(n210), .Y(
        n1317) );
  oa21d1_hd U2064 ( .A(n573), .B(n112), .C(n1317), .Y(n292) );
  ao22d1_hd U2065 ( .A(n479), .B(b[15]), .C(intadd_3_B_11_), .D(n213), .Y(
        n1318) );
  oa21d1_hd U2066 ( .A(n568), .B(n113), .C(n1318), .Y(n293) );
  ao22d1_hd U2067 ( .A(n479), .B(b[14]), .C(intadd_3_B_10_), .D(n213), .Y(
        n1319) );
  ao22d1_hd U2068 ( .A(n479), .B(b[13]), .C(intadd_3_B_9_), .D(n212), .Y(n1320) );
  oa21d1_hd U2069 ( .A(n559), .B(n1335), .C(n1320), .Y(n295) );
  ao22d1_hd U2070 ( .A(n479), .B(b[12]), .C(intadd_3_B_8_), .D(n212), .Y(n1321) );
  ao22d1_hd U2071 ( .A(n479), .B(b[11]), .C(intadd_3_B_7_), .D(n211), .Y(n1322) );
  oa21d1_hd U2072 ( .A(n550), .B(n112), .C(n1322), .Y(n297) );
  ao22d1_hd U2073 ( .A(n479), .B(b[10]), .C(intadd_3_B_6_), .D(n210), .Y(n1323) );
  oa21d1_hd U2074 ( .A(n545), .B(n113), .C(n1323), .Y(n298) );
  ao22d1_hd U2075 ( .A(n478), .B(b[9]), .C(intadd_3_B_5_), .D(n213), .Y(n1324)
         );
  oa21d1_hd U2076 ( .A(n540), .B(n1335), .C(n1324), .Y(n299) );
  ao22d1_hd U2077 ( .A(n478), .B(b[8]), .C(intadd_3_B_4_), .D(n211), .Y(n1325)
         );
  ao22d1_hd U2078 ( .A(n478), .B(b[7]), .C(intadd_3_B_3_), .D(n212), .Y(n1326)
         );
  oa21d1_hd U2079 ( .A(n530), .B(n112), .C(n1326), .Y(n301) );
  ao22d1_hd U2080 ( .A(n478), .B(b[6]), .C(intadd_3_B_2_), .D(n210), .Y(n1327)
         );
  ao22d1_hd U2081 ( .A(n478), .B(b[5]), .C(intadd_3_B_1_), .D(n213), .Y(n1328)
         );
  ao22d1_hd U2082 ( .A(n486), .B(b[4]), .C(intadd_3_B_0_), .D(n211), .Y(n1329)
         );
  oa21d1_hd U2083 ( .A(n518), .B(n113), .C(n1329), .Y(n304) );
  ao22d1_hd U2084 ( .A(n486), .B(b[3]), .C(n503), .D(n210), .Y(n1330) );
  oa21d1_hd U2085 ( .A(n514), .B(n1335), .C(n1330), .Y(n305) );
  ao22d1_hd U2086 ( .A(n486), .B(b[2]), .C(b_m[1]), .D(n213), .Y(n1331) );
  oa21d1_hd U2087 ( .A(n508), .B(n112), .C(n1331), .Y(n306) );
  ao22d1_hd U2088 ( .A(n1332), .B(b[1]), .C(b_m[0]), .D(n212), .Y(n1333) );
  oa21d1_hd U2089 ( .A(n93), .B(n113), .C(n1333), .Y(n307) );
  ao22d1_hd U2090 ( .A(n486), .B(b[21]), .C(intadd_3_B_17_), .D(n211), .Y(
        n1337) );
  oa21d1_hd U2091 ( .A(n596), .B(n1335), .C(n1337), .Y(n309) );
  ivd1_hd U2092 ( .A(n1338), .Y(n1407) );
  ao22d1_hd U2093 ( .A(n106), .B(n598), .C(n108), .D(n379), .Y(n1339) );
  oa21d1_hd U2094 ( .A(n1340), .B(n1407), .C(n1339), .Y(n310) );
  oa211d1_hd U2095 ( .A(n1349), .B(n1342), .C(n1347), .D(n1341), .Y(n1344) );
  ao211d1_hd U2096 ( .A(a_e[8]), .B(n102), .C(DP_OP_113J2_124_6892_n3), .D(
        n1343), .Y(n1353) );
  ao22d1_hd U2097 ( .A(a_e[8]), .B(n1344), .C(n1353), .D(n78), .Y(n1345) );
  ao22d1_hd U2098 ( .A(a_e[1]), .B(n79), .C(C81_DATA2_1), .D(n77), .Y(n1346)
         );
  nr2d1_hd U2099 ( .A(n1349), .B(n1355), .Y(n1352) );
  oa211d1_hd U2100 ( .A(n1353), .B(n1352), .C(n77), .D(n1350), .Y(n1354) );
  oa211d1_hd U2101 ( .A(n1347), .B(n1355), .C(n138), .D(n1354), .Y(n319) );
  ivd1_hd U2102 ( .A(n1356), .Y(n1358) );
  nr2d1_hd U2103 ( .A(DP_OP_116J2_127_7148_n3), .B(n1358), .Y(n1357) );
  oa21d1_hd U2104 ( .A(n1357), .B(n1409), .C(n1362), .Y(n1359) );
  ao211d1_hd U2105 ( .A(n103), .B(b_e[8]), .C(DP_OP_116J2_127_7148_n3), .D(
        n1358), .Y(n1413) );
  ao22d1_hd U2106 ( .A(b_e[8]), .B(n1359), .C(n1413), .D(n82), .Y(n1360) );
  ao22d1_hd U2107 ( .A(b_e[1]), .B(n83), .C(C82_DATA2_1), .D(n81), .Y(n1361)
         );
  oa22d1_hd U2108 ( .A(n164), .B(n114), .C(n1377), .D(n1404), .Y(n328) );
  ao22d1_hd U2109 ( .A(n1332), .B(a[20]), .C(n120), .D(n203), .Y(n1365) );
  oa21d1_hd U2110 ( .A(n164), .B(n1366), .C(n1365), .Y(n329) );
  ao22d1_hd U2111 ( .A(n477), .B(a[19]), .C(n122), .D(a_m[19]), .Y(n1367) );
  oa21d1_hd U2112 ( .A(n165), .B(n1368), .C(n1367), .Y(n330) );
  oa22d1_hd U2113 ( .A(n163), .B(n460), .C(n1377), .D(n1368), .Y(n331) );
  ao22d1_hd U2114 ( .A(n477), .B(a[17]), .C(n122), .D(n92), .Y(n1370) );
  oa21d1_hd U2115 ( .A(n164), .B(n1371), .C(n1370), .Y(n332) );
  ao22d1_hd U2116 ( .A(n478), .B(a[16]), .C(n123), .D(a_m[16]), .Y(n1372) );
  oa21d1_hd U2117 ( .A(n163), .B(n1373), .C(n1372), .Y(n333) );
  ao22d1_hd U2118 ( .A(n477), .B(a[15]), .C(n122), .D(a_m[15]), .Y(n1374) );
  oa21d1_hd U2119 ( .A(n162), .B(n125), .C(n1374), .Y(n334) );
  ao22d1_hd U2120 ( .A(n477), .B(a[14]), .C(n121), .D(a_m[14]), .Y(n1375) );
  oa21d1_hd U2121 ( .A(n163), .B(n1376), .C(n1375), .Y(n335) );
  oa22d1_hd U2122 ( .A(n162), .B(n1378), .C(n1377), .D(n1376), .Y(n336) );
  ao22d1_hd U2123 ( .A(n477), .B(a[12]), .C(n123), .D(a_m[12]), .Y(n1379) );
  oa21d1_hd U2124 ( .A(n165), .B(n462), .C(n1379), .Y(n337) );
  ao22d1_hd U2125 ( .A(n476), .B(a[11]), .C(n120), .D(n193), .Y(n1381) );
  oa21d1_hd U2126 ( .A(n164), .B(n1382), .C(n1381), .Y(n338) );
  ao22d1_hd U2127 ( .A(n476), .B(a[10]), .C(n121), .D(a_m[10]), .Y(n1383) );
  oa21d1_hd U2128 ( .A(n163), .B(n1384), .C(n1383), .Y(n339) );
  ao22d1_hd U2129 ( .A(n476), .B(a[9]), .C(n123), .D(a_m[9]), .Y(n1385) );
  oa21d1_hd U2130 ( .A(n162), .B(n608), .C(n1385), .Y(n340) );
  ao22d1_hd U2131 ( .A(n476), .B(a[8]), .C(n120), .D(n604), .Y(n1386) );
  oa21d1_hd U2132 ( .A(n165), .B(n1387), .C(n1386), .Y(n341) );
  ao22d1_hd U2133 ( .A(n476), .B(a[7]), .C(n122), .D(a_m[7]), .Y(n1388) );
  oa21d1_hd U2134 ( .A(n164), .B(n1389), .C(n1388), .Y(n342) );
  ao22d1_hd U2135 ( .A(n476), .B(a[6]), .C(n123), .D(a_m[6]), .Y(n1390) );
  oa21d1_hd U2136 ( .A(n163), .B(n85), .C(n1390), .Y(n343) );
  ao22d1_hd U2137 ( .A(n1332), .B(a[5]), .C(n120), .D(a_m[5]), .Y(n1392) );
  oa21d1_hd U2138 ( .A(n162), .B(n1393), .C(n1392), .Y(n344) );
  ao22d1_hd U2139 ( .A(n485), .B(a[4]), .C(n121), .D(a_m[4]), .Y(n1394) );
  oa21d1_hd U2140 ( .A(n165), .B(n1395), .C(n1394), .Y(n345) );
  ao22d1_hd U2141 ( .A(n477), .B(a[3]), .C(n120), .D(a_m[3]), .Y(n1396) );
  oa21d1_hd U2142 ( .A(n164), .B(n471), .C(n1396), .Y(n346) );
  ao22d1_hd U2143 ( .A(n484), .B(a[2]), .C(n121), .D(n196), .Y(n1398) );
  oa21d1_hd U2144 ( .A(n163), .B(n1399), .C(n1398), .Y(n347) );
  ao22d1_hd U2145 ( .A(n485), .B(a[1]), .C(n121), .D(a_m[1]), .Y(n1400) );
  oa21d1_hd U2146 ( .A(n162), .B(n1401), .C(n1400), .Y(n348) );
  ao22d1_hd U2147 ( .A(n485), .B(a[22]), .C(n122), .D(a_m[22]), .Y(n1403) );
  oa21d1_hd U2148 ( .A(n165), .B(n1404), .C(n1403), .Y(n354) );
  ao22d1_hd U2149 ( .A(a_m[22]), .B(n102), .C(n618), .D(n380), .Y(n1406) );
  oa21d1_hd U2150 ( .A(n1408), .B(n1407), .C(n1406), .Y(n355) );
  nr2d1_hd U2151 ( .A(n1415), .B(n1409), .Y(n1412) );
  oa211d1_hd U2152 ( .A(n1413), .B(n1412), .C(n81), .D(n1410), .Y(n1414) );
  oa211d1_hd U2153 ( .A(n1362), .B(n1415), .C(n148), .D(n1414), .Y(n356) );
  ivd1_hd U2154 ( .A(state[3]), .Y(n1614) );
  ivd1_hd U2155 ( .A(n3277), .Y(n1613) );
  ivd1_hd U2156 ( .A(o_AB_ACK), .Y(n1544) );
endmodule


module float_multiplier_0 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, 
        i_Z_ACK, i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N34, a_s, b_s, N35, round_bit, sticky, z_s, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201,
         N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212,
         N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223,
         N467, N468, N469, N470, N471, N472, N473, N474, N475, C82_DATA2_1,
         C82_DATA2_2, C82_DATA2_3, C82_DATA2_4, C82_DATA2_5, C82_DATA2_6,
         C81_DATA2_1, C81_DATA2_2, C81_DATA2_3, C81_DATA2_4, C81_DATA2_5,
         C81_DATA2_6, net908, n10, n14, n36, n104, n105, n138, n141, n146,
         n148, n151, n155, n156, n157, n158, n160, n161, n171, n172, n173,
         n174, n177, n179, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, DP_OP_116J2_127_7148_n3, DP_OP_116J2_127_7148_n4,
         DP_OP_116J2_127_7148_n5, DP_OP_116J2_127_7148_n6,
         DP_OP_116J2_127_7148_n7, DP_OP_116J2_127_7148_n8,
         DP_OP_113J2_124_6892_n3, DP_OP_113J2_124_6892_n4,
         DP_OP_113J2_124_6892_n5, DP_OP_113J2_124_6892_n6,
         DP_OP_113J2_124_6892_n7, DP_OP_113J2_124_6892_n8, C1_Z_6, C1_Z_5,
         C1_Z_4, C1_Z_3, C1_Z_2, C1_Z_1, DP_OP_125J2_130_6300_n42,
         DP_OP_125J2_130_6300_n41, DP_OP_125J2_130_6300_n40,
         DP_OP_125J2_130_6300_n39, DP_OP_125J2_130_6300_n38,
         DP_OP_125J2_130_6300_n37, DP_OP_125J2_130_6300_n36,
         DP_OP_125J2_130_6300_n35, DP_OP_125J2_130_6300_n34,
         DP_OP_125J2_130_6300_n32, DP_OP_125J2_130_6300_n31,
         DP_OP_125J2_130_6300_n30, DP_OP_125J2_130_6300_n29,
         DP_OP_125J2_130_6300_n28, DP_OP_125J2_130_6300_n27,
         DP_OP_125J2_130_6300_n26, DP_OP_125J2_130_6300_n25,
         DP_OP_125J2_130_6300_n20, DP_OP_125J2_130_6300_n19,
         DP_OP_125J2_130_6300_n18, DP_OP_125J2_130_6300_n17,
         DP_OP_125J2_130_6300_n16, DP_OP_125J2_130_6300_n15,
         DP_OP_125J2_130_6300_n14, DP_OP_125J2_130_6300_n13,
         DP_OP_125J2_130_6300_n12, DP_OP_125J2_130_6300_n9,
         DP_OP_125J2_130_6300_n8, DP_OP_125J2_130_6300_n7,
         DP_OP_125J2_130_6300_n6, DP_OP_125J2_130_6300_n5,
         DP_OP_125J2_130_6300_n4, DP_OP_125J2_130_6300_n3,
         DP_OP_125J2_130_6300_n2, n381, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1332, intadd_24_A_16_, intadd_24_A_15_,
         intadd_24_A_13_, intadd_24_A_12_, intadd_24_A_11_, intadd_24_A_10_,
         intadd_24_A_9_, intadd_24_A_8_, intadd_24_A_7_, intadd_24_A_6_,
         intadd_24_A_5_, intadd_24_A_4_, intadd_24_A_3_, intadd_24_A_2_,
         intadd_24_A_1_, intadd_24_A_0_, intadd_24_B_16_, intadd_24_B_15_,
         intadd_24_B_14_, intadd_24_B_13_, intadd_24_B_12_, intadd_24_B_11_,
         intadd_24_B_10_, intadd_24_B_9_, intadd_24_B_8_, intadd_24_B_7_,
         intadd_24_B_6_, intadd_24_B_5_, intadd_24_B_4_, intadd_24_B_3_,
         intadd_24_B_2_, intadd_24_B_1_, intadd_24_B_0_, intadd_24_CI,
         intadd_24_SUM_16_, intadd_24_SUM_15_, intadd_24_SUM_14_,
         intadd_24_SUM_13_, intadd_24_SUM_12_, intadd_24_SUM_11_,
         intadd_24_SUM_10_, intadd_24_SUM_9_, intadd_24_SUM_8_,
         intadd_24_SUM_7_, intadd_24_SUM_6_, intadd_24_SUM_5_,
         intadd_24_SUM_4_, intadd_24_SUM_3_, intadd_24_SUM_2_,
         intadd_24_SUM_1_, intadd_24_SUM_0_, intadd_24_n17, intadd_24_n16,
         intadd_24_n15, intadd_24_n14, intadd_24_n13, intadd_24_n12,
         intadd_24_n11, intadd_24_n10, intadd_24_n9, intadd_24_n8,
         intadd_24_n7, intadd_24_n6, intadd_24_n5, intadd_24_n4, intadd_24_n3,
         intadd_24_n2, intadd_24_n1, intadd_25_A_11_, intadd_25_A_10_,
         intadd_25_A_9_, intadd_25_A_8_, intadd_25_A_7_, intadd_25_A_6_,
         intadd_25_A_5_, intadd_25_A_4_, intadd_25_A_3_, intadd_25_A_2_,
         intadd_25_A_1_, intadd_25_A_0_, intadd_25_B_11_, intadd_25_B_10_,
         intadd_25_B_9_, intadd_25_B_8_, intadd_25_B_7_, intadd_25_B_6_,
         intadd_25_B_5_, intadd_25_B_4_, intadd_25_B_3_, intadd_25_B_2_,
         intadd_25_B_1_, intadd_25_B_0_, intadd_25_CI, intadd_25_SUM_11_,
         intadd_25_SUM_10_, intadd_25_SUM_9_, intadd_25_SUM_8_,
         intadd_25_SUM_7_, intadd_25_SUM_6_, intadd_25_SUM_5_,
         intadd_25_SUM_4_, intadd_25_SUM_3_, intadd_25_SUM_2_,
         intadd_25_SUM_1_, intadd_25_SUM_0_, intadd_25_n12, intadd_25_n11,
         intadd_25_n10, intadd_25_n9, intadd_25_n8, intadd_25_n7, intadd_25_n6,
         intadd_25_n5, intadd_25_n4, intadd_25_n3, intadd_25_n2, intadd_25_n1,
         intadd_26_A_10_, intadd_26_A_8_, intadd_26_A_7_, intadd_26_A_6_,
         intadd_26_A_5_, intadd_26_A_3_, intadd_26_A_2_, intadd_26_A_1_,
         intadd_26_A_0_, intadd_26_B_9_, intadd_26_B_4_, intadd_26_B_2_,
         intadd_26_B_1_, intadd_26_B_0_, intadd_26_CI, intadd_26_n11,
         intadd_26_n10, intadd_26_n9, intadd_26_n8, intadd_26_n7, intadd_26_n6,
         intadd_26_n5, intadd_26_n4, intadd_26_n3, intadd_26_n2, intadd_26_n1,
         intadd_27_A_10_, intadd_27_A_9_, intadd_27_A_8_, intadd_27_A_7_,
         intadd_27_A_6_, intadd_27_A_5_, intadd_27_A_4_, intadd_27_A_3_,
         intadd_27_A_2_, intadd_27_A_1_, intadd_27_A_0_, intadd_27_B_10_,
         intadd_27_B_9_, intadd_27_B_8_, intadd_27_B_7_, intadd_27_B_6_,
         intadd_27_B_5_, intadd_27_B_4_, intadd_27_B_3_, intadd_27_B_2_,
         intadd_27_B_1_, intadd_27_B_0_, intadd_27_CI, intadd_27_SUM_10_,
         intadd_27_SUM_9_, intadd_27_SUM_8_, intadd_27_SUM_7_,
         intadd_27_SUM_6_, intadd_27_SUM_5_, intadd_27_SUM_4_,
         intadd_27_SUM_3_, intadd_27_SUM_2_, intadd_27_SUM_1_,
         intadd_27_SUM_0_, intadd_27_n11, intadd_27_n10, intadd_27_n9,
         intadd_27_n8, intadd_27_n7, intadd_27_n6, intadd_27_n5, intadd_27_n4,
         intadd_27_n3, intadd_27_n2, intadd_27_n1, intadd_28_A_8_,
         intadd_28_A_7_, intadd_28_A_6_, intadd_28_A_5_, intadd_28_A_3_,
         intadd_28_A_2_, intadd_28_A_1_, intadd_28_B_8_, intadd_28_B_7_,
         intadd_28_B_6_, intadd_28_B_5_, intadd_28_B_4_, intadd_28_B_3_,
         intadd_28_B_2_, intadd_28_B_1_, intadd_28_B_0_, intadd_28_CI,
         intadd_28_SUM_8_, intadd_28_SUM_7_, intadd_28_SUM_6_,
         intadd_28_SUM_5_, intadd_28_SUM_4_, intadd_28_SUM_0_, intadd_28_n9,
         intadd_28_n8, intadd_28_n7, intadd_28_n6, intadd_28_n5, intadd_28_n4,
         intadd_28_n3, intadd_28_n2, intadd_28_n1, intadd_29_A_7_,
         intadd_29_A_6_, intadd_29_A_5_, intadd_29_A_4_, intadd_29_A_3_,
         intadd_29_A_2_, intadd_29_A_1_, intadd_29_B_7_, intadd_29_B_6_,
         intadd_29_B_5_, intadd_29_B_4_, intadd_29_B_3_, intadd_29_B_2_,
         intadd_29_B_1_, intadd_29_CI, intadd_29_SUM_7_, intadd_29_SUM_6_,
         intadd_29_SUM_5_, intadd_29_SUM_4_, intadd_29_SUM_3_,
         intadd_29_SUM_2_, intadd_29_SUM_1_, intadd_29_SUM_0_, intadd_29_n8,
         intadd_29_n7, intadd_29_n6, intadd_29_n5, intadd_29_n4, intadd_29_n3,
         intadd_29_n2, intadd_29_n1, intadd_30_A_5_, intadd_30_A_4_,
         intadd_30_A_3_, intadd_30_A_2_, intadd_30_A_1_, intadd_30_A_0_,
         intadd_30_B_5_, intadd_30_B_4_, intadd_30_B_3_, intadd_30_B_2_,
         intadd_30_B_1_, intadd_30_B_0_, intadd_30_CI, intadd_30_SUM_5_,
         intadd_30_SUM_4_, intadd_30_SUM_3_, intadd_30_SUM_2_,
         intadd_30_SUM_1_, intadd_30_SUM_0_, intadd_30_n6, intadd_30_n5,
         intadd_30_n4, intadd_30_n3, intadd_30_n2, intadd_30_n1,
         intadd_31_A_4_, intadd_31_A_3_, intadd_31_A_2_, intadd_31_A_1_,
         intadd_31_A_0_, intadd_31_B_4_, intadd_31_B_3_, intadd_31_B_2_,
         intadd_31_B_1_, intadd_31_B_0_, intadd_31_CI, intadd_31_SUM_4_,
         intadd_31_SUM_3_, intadd_31_SUM_2_, intadd_31_SUM_1_,
         intadd_31_SUM_0_, intadd_31_n5, intadd_31_n4, intadd_31_n3,
         intadd_31_n2, intadd_31_n1, intadd_32_A_2_, intadd_32_A_1_,
         intadd_32_B_2_, intadd_32_B_1_, intadd_32_B_0_, intadd_32_CI,
         intadd_32_n3, intadd_32_n2, intadd_32_n1, intadd_33_A_2_,
         intadd_33_A_1_, intadd_33_A_0_, intadd_33_B_2_, intadd_33_B_1_,
         intadd_33_B_0_, intadd_33_CI, intadd_33_SUM_2_, intadd_33_SUM_1_,
         intadd_33_SUM_0_, intadd_33_n3, intadd_33_n2, intadd_33_n1,
         intadd_34_A_2_, intadd_34_A_1_, intadd_34_A_0_, intadd_34_B_2_,
         intadd_34_B_1_, intadd_34_B_0_, intadd_34_CI, intadd_34_SUM_2_,
         intadd_34_SUM_1_, intadd_34_SUM_0_, intadd_34_n3, intadd_34_n2,
         intadd_34_n1, intadd_35_A_0_, intadd_35_B_2_, intadd_35_B_1_,
         intadd_35_B_0_, intadd_35_SUM_2_, intadd_35_SUM_1_, intadd_35_SUM_0_,
         intadd_35_n3, intadd_35_n2, intadd_35_n1, intadd_36_B_2_,
         intadd_36_B_1_, intadd_36_B_0_, intadd_36_CI, intadd_36_SUM_2_,
         intadd_36_SUM_1_, intadd_36_SUM_0_, intadd_36_n3, intadd_36_n2,
         intadd_36_n1, intadd_37_A_2_, intadd_37_A_1_, intadd_37_A_0_,
         intadd_37_B_2_, intadd_37_B_1_, intadd_37_B_0_, intadd_37_CI,
         intadd_37_SUM_2_, intadd_37_SUM_1_, intadd_37_SUM_0_, intadd_37_n3,
         intadd_37_n2, intadd_37_n1, intadd_38_B_2_, intadd_38_B_1_,
         intadd_38_B_0_, intadd_38_CI, intadd_38_SUM_2_, intadd_38_SUM_1_,
         intadd_38_SUM_0_, intadd_38_n3, intadd_38_n2, intadd_38_n1,
         intadd_39_A_1_, intadd_39_A_0_, intadd_39_B_2_, intadd_39_CI,
         intadd_39_SUM_2_, intadd_39_n3, intadd_39_n2, intadd_39_n1,
         intadd_20_A_36_, intadd_20_A_35_, intadd_20_A_34_, intadd_20_A_33_,
         intadd_20_A_31_, intadd_20_A_30_, intadd_20_A_29_, intadd_20_A_27_,
         intadd_20_A_26_, intadd_20_A_24_, intadd_20_A_23_, intadd_20_A_21_,
         intadd_20_A_20_, intadd_20_A_19_, intadd_20_A_18_, intadd_20_A_17_,
         intadd_20_A_16_, intadd_20_A_15_, intadd_20_A_14_, intadd_20_A_13_,
         intadd_20_A_12_, intadd_20_A_11_, intadd_20_A_10_, intadd_20_A_9_,
         intadd_20_A_8_, intadd_20_A_7_, intadd_20_A_6_, intadd_20_A_5_,
         intadd_20_A_4_, intadd_20_A_3_, intadd_20_A_2_, intadd_20_A_1_,
         intadd_20_A_0_, intadd_20_B_36_, intadd_20_B_35_, intadd_20_B_34_,
         intadd_20_B_32_, intadd_20_B_31_, intadd_20_B_30_, intadd_20_B_28_,
         intadd_20_B_27_, intadd_20_B_25_, intadd_20_B_24_, intadd_20_B_22_,
         intadd_20_B_21_, intadd_20_B_20_, intadd_20_B_19_, intadd_20_B_18_,
         intadd_20_B_17_, intadd_20_B_16_, intadd_20_B_15_, intadd_20_B_14_,
         intadd_20_B_13_, intadd_20_B_12_, intadd_20_B_11_, intadd_20_B_10_,
         intadd_20_B_9_, intadd_20_B_8_, intadd_20_B_7_, intadd_20_B_6_,
         intadd_20_B_5_, intadd_20_B_4_, intadd_20_B_3_, intadd_20_B_2_,
         intadd_20_B_1_, intadd_20_B_0_, intadd_20_CI, intadd_20_SUM_16_,
         intadd_20_SUM_15_, intadd_20_SUM_14_, intadd_20_SUM_13_,
         intadd_20_SUM_12_, intadd_20_SUM_11_, intadd_20_SUM_10_,
         intadd_20_SUM_9_, intadd_20_SUM_8_, intadd_20_SUM_7_,
         intadd_20_SUM_6_, intadd_20_SUM_5_, intadd_20_SUM_4_,
         intadd_20_SUM_3_, intadd_20_SUM_2_, intadd_20_SUM_1_,
         intadd_20_SUM_0_, intadd_20_n37, intadd_20_n36, intadd_20_n35,
         intadd_20_n34, intadd_20_n33, intadd_20_n32, intadd_20_n31,
         intadd_20_n30, intadd_20_n29, intadd_20_n28, intadd_20_n27,
         intadd_20_n26, intadd_20_n25, intadd_20_n24, intadd_20_n23,
         intadd_20_n22, intadd_20_n21, intadd_20_n20, intadd_20_n19,
         intadd_20_n18, intadd_20_n17, intadd_20_n16, intadd_20_n15,
         intadd_20_n14, intadd_20_n13, intadd_20_n12, intadd_20_n11,
         intadd_20_n10, intadd_20_n9, intadd_20_n8, intadd_20_n7, intadd_20_n6,
         intadd_20_n5, intadd_20_n4, intadd_20_n3, intadd_20_n2, intadd_20_n1,
         intadd_21_A_21_, intadd_21_A_20_, intadd_21_A_19_, intadd_21_A_18_,
         intadd_21_A_17_, intadd_21_A_16_, intadd_21_A_15_, intadd_21_A_14_,
         intadd_21_A_13_, intadd_21_A_12_, intadd_21_A_11_, intadd_21_A_10_,
         intadd_21_A_9_, intadd_21_A_8_, intadd_21_A_7_, intadd_21_A_6_,
         intadd_21_A_5_, intadd_21_A_4_, intadd_21_A_3_, intadd_21_A_2_,
         intadd_21_A_1_, intadd_21_A_0_, intadd_21_B_22_, intadd_21_B_21_,
         intadd_21_B_20_, intadd_21_B_19_, intadd_21_B_18_, intadd_21_B_17_,
         intadd_21_B_16_, intadd_21_B_15_, intadd_21_B_14_, intadd_21_B_13_,
         intadd_21_B_12_, intadd_21_B_11_, intadd_21_B_10_, intadd_21_B_9_,
         intadd_21_B_8_, intadd_21_B_7_, intadd_21_B_6_, intadd_21_B_5_,
         intadd_21_B_4_, intadd_21_B_3_, intadd_21_B_2_, intadd_21_B_1_,
         intadd_21_B_0_, intadd_21_CI, intadd_21_SUM_22_, intadd_21_SUM_21_,
         intadd_21_SUM_20_, intadd_21_SUM_19_, intadd_21_SUM_18_,
         intadd_21_SUM_17_, intadd_21_SUM_16_, intadd_21_SUM_15_,
         intadd_21_SUM_14_, intadd_21_SUM_13_, intadd_21_SUM_12_,
         intadd_21_SUM_11_, intadd_21_SUM_10_, intadd_21_SUM_9_,
         intadd_21_SUM_8_, intadd_21_SUM_7_, intadd_21_SUM_6_,
         intadd_21_SUM_5_, intadd_21_SUM_4_, intadd_21_SUM_3_,
         intadd_21_SUM_2_, intadd_21_SUM_1_, intadd_21_SUM_0_, intadd_21_n23,
         intadd_21_n22, intadd_21_n21, intadd_21_n20, intadd_21_n19,
         intadd_21_n18, intadd_21_n17, intadd_21_n16, intadd_21_n15,
         intadd_21_n14, intadd_21_n13, intadd_21_n12, intadd_21_n11,
         intadd_21_n10, intadd_21_n9, intadd_21_n8, intadd_21_n7, intadd_21_n6,
         intadd_21_n5, intadd_21_n4, intadd_21_n3, intadd_21_n2, intadd_21_n1,
         intadd_22_A_18_, intadd_22_A_17_, intadd_22_A_16_, intadd_22_A_15_,
         intadd_22_A_14_, intadd_22_A_13_, intadd_22_A_12_, intadd_22_A_11_,
         intadd_22_A_10_, intadd_22_A_9_, intadd_22_A_8_, intadd_22_A_7_,
         intadd_22_A_6_, intadd_22_A_5_, intadd_22_A_4_, intadd_22_A_3_,
         intadd_22_A_2_, intadd_22_A_1_, intadd_22_A_0_, intadd_22_B_18_,
         intadd_22_B_17_, intadd_22_B_16_, intadd_22_B_15_, intadd_22_B_14_,
         intadd_22_B_13_, intadd_22_B_12_, intadd_22_B_11_, intadd_22_B_10_,
         intadd_22_B_9_, intadd_22_B_8_, intadd_22_B_7_, intadd_22_B_6_,
         intadd_22_B_5_, intadd_22_B_4_, intadd_22_B_3_, intadd_22_B_2_,
         intadd_22_B_1_, intadd_22_B_0_, intadd_22_CI, intadd_22_n19,
         intadd_22_n18, intadd_22_n17, intadd_22_n16, intadd_22_n15,
         intadd_22_n14, intadd_22_n13, intadd_22_n12, intadd_22_n11,
         intadd_22_n10, intadd_22_n9, intadd_22_n8, intadd_22_n7, intadd_22_n6,
         intadd_22_n5, intadd_22_n4, intadd_22_n3, intadd_22_n2, intadd_22_n1,
         intadd_23_A_17_, intadd_23_B_17_, intadd_23_B_16_, intadd_23_B_15_,
         intadd_23_B_14_, intadd_23_B_13_, intadd_23_B_12_, intadd_23_B_11_,
         intadd_23_B_10_, intadd_23_B_9_, intadd_23_B_8_, intadd_23_B_7_,
         intadd_23_B_6_, intadd_23_B_5_, intadd_23_B_4_, intadd_23_B_3_,
         intadd_23_B_2_, intadd_23_B_1_, intadd_23_B_0_, intadd_23_CI,
         intadd_23_SUM_17_, intadd_23_SUM_16_, intadd_23_SUM_15_,
         intadd_23_SUM_14_, intadd_23_SUM_13_, intadd_23_SUM_12_,
         intadd_23_SUM_11_, intadd_23_SUM_10_, intadd_23_SUM_9_,
         intadd_23_SUM_8_, intadd_23_SUM_7_, intadd_23_SUM_6_,
         intadd_23_SUM_5_, intadd_23_SUM_4_, intadd_23_SUM_3_,
         intadd_23_SUM_2_, intadd_23_SUM_1_, intadd_23_SUM_0_, intadd_23_n18,
         intadd_23_n17, intadd_23_n16, intadd_23_n15, intadd_23_n14,
         intadd_23_n13, intadd_23_n12, intadd_23_n11, intadd_23_n10,
         intadd_23_n9, intadd_23_n8, intadd_23_n7, intadd_23_n6, intadd_23_n5,
         intadd_23_n4, intadd_23_n3, intadd_23_n2, intadd_23_n1, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n11, n12, n13, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n139, n140,
         n142, n143, n144, n145, n147, n149, n150, n152, n153, n154, n159,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n175, n176,
         n178, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [23:0] a_m;
  wire   [9:0] b_e;
  wire   [23:0] b_m;
  wire   [49:2] product;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ao211d1_hd U246 ( .A(n1437), .B(n155), .C(i_RST), .D(n500), .Y(n350) );
  oa22d1_hd U247 ( .A(n156), .B(n157), .C(n1432), .D(n158), .Y(n351) );
  oa22d1_hd U249 ( .A(n160), .B(n157), .C(n78), .D(n158), .Y(n352) );
  oa22d1_hd U250 ( .A(n161), .B(n157), .C(n1431), .D(n158), .Y(n353) );
  oa22d1_hd U267 ( .A(n171), .B(n157), .C(n1435), .D(n158), .Y(n357) );
  nd4d1_hd U269 ( .A(n160), .B(n172), .C(n173), .D(n174), .Y(n158) );
  ao211d1_hd U270 ( .A(n1427), .B(n36), .C(i_RST), .D(n500), .Y(n174) );
  ao211d1_hd U281 ( .A(n476), .B(n177), .C(i_RST), .D(n179), .Y(n358) );
  ivd1_hd U364 ( .A(i_RST), .Y(N34) );
  fad1_hd DP_OP_116J2_127_7148_U6 ( .A(n116), .B(n1213), .CI(
        DP_OP_116J2_127_7148_n4), .CO(DP_OP_116J2_127_7148_n3), .S(C82_DATA2_6) );
  fad1_hd DP_OP_116J2_127_7148_U7 ( .A(n117), .B(n1212), .CI(
        DP_OP_116J2_127_7148_n5), .CO(DP_OP_116J2_127_7148_n4), .S(C82_DATA2_5) );
  fad1_hd DP_OP_116J2_127_7148_U8 ( .A(n118), .B(n1211), .CI(
        DP_OP_116J2_127_7148_n6), .CO(DP_OP_116J2_127_7148_n5), .S(C82_DATA2_4) );
  fad1_hd DP_OP_116J2_127_7148_U9 ( .A(n116), .B(n1210), .CI(
        DP_OP_116J2_127_7148_n7), .CO(DP_OP_116J2_127_7148_n6), .S(C82_DATA2_3) );
  fad1_hd DP_OP_116J2_127_7148_U10 ( .A(n116), .B(n1209), .CI(
        DP_OP_116J2_127_7148_n8), .CO(DP_OP_116J2_127_7148_n7), .S(C82_DATA2_2) );
  fad1_hd DP_OP_116J2_127_7148_U11 ( .A(n117), .B(n1208), .CI(n1207), .CO(
        DP_OP_116J2_127_7148_n8), .S(C82_DATA2_1) );
  fad1_hd DP_OP_113J2_124_6892_U6 ( .A(n117), .B(C1_Z_6), .CI(
        DP_OP_113J2_124_6892_n4), .CO(DP_OP_113J2_124_6892_n3), .S(C81_DATA2_6) );
  fad1_hd DP_OP_113J2_124_6892_U7 ( .A(n118), .B(C1_Z_5), .CI(
        DP_OP_113J2_124_6892_n5), .CO(DP_OP_113J2_124_6892_n4), .S(C81_DATA2_5) );
  fad1_hd DP_OP_113J2_124_6892_U8 ( .A(n116), .B(C1_Z_4), .CI(
        DP_OP_113J2_124_6892_n6), .CO(DP_OP_113J2_124_6892_n5), .S(C81_DATA2_4) );
  fad1_hd DP_OP_113J2_124_6892_U9 ( .A(n117), .B(C1_Z_3), .CI(
        DP_OP_113J2_124_6892_n7), .CO(DP_OP_113J2_124_6892_n6), .S(C81_DATA2_3) );
  fad1_hd DP_OP_113J2_124_6892_U10 ( .A(n117), .B(C1_Z_2), .CI(
        DP_OP_113J2_124_6892_n8), .CO(DP_OP_113J2_124_6892_n7), .S(C81_DATA2_2) );
  fad1_hd DP_OP_113J2_124_6892_U11 ( .A(n118), .B(C1_Z_1), .CI(n1206), .CO(
        DP_OP_113J2_124_6892_n8), .S(C81_DATA2_1) );
  had1_hd DP_OP_125J2_130_6300_U32 ( .A(b_e[0]), .B(a_e[0]), .CO(
        DP_OP_125J2_130_6300_n20), .S(DP_OP_125J2_130_6300_n34) );
  fad1_hd DP_OP_125J2_130_6300_U31 ( .A(a_e[1]), .B(b_e[1]), .CI(
        DP_OP_125J2_130_6300_n20), .CO(DP_OP_125J2_130_6300_n19), .S(
        DP_OP_125J2_130_6300_n35) );
  fad1_hd DP_OP_125J2_130_6300_U30 ( .A(a_e[2]), .B(b_e[2]), .CI(
        DP_OP_125J2_130_6300_n19), .CO(DP_OP_125J2_130_6300_n18), .S(
        DP_OP_125J2_130_6300_n36) );
  fad1_hd DP_OP_125J2_130_6300_U29 ( .A(a_e[3]), .B(b_e[3]), .CI(
        DP_OP_125J2_130_6300_n18), .CO(DP_OP_125J2_130_6300_n17), .S(
        DP_OP_125J2_130_6300_n37) );
  fad1_hd DP_OP_125J2_130_6300_U28 ( .A(a_e[4]), .B(b_e[4]), .CI(
        DP_OP_125J2_130_6300_n17), .CO(DP_OP_125J2_130_6300_n16), .S(
        DP_OP_125J2_130_6300_n38) );
  fad1_hd DP_OP_125J2_130_6300_U27 ( .A(a_e[5]), .B(b_e[5]), .CI(
        DP_OP_125J2_130_6300_n16), .CO(DP_OP_125J2_130_6300_n15), .S(
        DP_OP_125J2_130_6300_n39) );
  fad1_hd DP_OP_125J2_130_6300_U26 ( .A(a_e[6]), .B(b_e[6]), .CI(
        DP_OP_125J2_130_6300_n15), .CO(DP_OP_125J2_130_6300_n14), .S(
        DP_OP_125J2_130_6300_n40) );
  fad1_hd DP_OP_125J2_130_6300_U25 ( .A(a_e[7]), .B(b_e[7]), .CI(
        DP_OP_125J2_130_6300_n14), .CO(DP_OP_125J2_130_6300_n13), .S(
        DP_OP_125J2_130_6300_n41) );
  fad1_hd DP_OP_125J2_130_6300_U24 ( .A(a_e[8]), .B(b_e[8]), .CI(
        DP_OP_125J2_130_6300_n13), .CO(DP_OP_125J2_130_6300_n12), .S(
        DP_OP_125J2_130_6300_n42) );
  fad1_hd DP_OP_125J2_130_6300_U10 ( .A(n1436), .B(n378), .CI(
        DP_OP_125J2_130_6300_n25), .CO(DP_OP_125J2_130_6300_n9), .S(N467) );
  fad1_hd DP_OP_125J2_130_6300_U9 ( .A(DP_OP_125J2_130_6300_n26), .B(n379), 
        .CI(DP_OP_125J2_130_6300_n9), .CO(DP_OP_125J2_130_6300_n8), .S(N468)
         );
  fad1_hd DP_OP_125J2_130_6300_U8 ( .A(DP_OP_125J2_130_6300_n27), .B(n378), 
        .CI(DP_OP_125J2_130_6300_n8), .CO(DP_OP_125J2_130_6300_n7), .S(N469)
         );
  fad1_hd DP_OP_125J2_130_6300_U7 ( .A(DP_OP_125J2_130_6300_n28), .B(n379), 
        .CI(DP_OP_125J2_130_6300_n7), .CO(DP_OP_125J2_130_6300_n6), .S(N470)
         );
  fad1_hd DP_OP_125J2_130_6300_U6 ( .A(DP_OP_125J2_130_6300_n29), .B(n378), 
        .CI(DP_OP_125J2_130_6300_n6), .CO(DP_OP_125J2_130_6300_n5), .S(N471)
         );
  fad1_hd DP_OP_125J2_130_6300_U5 ( .A(DP_OP_125J2_130_6300_n30), .B(n379), 
        .CI(DP_OP_125J2_130_6300_n5), .CO(DP_OP_125J2_130_6300_n4), .S(N472)
         );
  fad1_hd DP_OP_125J2_130_6300_U4 ( .A(DP_OP_125J2_130_6300_n31), .B(n378), 
        .CI(DP_OP_125J2_130_6300_n4), .CO(DP_OP_125J2_130_6300_n3), .S(N473)
         );
  fad1_hd DP_OP_125J2_130_6300_U3 ( .A(DP_OP_125J2_130_6300_n32), .B(n379), 
        .CI(DP_OP_125J2_130_6300_n3), .CO(DP_OP_125J2_130_6300_n2), .S(N474)
         );
  fds2d1_hd a_e_reg_7_ ( .CRN(n141), .D(n138), .CK(i_CLK), .Q(n10), .QN(a_e[7]) );
  fds2d1_hd b_e_reg_7_ ( .CRN(n151), .D(n148), .CK(i_CLK), .Q(n14), .QN(b_e[7]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n319), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n356), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n309), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n306), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n290), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n291), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n292), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n295), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n296), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n299), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n305), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n294), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n289), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n297), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n298), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n302), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n301), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n287), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n304), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n293), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n303), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n300), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n288), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n326), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n317), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n327), .CK(i_CLK), .Q(b_e[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n318), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n325), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n316), .CK(i_CLK), .Q(a_e[2]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n315), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n324), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n323), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n314), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n282), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n322), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n313), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n281), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n285), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n312), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n321), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n262), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n276), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n264), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n280), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n268), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n272), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n261), .CK(i_CLK), .Q(z_m[22]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n270), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n266), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n274), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n278), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n269), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n265), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n277), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n273), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n275), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n267), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n279), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n271), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n263), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n286), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n320), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n311), .CK(i_CLK), .Q(a_e[8]) );
  clknd2d1_hd U552 ( .A(N34), .B(n158), .Y(n157) );
  fad1_hd intadd_24_U18 ( .A(intadd_24_A_0_), .B(intadd_24_B_0_), .CI(
        intadd_24_CI), .CO(intadd_24_n17), .S(intadd_24_SUM_0_) );
  fad1_hd intadd_24_U17 ( .A(intadd_24_A_1_), .B(intadd_24_B_1_), .CI(
        intadd_24_n17), .CO(intadd_24_n16), .S(intadd_24_SUM_1_) );
  fad1_hd intadd_24_U16 ( .A(intadd_24_A_2_), .B(intadd_24_B_2_), .CI(
        intadd_24_n16), .CO(intadd_24_n15), .S(intadd_24_SUM_2_) );
  fad1_hd intadd_24_U15 ( .A(intadd_24_A_3_), .B(intadd_24_B_3_), .CI(
        intadd_24_n15), .CO(intadd_24_n14), .S(intadd_24_SUM_3_) );
  fad1_hd intadd_24_U14 ( .A(intadd_24_A_4_), .B(intadd_24_B_4_), .CI(
        intadd_24_n14), .CO(intadd_24_n13), .S(intadd_24_SUM_4_) );
  fad1_hd intadd_24_U13 ( .A(intadd_24_A_5_), .B(intadd_24_B_5_), .CI(
        intadd_24_n13), .CO(intadd_24_n12), .S(intadd_24_SUM_5_) );
  fad1_hd intadd_24_U12 ( .A(intadd_24_A_6_), .B(intadd_24_B_6_), .CI(
        intadd_24_n12), .CO(intadd_24_n11), .S(intadd_24_SUM_6_) );
  fad1_hd intadd_24_U11 ( .A(intadd_24_A_7_), .B(intadd_24_B_7_), .CI(
        intadd_24_n11), .CO(intadd_24_n10), .S(intadd_24_SUM_7_) );
  fad1_hd intadd_24_U10 ( .A(intadd_24_A_8_), .B(intadd_24_B_8_), .CI(
        intadd_24_n10), .CO(intadd_24_n9), .S(intadd_24_SUM_8_) );
  fad1_hd intadd_24_U9 ( .A(intadd_24_A_9_), .B(intadd_24_B_9_), .CI(
        intadd_24_n9), .CO(intadd_24_n8), .S(intadd_24_SUM_9_) );
  fad1_hd intadd_24_U8 ( .A(intadd_24_A_10_), .B(intadd_24_B_10_), .CI(
        intadd_24_n8), .CO(intadd_24_n7), .S(intadd_24_SUM_10_) );
  fad1_hd intadd_24_U7 ( .A(intadd_24_A_11_), .B(intadd_24_B_11_), .CI(
        intadd_24_n7), .CO(intadd_24_n6), .S(intadd_24_SUM_11_) );
  fad1_hd intadd_24_U6 ( .A(intadd_24_A_12_), .B(intadd_24_B_12_), .CI(
        intadd_24_n6), .CO(intadd_24_n5), .S(intadd_24_SUM_12_) );
  fad1_hd intadd_24_U5 ( .A(intadd_24_A_13_), .B(intadd_24_B_13_), .CI(
        intadd_24_n5), .CO(intadd_24_n4), .S(intadd_24_SUM_13_) );
  fad1_hd intadd_24_U4 ( .A(intadd_26_n1), .B(intadd_24_B_14_), .CI(
        intadd_24_n4), .CO(intadd_24_n3), .S(intadd_24_SUM_14_) );
  fad1_hd intadd_24_U3 ( .A(intadd_24_A_15_), .B(intadd_24_B_15_), .CI(
        intadd_24_n3), .CO(intadd_24_n2), .S(intadd_24_SUM_15_) );
  fad1_hd intadd_25_U13 ( .A(intadd_25_A_0_), .B(intadd_25_B_0_), .CI(
        intadd_25_CI), .CO(intadd_25_n12), .S(intadd_25_SUM_0_) );
  fad1_hd intadd_25_U12 ( .A(intadd_25_A_1_), .B(intadd_25_B_1_), .CI(
        intadd_25_n12), .CO(intadd_25_n11), .S(intadd_25_SUM_1_) );
  fad1_hd intadd_25_U11 ( .A(intadd_25_A_2_), .B(intadd_25_B_2_), .CI(
        intadd_25_n11), .CO(intadd_25_n10), .S(intadd_25_SUM_2_) );
  fad1_hd intadd_25_U10 ( .A(intadd_25_A_3_), .B(intadd_25_B_3_), .CI(
        intadd_25_n10), .CO(intadd_25_n9), .S(intadd_25_SUM_3_) );
  fad1_hd intadd_25_U9 ( .A(intadd_25_A_4_), .B(intadd_25_B_4_), .CI(
        intadd_25_n9), .CO(intadd_25_n8), .S(intadd_25_SUM_4_) );
  fad1_hd intadd_25_U8 ( .A(intadd_25_A_5_), .B(intadd_25_B_5_), .CI(
        intadd_25_n8), .CO(intadd_25_n7), .S(intadd_25_SUM_5_) );
  fad1_hd intadd_25_U7 ( .A(intadd_25_A_6_), .B(intadd_25_B_6_), .CI(
        intadd_25_n7), .CO(intadd_25_n6), .S(intadd_25_SUM_6_) );
  fad1_hd intadd_25_U6 ( .A(intadd_25_A_7_), .B(intadd_25_B_7_), .CI(
        intadd_25_n6), .CO(intadd_25_n5), .S(intadd_25_SUM_7_) );
  fad1_hd intadd_25_U5 ( .A(intadd_25_A_8_), .B(intadd_25_B_8_), .CI(
        intadd_25_n5), .CO(intadd_25_n4), .S(intadd_25_SUM_8_) );
  fad1_hd intadd_25_U4 ( .A(intadd_25_A_9_), .B(intadd_25_B_9_), .CI(
        intadd_25_n4), .CO(intadd_25_n3), .S(intadd_25_SUM_9_) );
  fad1_hd intadd_25_U3 ( .A(intadd_25_A_10_), .B(intadd_25_B_10_), .CI(
        intadd_25_n3), .CO(intadd_25_n2), .S(intadd_25_SUM_10_) );
  fad1_hd intadd_25_U2 ( .A(intadd_25_A_11_), .B(intadd_25_B_11_), .CI(
        intadd_25_n2), .CO(intadd_25_n1), .S(intadd_25_SUM_11_) );
  fad1_hd intadd_26_U12 ( .A(intadd_26_A_0_), .B(intadd_26_B_0_), .CI(
        intadd_26_CI), .CO(intadd_26_n11), .S(intadd_24_A_3_) );
  fad1_hd intadd_26_U11 ( .A(intadd_26_A_1_), .B(intadd_26_B_1_), .CI(
        intadd_26_n11), .CO(intadd_26_n10), .S(intadd_24_A_4_) );
  fad1_hd intadd_26_U10 ( .A(intadd_26_A_2_), .B(intadd_26_B_2_), .CI(
        intadd_26_n10), .CO(intadd_26_n9), .S(intadd_24_A_5_) );
  fad1_hd intadd_26_U9 ( .A(intadd_26_A_3_), .B(intadd_25_SUM_0_), .CI(
        intadd_26_n9), .CO(intadd_26_n8), .S(intadd_24_A_6_) );
  fad1_hd intadd_26_U8 ( .A(intadd_25_SUM_1_), .B(intadd_26_B_4_), .CI(
        intadd_26_n8), .CO(intadd_26_n7), .S(intadd_24_A_7_) );
  fad1_hd intadd_26_U7 ( .A(intadd_26_A_5_), .B(intadd_25_SUM_2_), .CI(
        intadd_26_n7), .CO(intadd_26_n6), .S(intadd_24_A_8_) );
  fad1_hd intadd_26_U6 ( .A(intadd_26_A_6_), .B(intadd_25_SUM_3_), .CI(
        intadd_26_n6), .CO(intadd_26_n5), .S(intadd_24_A_9_) );
  fad1_hd intadd_26_U5 ( .A(intadd_26_A_7_), .B(intadd_25_SUM_4_), .CI(
        intadd_26_n5), .CO(intadd_26_n4), .S(intadd_24_A_10_) );
  fad1_hd intadd_26_U4 ( .A(intadd_26_A_8_), .B(intadd_25_SUM_5_), .CI(
        intadd_26_n4), .CO(intadd_26_n3), .S(intadd_24_A_11_) );
  fad1_hd intadd_26_U3 ( .A(intadd_25_SUM_6_), .B(intadd_26_B_9_), .CI(
        intadd_26_n3), .CO(intadd_26_n2), .S(intadd_24_A_12_) );
  fad1_hd intadd_26_U2 ( .A(intadd_26_A_10_), .B(intadd_25_SUM_7_), .CI(
        intadd_26_n2), .CO(intadd_26_n1), .S(intadd_24_B_13_) );
  fad1_hd intadd_27_U12 ( .A(intadd_27_A_0_), .B(intadd_27_B_0_), .CI(
        intadd_27_CI), .CO(intadd_27_n11), .S(intadd_27_SUM_0_) );
  fad1_hd intadd_27_U11 ( .A(intadd_27_A_1_), .B(intadd_27_B_1_), .CI(
        intadd_27_n11), .CO(intadd_27_n10), .S(intadd_27_SUM_1_) );
  fad1_hd intadd_27_U10 ( .A(intadd_27_A_2_), .B(intadd_27_B_2_), .CI(
        intadd_27_n10), .CO(intadd_27_n9), .S(intadd_27_SUM_2_) );
  fad1_hd intadd_27_U9 ( .A(intadd_27_A_3_), .B(intadd_27_B_3_), .CI(
        intadd_27_n9), .CO(intadd_27_n8), .S(intadd_27_SUM_3_) );
  fad1_hd intadd_27_U8 ( .A(intadd_27_A_4_), .B(intadd_27_B_4_), .CI(
        intadd_27_n8), .CO(intadd_27_n7), .S(intadd_27_SUM_4_) );
  fad1_hd intadd_27_U7 ( .A(intadd_27_A_5_), .B(intadd_27_B_5_), .CI(
        intadd_27_n7), .CO(intadd_27_n6), .S(intadd_27_SUM_5_) );
  fad1_hd intadd_27_U6 ( .A(intadd_27_A_6_), .B(intadd_27_B_6_), .CI(
        intadd_27_n6), .CO(intadd_27_n5), .S(intadd_27_SUM_6_) );
  fad1_hd intadd_27_U5 ( .A(intadd_27_A_7_), .B(intadd_27_B_7_), .CI(
        intadd_27_n5), .CO(intadd_27_n4), .S(intadd_27_SUM_7_) );
  fad1_hd intadd_27_U4 ( .A(intadd_27_A_8_), .B(intadd_27_B_8_), .CI(
        intadd_27_n4), .CO(intadd_27_n3), .S(intadd_27_SUM_8_) );
  fad1_hd intadd_27_U3 ( .A(intadd_27_A_9_), .B(intadd_27_B_9_), .CI(
        intadd_27_n3), .CO(intadd_27_n2), .S(intadd_27_SUM_9_) );
  fad1_hd intadd_28_U10 ( .A(a_m[2]), .B(intadd_28_B_0_), .CI(intadd_28_CI), 
        .CO(intadd_28_n9), .S(intadd_28_SUM_0_) );
  fad1_hd intadd_28_U9 ( .A(intadd_28_A_1_), .B(intadd_28_B_1_), .CI(
        intadd_28_n9), .CO(intadd_28_n8), .S(intadd_27_A_6_) );
  fad1_hd intadd_28_U8 ( .A(intadd_28_A_2_), .B(intadd_28_B_2_), .CI(
        intadd_28_n8), .CO(intadd_28_n7), .S(intadd_27_A_7_) );
  fad1_hd intadd_28_U7 ( .A(intadd_28_A_3_), .B(intadd_28_B_3_), .CI(
        intadd_28_n7), .CO(intadd_28_n6), .S(intadd_27_A_8_) );
  fad1_hd intadd_28_U6 ( .A(intadd_32_n1), .B(intadd_28_B_4_), .CI(
        intadd_28_n6), .CO(intadd_28_n5), .S(intadd_28_SUM_4_) );
  fad1_hd intadd_28_U5 ( .A(intadd_28_A_5_), .B(intadd_28_B_5_), .CI(
        intadd_28_n5), .CO(intadd_28_n4), .S(intadd_28_SUM_5_) );
  fad1_hd intadd_28_U4 ( .A(intadd_28_A_6_), .B(intadd_28_B_6_), .CI(
        intadd_28_n4), .CO(intadd_28_n3), .S(intadd_28_SUM_6_) );
  fad1_hd intadd_28_U3 ( .A(intadd_28_A_7_), .B(intadd_28_B_7_), .CI(
        intadd_28_n3), .CO(intadd_28_n2), .S(intadd_28_SUM_7_) );
  fad1_hd intadd_29_U9 ( .A(a_m[5]), .B(n107), .CI(intadd_29_CI), .CO(
        intadd_29_n8), .S(intadd_29_SUM_0_) );
  fad1_hd intadd_29_U8 ( .A(intadd_29_A_1_), .B(intadd_29_B_1_), .CI(
        intadd_29_n8), .CO(intadd_29_n7), .S(intadd_29_SUM_1_) );
  fad1_hd intadd_29_U7 ( .A(intadd_29_A_2_), .B(intadd_29_B_2_), .CI(
        intadd_29_n7), .CO(intadd_29_n6), .S(intadd_29_SUM_2_) );
  fad1_hd intadd_29_U6 ( .A(intadd_29_A_3_), .B(intadd_29_B_3_), .CI(
        intadd_29_n6), .CO(intadd_29_n5), .S(intadd_29_SUM_3_) );
  fad1_hd intadd_29_U5 ( .A(intadd_29_A_4_), .B(intadd_29_B_4_), .CI(
        intadd_29_n5), .CO(intadd_29_n4), .S(intadd_29_SUM_4_) );
  fad1_hd intadd_29_U4 ( .A(intadd_29_A_5_), .B(intadd_29_B_5_), .CI(
        intadd_29_n4), .CO(intadd_29_n3), .S(intadd_29_SUM_5_) );
  fad1_hd intadd_29_U3 ( .A(intadd_29_A_6_), .B(intadd_29_B_6_), .CI(
        intadd_29_n3), .CO(intadd_29_n2), .S(intadd_29_SUM_6_) );
  fad1_hd intadd_29_U2 ( .A(intadd_29_A_7_), .B(intadd_29_B_7_), .CI(
        intadd_29_n2), .CO(intadd_29_n1), .S(intadd_29_SUM_7_) );
  fad1_hd intadd_30_U7 ( .A(intadd_30_A_0_), .B(intadd_30_B_0_), .CI(
        intadd_30_CI), .CO(intadd_30_n6), .S(intadd_30_SUM_0_) );
  fad1_hd intadd_30_U6 ( .A(intadd_30_A_1_), .B(intadd_30_B_1_), .CI(
        intadd_30_n6), .CO(intadd_30_n5), .S(intadd_30_SUM_1_) );
  fad1_hd intadd_30_U5 ( .A(intadd_30_A_2_), .B(intadd_30_B_2_), .CI(
        intadd_30_n5), .CO(intadd_30_n4), .S(intadd_30_SUM_2_) );
  fad1_hd intadd_30_U4 ( .A(intadd_30_A_3_), .B(intadd_30_B_3_), .CI(
        intadd_30_n4), .CO(intadd_30_n3), .S(intadd_30_SUM_3_) );
  fad1_hd intadd_30_U3 ( .A(intadd_30_A_4_), .B(intadd_30_B_4_), .CI(
        intadd_30_n3), .CO(intadd_30_n2), .S(intadd_30_SUM_4_) );
  fad1_hd intadd_31_U6 ( .A(intadd_31_A_0_), .B(intadd_31_B_0_), .CI(
        intadd_31_CI), .CO(intadd_31_n5), .S(intadd_31_SUM_0_) );
  fad1_hd intadd_31_U5 ( .A(intadd_31_A_1_), .B(intadd_31_B_1_), .CI(
        intadd_31_n5), .CO(intadd_31_n4), .S(intadd_31_SUM_1_) );
  fad1_hd intadd_31_U4 ( .A(intadd_31_A_2_), .B(intadd_31_B_2_), .CI(
        intadd_31_n4), .CO(intadd_31_n3), .S(intadd_31_SUM_2_) );
  fad1_hd intadd_31_U3 ( .A(intadd_31_A_3_), .B(intadd_31_B_3_), .CI(
        intadd_31_n3), .CO(intadd_31_n2), .S(intadd_31_SUM_3_) );
  fad1_hd intadd_32_U4 ( .A(n106), .B(intadd_32_B_0_), .CI(intadd_32_CI), .CO(
        intadd_32_n3), .S(intadd_28_B_1_) );
  fad1_hd intadd_32_U3 ( .A(intadd_32_A_1_), .B(intadd_32_B_1_), .CI(
        intadd_32_n3), .CO(intadd_32_n2), .S(intadd_28_A_2_) );
  fad1_hd intadd_32_U2 ( .A(intadd_32_A_2_), .B(intadd_32_B_2_), .CI(
        intadd_32_n2), .CO(intadd_32_n1), .S(intadd_28_A_3_) );
  fad1_hd intadd_33_U4 ( .A(intadd_33_A_0_), .B(intadd_33_B_0_), .CI(
        intadd_33_CI), .CO(intadd_33_n3), .S(intadd_33_SUM_0_) );
  fad1_hd intadd_33_U3 ( .A(intadd_33_A_1_), .B(intadd_33_B_1_), .CI(
        intadd_33_n3), .CO(intadd_33_n2), .S(intadd_33_SUM_1_) );
  fad1_hd intadd_34_U4 ( .A(intadd_34_A_0_), .B(intadd_34_B_0_), .CI(
        intadd_34_CI), .CO(intadd_34_n3), .S(intadd_34_SUM_0_) );
  fad1_hd intadd_34_U3 ( .A(intadd_34_A_1_), .B(intadd_34_B_1_), .CI(
        intadd_34_n3), .CO(intadd_34_n2), .S(intadd_34_SUM_1_) );
  fad1_hd intadd_34_U2 ( .A(intadd_34_A_2_), .B(intadd_34_B_2_), .CI(
        intadd_34_n2), .CO(intadd_34_n1), .S(intadd_34_SUM_2_) );
  fad1_hd intadd_35_U4 ( .A(intadd_35_A_0_), .B(intadd_35_B_0_), .CI(
        intadd_30_SUM_1_), .CO(intadd_35_n3), .S(intadd_35_SUM_0_) );
  fad1_hd intadd_35_U3 ( .A(intadd_30_SUM_2_), .B(intadd_35_B_1_), .CI(
        intadd_35_n3), .CO(intadd_35_n2), .S(intadd_35_SUM_1_) );
  fad1_hd intadd_36_U4 ( .A(intadd_29_SUM_5_), .B(intadd_36_B_0_), .CI(
        intadd_36_CI), .CO(intadd_36_n3), .S(intadd_36_SUM_0_) );
  fad1_hd intadd_36_U3 ( .A(intadd_29_SUM_6_), .B(intadd_36_B_1_), .CI(
        intadd_36_n3), .CO(intadd_36_n2), .S(intadd_36_SUM_1_) );
  fad1_hd intadd_37_U4 ( .A(intadd_37_A_0_), .B(intadd_37_B_0_), .CI(
        intadd_37_CI), .CO(intadd_37_n3), .S(intadd_37_SUM_0_) );
  fad1_hd intadd_37_U3 ( .A(intadd_37_A_1_), .B(intadd_37_B_1_), .CI(
        intadd_37_n3), .CO(intadd_37_n2), .S(intadd_37_SUM_1_) );
  fad1_hd intadd_38_U4 ( .A(intadd_29_SUM_2_), .B(intadd_38_B_0_), .CI(
        intadd_38_CI), .CO(intadd_38_n3), .S(intadd_38_SUM_0_) );
  fad1_hd intadd_38_U3 ( .A(intadd_29_SUM_3_), .B(intadd_38_B_1_), .CI(
        intadd_38_n3), .CO(intadd_38_n2), .S(intadd_38_SUM_1_) );
  fad1_hd intadd_38_U2 ( .A(intadd_29_SUM_4_), .B(intadd_38_B_2_), .CI(
        intadd_38_n2), .CO(intadd_38_n1), .S(intadd_38_SUM_2_) );
  fad1_hd intadd_39_U4 ( .A(intadd_39_A_0_), .B(intadd_25_SUM_9_), .CI(
        intadd_39_CI), .CO(intadd_39_n3), .S(intadd_24_A_15_) );
  fad1_hd intadd_39_U3 ( .A(intadd_39_A_1_), .B(intadd_25_SUM_10_), .CI(
        intadd_39_n3), .CO(intadd_39_n2), .S(intadd_24_A_16_) );
  fad1_hd intadd_39_U2 ( .A(intadd_25_SUM_11_), .B(intadd_39_B_2_), .CI(
        intadd_39_n2), .CO(intadd_39_n1), .S(intadd_39_SUM_2_) );
  fad1_hd intadd_20_U38 ( .A(intadd_20_A_0_), .B(intadd_20_B_0_), .CI(
        intadd_20_CI), .CO(intadd_20_n37), .S(intadd_20_SUM_0_) );
  fad1_hd intadd_20_U37 ( .A(intadd_20_A_1_), .B(intadd_20_B_1_), .CI(
        intadd_20_n37), .CO(intadd_20_n36), .S(intadd_20_SUM_1_) );
  fad1_hd intadd_20_U36 ( .A(intadd_20_A_2_), .B(intadd_20_B_2_), .CI(
        intadd_20_n36), .CO(intadd_20_n35), .S(intadd_20_SUM_2_) );
  fad1_hd intadd_20_U35 ( .A(intadd_20_A_3_), .B(intadd_20_B_3_), .CI(
        intadd_20_n35), .CO(intadd_20_n34), .S(intadd_20_SUM_3_) );
  fad1_hd intadd_20_U34 ( .A(intadd_20_A_4_), .B(intadd_20_B_4_), .CI(
        intadd_20_n34), .CO(intadd_20_n33), .S(intadd_20_SUM_4_) );
  fad1_hd intadd_20_U33 ( .A(intadd_20_A_5_), .B(intadd_20_B_5_), .CI(
        intadd_20_n33), .CO(intadd_20_n32), .S(intadd_20_SUM_5_) );
  fad1_hd intadd_20_U32 ( .A(intadd_20_A_6_), .B(intadd_20_B_6_), .CI(
        intadd_20_n32), .CO(intadd_20_n31), .S(intadd_20_SUM_6_) );
  fad1_hd intadd_20_U31 ( .A(intadd_20_A_7_), .B(intadd_20_B_7_), .CI(
        intadd_20_n31), .CO(intadd_20_n30), .S(intadd_20_SUM_7_) );
  fad1_hd intadd_20_U30 ( .A(intadd_20_A_8_), .B(intadd_20_B_8_), .CI(
        intadd_20_n30), .CO(intadd_20_n29), .S(intadd_20_SUM_8_) );
  fad1_hd intadd_20_U29 ( .A(intadd_20_A_9_), .B(intadd_20_B_9_), .CI(
        intadd_20_n29), .CO(intadd_20_n28), .S(intadd_20_SUM_9_) );
  fad1_hd intadd_20_U28 ( .A(intadd_20_A_10_), .B(intadd_20_B_10_), .CI(
        intadd_20_n28), .CO(intadd_20_n27), .S(intadd_20_SUM_10_) );
  fad1_hd intadd_20_U27 ( .A(intadd_20_A_11_), .B(intadd_20_B_11_), .CI(
        intadd_20_n27), .CO(intadd_20_n26), .S(intadd_20_SUM_11_) );
  fad1_hd intadd_20_U26 ( .A(intadd_20_A_12_), .B(intadd_20_B_12_), .CI(
        intadd_20_n26), .CO(intadd_20_n25), .S(intadd_20_SUM_12_) );
  fad1_hd intadd_20_U25 ( .A(intadd_20_A_13_), .B(intadd_20_B_13_), .CI(
        intadd_20_n25), .CO(intadd_20_n24), .S(intadd_20_SUM_13_) );
  fad1_hd intadd_20_U24 ( .A(intadd_20_A_14_), .B(intadd_20_B_14_), .CI(
        intadd_20_n24), .CO(intadd_20_n23), .S(intadd_20_SUM_14_) );
  fad1_hd intadd_20_U23 ( .A(intadd_20_A_15_), .B(intadd_20_B_15_), .CI(
        intadd_20_n23), .CO(intadd_20_n22), .S(intadd_20_SUM_15_) );
  fad1_hd intadd_20_U22 ( .A(intadd_20_A_16_), .B(intadd_20_B_16_), .CI(
        intadd_20_n22), .CO(intadd_20_n21), .S(intadd_20_SUM_16_) );
  fad1_hd intadd_21_U24 ( .A(intadd_21_A_0_), .B(intadd_21_B_0_), .CI(
        intadd_21_CI), .CO(intadd_21_n23), .S(intadd_21_SUM_0_) );
  fad1_hd intadd_21_U23 ( .A(intadd_21_A_1_), .B(intadd_21_B_1_), .CI(
        intadd_21_n23), .CO(intadd_21_n22), .S(intadd_21_SUM_1_) );
  fad1_hd intadd_21_U22 ( .A(intadd_21_A_2_), .B(intadd_21_B_2_), .CI(
        intadd_21_n22), .CO(intadd_21_n21), .S(intadd_21_SUM_2_) );
  fad1_hd intadd_21_U21 ( .A(intadd_21_A_3_), .B(intadd_21_B_3_), .CI(
        intadd_21_n21), .CO(intadd_21_n20), .S(intadd_21_SUM_3_) );
  fad1_hd intadd_21_U20 ( .A(intadd_21_A_4_), .B(intadd_21_B_4_), .CI(
        intadd_21_n20), .CO(intadd_21_n19), .S(intadd_21_SUM_4_) );
  fad1_hd intadd_21_U19 ( .A(intadd_21_A_5_), .B(intadd_21_B_5_), .CI(
        intadd_21_n19), .CO(intadd_21_n18), .S(intadd_21_SUM_5_) );
  fad1_hd intadd_21_U18 ( .A(intadd_21_A_6_), .B(intadd_21_B_6_), .CI(
        intadd_21_n18), .CO(intadd_21_n17), .S(intadd_21_SUM_6_) );
  fad1_hd intadd_21_U17 ( .A(intadd_21_A_7_), .B(intadd_21_B_7_), .CI(
        intadd_21_n17), .CO(intadd_21_n16), .S(intadd_21_SUM_7_) );
  fad1_hd intadd_21_U16 ( .A(intadd_21_A_8_), .B(intadd_21_B_8_), .CI(
        intadd_21_n16), .CO(intadd_21_n15), .S(intadd_21_SUM_8_) );
  fad1_hd intadd_21_U15 ( .A(intadd_21_A_9_), .B(intadd_21_B_9_), .CI(
        intadd_21_n15), .CO(intadd_21_n14), .S(intadd_21_SUM_9_) );
  fad1_hd intadd_21_U14 ( .A(intadd_21_A_10_), .B(intadd_21_B_10_), .CI(
        intadd_21_n14), .CO(intadd_21_n13), .S(intadd_21_SUM_10_) );
  fad1_hd intadd_21_U13 ( .A(intadd_21_A_11_), .B(intadd_21_B_11_), .CI(
        intadd_21_n13), .CO(intadd_21_n12), .S(intadd_21_SUM_11_) );
  fad1_hd intadd_21_U12 ( .A(intadd_21_A_12_), .B(intadd_21_B_12_), .CI(
        intadd_21_n12), .CO(intadd_21_n11), .S(intadd_21_SUM_12_) );
  fad1_hd intadd_21_U11 ( .A(intadd_21_A_13_), .B(intadd_21_B_13_), .CI(
        intadd_21_n11), .CO(intadd_21_n10), .S(intadd_21_SUM_13_) );
  fad1_hd intadd_21_U10 ( .A(intadd_21_A_14_), .B(intadd_21_B_14_), .CI(
        intadd_21_n10), .CO(intadd_21_n9), .S(intadd_21_SUM_14_) );
  fad1_hd intadd_21_U9 ( .A(intadd_21_A_15_), .B(intadd_21_B_15_), .CI(
        intadd_21_n9), .CO(intadd_21_n8), .S(intadd_21_SUM_15_) );
  fad1_hd intadd_21_U8 ( .A(intadd_21_A_16_), .B(intadd_21_B_16_), .CI(
        intadd_21_n8), .CO(intadd_21_n7), .S(intadd_21_SUM_16_) );
  fad1_hd intadd_21_U7 ( .A(intadd_21_A_17_), .B(intadd_21_B_17_), .CI(
        intadd_21_n7), .CO(intadd_21_n6), .S(intadd_21_SUM_17_) );
  fad1_hd intadd_21_U6 ( .A(intadd_21_A_18_), .B(intadd_21_B_18_), .CI(
        intadd_21_n6), .CO(intadd_21_n5), .S(intadd_21_SUM_18_) );
  fad1_hd intadd_21_U5 ( .A(intadd_21_A_19_), .B(intadd_21_B_19_), .CI(
        intadd_21_n5), .CO(intadd_21_n4), .S(intadd_21_SUM_19_) );
  fad1_hd intadd_21_U4 ( .A(intadd_21_A_20_), .B(intadd_21_B_20_), .CI(
        intadd_21_n4), .CO(intadd_21_n3), .S(intadd_21_SUM_20_) );
  fad1_hd intadd_21_U3 ( .A(intadd_21_A_21_), .B(intadd_21_B_21_), .CI(
        intadd_21_n3), .CO(intadd_21_n2), .S(intadd_21_SUM_21_) );
  fad1_hd intadd_21_U2 ( .A(intadd_22_n1), .B(intadd_21_B_22_), .CI(
        intadd_21_n2), .CO(intadd_21_n1), .S(intadd_21_SUM_22_) );
  fad1_hd intadd_22_U20 ( .A(intadd_22_A_0_), .B(intadd_22_B_0_), .CI(
        intadd_22_CI), .CO(intadd_22_n19), .S(intadd_21_A_3_) );
  fad1_hd intadd_22_U19 ( .A(intadd_22_A_1_), .B(intadd_22_B_1_), .CI(
        intadd_22_n19), .CO(intadd_22_n18), .S(intadd_21_A_4_) );
  fad1_hd intadd_22_U17 ( .A(intadd_22_A_3_), .B(intadd_22_B_3_), .CI(
        intadd_22_n17), .CO(intadd_22_n16), .S(intadd_21_A_6_) );
  fad1_hd intadd_22_U16 ( .A(intadd_22_A_4_), .B(intadd_22_B_4_), .CI(
        intadd_22_n16), .CO(intadd_22_n15), .S(intadd_21_A_7_) );
  fad1_hd intadd_22_U15 ( .A(intadd_22_A_5_), .B(intadd_22_B_5_), .CI(
        intadd_22_n15), .CO(intadd_22_n14), .S(intadd_21_A_8_) );
  fad1_hd intadd_22_U14 ( .A(intadd_22_A_6_), .B(intadd_22_B_6_), .CI(
        intadd_22_n14), .CO(intadd_22_n13), .S(intadd_21_A_9_) );
  fad1_hd intadd_22_U13 ( .A(intadd_22_A_7_), .B(intadd_22_B_7_), .CI(
        intadd_22_n13), .CO(intadd_22_n12), .S(intadd_21_A_10_) );
  fad1_hd intadd_22_U12 ( .A(intadd_22_A_8_), .B(intadd_22_B_8_), .CI(
        intadd_22_n12), .CO(intadd_22_n11), .S(intadd_21_A_11_) );
  fad1_hd intadd_22_U11 ( .A(intadd_22_A_9_), .B(intadd_22_B_9_), .CI(
        intadd_22_n11), .CO(intadd_22_n10), .S(intadd_21_A_12_) );
  fad1_hd intadd_22_U10 ( .A(intadd_22_A_10_), .B(intadd_22_B_10_), .CI(
        intadd_22_n10), .CO(intadd_22_n9), .S(intadd_21_B_13_) );
  fad1_hd intadd_22_U7 ( .A(intadd_22_A_13_), .B(intadd_22_B_13_), .CI(
        intadd_22_n7), .CO(intadd_22_n6), .S(intadd_21_A_16_) );
  fad1_hd intadd_22_U6 ( .A(intadd_22_A_14_), .B(intadd_22_B_14_), .CI(
        intadd_22_n6), .CO(intadd_22_n5), .S(intadd_21_B_17_) );
  fad1_hd intadd_22_U5 ( .A(intadd_22_A_15_), .B(intadd_22_B_15_), .CI(
        intadd_22_n5), .CO(intadd_22_n4), .S(intadd_21_B_18_) );
  fad1_hd intadd_22_U4 ( .A(intadd_22_A_16_), .B(intadd_22_B_16_), .CI(
        intadd_22_n4), .CO(intadd_22_n3), .S(intadd_21_B_19_) );
  fd1qd1_hd b_m_reg_1_ ( .D(n307), .CK(i_CLK), .Q(b_m[1]) );
  fad1_hd intadd_30_U2 ( .A(intadd_30_A_5_), .B(intadd_30_B_5_), .CI(
        intadd_30_n2), .CO(intadd_30_n1), .S(intadd_30_SUM_5_) );
  fad1_hd intadd_24_U2 ( .A(intadd_24_A_16_), .B(intadd_24_B_16_), .CI(
        intadd_24_n2), .CO(intadd_24_n1), .S(intadd_24_SUM_16_) );
  fad1_hd intadd_31_U2 ( .A(intadd_31_A_4_), .B(intadd_31_B_4_), .CI(
        intadd_31_n2), .CO(intadd_31_n1), .S(intadd_31_SUM_4_) );
  fad1_hd intadd_28_U2 ( .A(intadd_28_A_8_), .B(intadd_28_B_8_), .CI(
        intadd_28_n2), .CO(intadd_28_n1), .S(intadd_28_SUM_8_) );
  fad1_hd intadd_27_U2 ( .A(intadd_27_A_10_), .B(intadd_27_B_10_), .CI(
        intadd_27_n2), .CO(intadd_27_n1), .S(intadd_27_SUM_10_) );
  fad1_hd intadd_33_U2 ( .A(intadd_33_A_2_), .B(intadd_33_B_2_), .CI(
        intadd_33_n2), .CO(intadd_33_n1), .S(intadd_33_SUM_2_) );
  fad1_hd intadd_23_U15 ( .A(intadd_23_B_5_), .B(intadd_23_B_4_), .CI(
        intadd_23_n15), .CO(intadd_23_n14), .S(intadd_23_SUM_4_) );
  fad1_hd intadd_23_U16 ( .A(intadd_23_B_4_), .B(intadd_23_B_3_), .CI(
        intadd_23_n16), .CO(intadd_23_n15), .S(intadd_23_SUM_3_) );
  fad1_hd intadd_23_U18 ( .A(intadd_23_B_2_), .B(intadd_23_B_1_), .CI(
        intadd_23_n18), .CO(intadd_23_n17), .S(intadd_23_SUM_1_) );
  fad1_hd intadd_23_U17 ( .A(intadd_23_B_3_), .B(intadd_23_B_2_), .CI(
        intadd_23_n17), .CO(intadd_23_n16), .S(intadd_23_SUM_2_) );
  fad1_hd intadd_23_U19 ( .A(intadd_23_B_1_), .B(intadd_23_B_0_), .CI(
        intadd_23_CI), .CO(intadd_23_n18), .S(intadd_23_SUM_0_) );
  fad2_hd intadd_20_U12 ( .A(intadd_20_A_26_), .B(intadd_28_n1), .CI(
        intadd_20_n12), .CO(intadd_20_n11), .S(N212) );
  fad2_hd intadd_20_U10 ( .A(intadd_31_SUM_4_), .B(intadd_20_B_28_), .CI(
        intadd_20_n10), .CO(intadd_20_n9), .S(N214) );
  fad2_hd intadd_20_U8 ( .A(intadd_20_A_30_), .B(intadd_20_B_30_), .CI(
        intadd_20_n8), .CO(intadd_20_n7), .S(N216) );
  fad2_hd intadd_20_U4 ( .A(intadd_20_A_34_), .B(intadd_20_B_34_), .CI(
        intadd_20_n4), .CO(intadd_20_n3), .S(N220) );
  fad1_hd intadd_35_U2 ( .A(intadd_30_SUM_3_), .B(intadd_35_B_2_), .CI(
        intadd_35_n2), .CO(intadd_35_n1), .S(intadd_35_SUM_2_) );
  fad2_hd intadd_20_U18 ( .A(intadd_20_A_20_), .B(intadd_20_B_20_), .CI(
        intadd_20_n18), .CO(intadd_20_n17), .S(N206) );
  fad1_hd intadd_23_U14 ( .A(intadd_23_B_6_), .B(intadd_23_B_5_), .CI(
        intadd_23_n14), .CO(intadd_23_n13), .S(intadd_23_SUM_5_) );
  fad1_hd intadd_36_U2 ( .A(intadd_29_SUM_7_), .B(intadd_36_B_2_), .CI(
        intadd_36_n2), .CO(intadd_36_n1), .S(intadd_36_SUM_2_) );
  fad1_hd intadd_37_U2 ( .A(intadd_37_A_2_), .B(intadd_37_B_2_), .CI(
        intadd_37_n2), .CO(intadd_37_n1), .S(intadd_37_SUM_2_) );
  fad1_hd intadd_20_U20 ( .A(intadd_20_A_18_), .B(intadd_20_B_18_), .CI(
        intadd_20_n20), .CO(intadd_20_n19), .S(N204) );
  fd1qd1_hd sticky_reg ( .D(n283), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n350), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd o_Z_STB_reg ( .D(n358), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_reg_30_ ( .D(n230), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n355), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n310), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n331), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n334), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n337), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n340), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd round_bit_reg ( .D(n284), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd z_reg_31_ ( .D(n229), .CK(i_CLK), .Q(z[31]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n308), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd z_reg_21_ ( .D(n239), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n240), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n241), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n242), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_25_ ( .D(n235), .CK(i_CLK), .Q(z[25]) );
  fd1qd1_hd z_reg_22_ ( .D(n238), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd state_reg_3_ ( .D(n357), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd state_reg_2_ ( .D(n351), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_1_ ( .D(n352), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n353), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd z_reg_15_ ( .D(n245), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n246), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_11_ ( .D(n249), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n250), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_7_ ( .D(n253), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n254), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_3_ ( .D(n257), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_2_ ( .D(n258), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_17_ ( .D(n243), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n244), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_13_ ( .D(n247), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n248), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_9_ ( .D(n251), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n252), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_5_ ( .D(n255), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_4_ ( .D(n256), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_1_ ( .D(n259), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_0_ ( .D(n260), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_28_ ( .D(n232), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n234), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n236), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n237), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n336), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n342), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n348), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd z_reg_29_ ( .D(n231), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n233), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n328), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n347), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n329), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n332), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n349), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n335), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n346), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n341), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n344), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n354), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n345), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n333), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n339), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n343), .CK(i_CLK), .Q(a_m[6]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n330), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n338), .CK(i_CLK), .Q(a_m[11]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n17), .CK(i_CLK), .Q(b[28]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n5), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n2), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n6), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n12), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n12), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n4), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n476), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n6), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n16), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd z_s_reg ( .D(N35), .E(n491), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd product_reg_2_ ( .D(N176), .E(n491), .CK(i_CLK), .Q(product[2])
         );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n501), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n7), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n7), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n11), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n11), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n9), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n3), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n476), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n4), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n12), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n4), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1434), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n5), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n16), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n17), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n7), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n6), .CK(i_CLK), .Q(b[23]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n16), .CK(i_CLK), .Q(b[22]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n7), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n1), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n13), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n17), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n6), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n15), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n501), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n501), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n17), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n500), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n500), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n17), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n13), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n7), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n15), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n3), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n3), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n13), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n2), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n2), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n16), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n16), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n6), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n15), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n2), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n5), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n146), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n11), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n9), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n4), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n4), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n3), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n12), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n9), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n9), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n3), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n11), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n12), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n12), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n4), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n476), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n11), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n11), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n9), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n3), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1434), .CK(i_CLK), .Q(a_s) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n7), .CK(i_CLK), .Q(b[26]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n5), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n15), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n5), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n15), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n500), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n6), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n2), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n5), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n2), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n15), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n13), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n501), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n501), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n17), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n146), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n13), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n16), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd guard_reg ( .D(n104), .E(n105), .CK(i_CLK), .Q(net908) );
  fd1eqd1_hd product_reg_3_ ( .D(N177), .E(n488), .CK(i_CLK), .Q(product[3])
         );
  fd1eqd1_hd product_reg_4_ ( .D(N178), .E(n491), .CK(i_CLK), .Q(product[4])
         );
  fd1eqd1_hd product_reg_5_ ( .D(N179), .E(n490), .CK(i_CLK), .Q(product[5])
         );
  fd1eqd1_hd product_reg_6_ ( .D(N180), .E(n492), .CK(i_CLK), .Q(product[6])
         );
  fd1eqd1_hd product_reg_7_ ( .D(N181), .E(n493), .CK(i_CLK), .Q(product[7])
         );
  fd1eqd1_hd product_reg_8_ ( .D(N182), .E(n489), .CK(i_CLK), .Q(product[8])
         );
  fd1eqd1_hd product_reg_9_ ( .D(N183), .E(n489), .CK(i_CLK), .Q(product[9])
         );
  fd1eqd1_hd product_reg_10_ ( .D(N184), .E(n496), .CK(i_CLK), .Q(product[10])
         );
  fd1eqd1_hd product_reg_11_ ( .D(N185), .E(n494), .CK(i_CLK), .Q(product[11])
         );
  fd1eqd1_hd z_e_reg_8_ ( .D(N474), .E(n8), .CK(i_CLK), .Q(z_e[8]) );
  fd1eqd1_hd z_e_reg_7_ ( .D(N473), .E(n8), .CK(i_CLK), .Q(z_e[7]) );
  fd1eqd1_hd z_e_reg_6_ ( .D(N472), .E(n8), .CK(i_CLK), .Q(z_e[6]) );
  fd1eqd1_hd z_e_reg_5_ ( .D(N471), .E(n8), .CK(i_CLK), .Q(z_e[5]) );
  fd1eqd1_hd z_e_reg_4_ ( .D(N470), .E(n8), .CK(i_CLK), .Q(z_e[4]) );
  fd1eqd1_hd z_e_reg_3_ ( .D(N469), .E(n1430), .CK(i_CLK), .Q(z_e[3]) );
  fd1eqd1_hd z_e_reg_2_ ( .D(N468), .E(n1430), .CK(i_CLK), .Q(z_e[2]) );
  fd1eqd1_hd z_e_reg_1_ ( .D(N467), .E(n1430), .CK(i_CLK), .Q(z_e[1]) );
  fd1eqd1_hd z_e_reg_0_ ( .D(n1429), .E(n1430), .CK(i_CLK), .Q(z_e[0]) );
  fd1eqd1_hd product_reg_12_ ( .D(N186), .E(n488), .CK(i_CLK), .Q(product[12])
         );
  fd1eqd1_hd z_e_reg_9_ ( .D(N475), .E(n1430), .CK(i_CLK), .Q(z_e[9]) );
  fd1eqd1_hd product_reg_13_ ( .D(N187), .E(n490), .CK(i_CLK), .Q(product[13])
         );
  fd1eqd1_hd product_reg_14_ ( .D(N188), .E(n495), .CK(i_CLK), .Q(product[14])
         );
  fd1eqd1_hd product_reg_15_ ( .D(N189), .E(n493), .CK(i_CLK), .Q(product[15])
         );
  fd1eqd1_hd product_reg_16_ ( .D(N190), .E(n495), .CK(i_CLK), .Q(product[16])
         );
  fd1eqd1_hd product_reg_17_ ( .D(N191), .E(n491), .CK(i_CLK), .Q(product[17])
         );
  fd1eqd1_hd product_reg_18_ ( .D(N192), .E(n490), .CK(i_CLK), .Q(product[18])
         );
  fd1eqd1_hd product_reg_19_ ( .D(N193), .E(n493), .CK(i_CLK), .Q(product[19])
         );
  fd1eqd1_hd product_reg_20_ ( .D(N194), .E(n494), .CK(i_CLK), .Q(product[20])
         );
  fd1eqd1_hd product_reg_21_ ( .D(N195), .E(n488), .CK(i_CLK), .Q(product[21])
         );
  fd1eqd1_hd product_reg_22_ ( .D(N196), .E(n489), .CK(i_CLK), .Q(product[22])
         );
  fd1eqd1_hd product_reg_23_ ( .D(N197), .E(n492), .CK(i_CLK), .Q(product[23])
         );
  fd1eqd1_hd product_reg_24_ ( .D(N198), .E(n495), .CK(i_CLK), .Q(product[24])
         );
  fd1eqd1_hd product_reg_25_ ( .D(N199), .E(n494), .CK(i_CLK), .Q(product[25])
         );
  fd1eqd1_hd product_reg_26_ ( .D(N200), .E(n490), .CK(i_CLK), .Q(product[26])
         );
  fd1eqd1_hd product_reg_27_ ( .D(N201), .E(n491), .CK(i_CLK), .Q(product[27])
         );
  fd1eqd1_hd product_reg_28_ ( .D(N202), .E(n491), .CK(i_CLK), .Q(product[28])
         );
  fd1eqd1_hd product_reg_29_ ( .D(N203), .E(n492), .CK(i_CLK), .Q(product[29])
         );
  fd1eqd1_hd product_reg_30_ ( .D(N204), .E(n488), .CK(i_CLK), .Q(product[30])
         );
  fd1eqd1_hd product_reg_31_ ( .D(N205), .E(n490), .CK(i_CLK), .Q(product[31])
         );
  fd1eqd1_hd product_reg_32_ ( .D(N206), .E(n495), .CK(i_CLK), .Q(product[32])
         );
  fd1eqd1_hd product_reg_33_ ( .D(N207), .E(n495), .CK(i_CLK), .Q(product[33])
         );
  fd1eqd1_hd product_reg_34_ ( .D(N208), .E(n492), .CK(i_CLK), .Q(product[34])
         );
  fd1eqd1_hd product_reg_35_ ( .D(N209), .E(n489), .CK(i_CLK), .Q(product[35])
         );
  fd1eqd1_hd product_reg_36_ ( .D(N210), .E(n488), .CK(i_CLK), .Q(product[36])
         );
  fd1eqd1_hd product_reg_37_ ( .D(N211), .E(n495), .CK(i_CLK), .Q(product[37])
         );
  fd1eqd1_hd product_reg_38_ ( .D(N212), .E(n493), .CK(i_CLK), .Q(product[38])
         );
  fd1eqd1_hd product_reg_39_ ( .D(N213), .E(n493), .CK(i_CLK), .Q(product[39])
         );
  fd1eqd1_hd product_reg_40_ ( .D(N214), .E(n489), .CK(i_CLK), .Q(product[40])
         );
  fd1eqd1_hd product_reg_41_ ( .D(N215), .E(n493), .CK(i_CLK), .Q(product[41])
         );
  fd1eqd1_hd product_reg_42_ ( .D(N216), .E(n494), .CK(i_CLK), .Q(product[42])
         );
  fd1eqd1_hd product_reg_43_ ( .D(N217), .E(n494), .CK(i_CLK), .Q(product[43])
         );
  fd1eqd1_hd product_reg_44_ ( .D(N218), .E(n490), .CK(i_CLK), .Q(product[44])
         );
  fd1eqd1_hd product_reg_45_ ( .D(N219), .E(n489), .CK(i_CLK), .Q(product[45])
         );
  fd1eqd1_hd product_reg_46_ ( .D(N220), .E(n492), .CK(i_CLK), .Q(product[46])
         );
  fd1eqd1_hd product_reg_47_ ( .D(N221), .E(n494), .CK(i_CLK), .Q(product[47])
         );
  fd1eqd1_hd product_reg_48_ ( .D(N222), .E(n492), .CK(i_CLK), .Q(product[48])
         );
  fd1eqd1_hd product_reg_49_ ( .D(N223), .E(n488), .CK(i_CLK), .Q(product[49])
         );
  fad1_hd intadd_23_U2 ( .A(intadd_23_A_17_), .B(intadd_23_B_17_), .CI(
        intadd_23_n2), .CO(intadd_23_n1), .S(intadd_23_SUM_17_) );
  fad1_hd intadd_23_U5 ( .A(intadd_23_B_15_), .B(intadd_23_B_14_), .CI(
        intadd_23_n5), .CO(intadd_23_n4), .S(intadd_23_SUM_14_) );
  fad1_hd intadd_23_U3 ( .A(intadd_23_B_17_), .B(intadd_23_B_16_), .CI(
        intadd_23_n3), .CO(intadd_23_n2), .S(intadd_23_SUM_16_) );
  fad1_hd intadd_23_U8 ( .A(intadd_23_B_12_), .B(intadd_23_B_11_), .CI(
        intadd_23_n8), .CO(intadd_23_n7), .S(intadd_23_SUM_11_) );
  fad1_hd intadd_23_U6 ( .A(intadd_23_B_14_), .B(intadd_23_B_13_), .CI(
        intadd_23_n6), .CO(intadd_23_n5), .S(intadd_23_SUM_13_) );
  fad1_hd intadd_23_U9 ( .A(intadd_23_B_11_), .B(intadd_23_B_10_), .CI(
        intadd_23_n9), .CO(intadd_23_n8), .S(intadd_23_SUM_10_) );
  fad1_hd intadd_23_U10 ( .A(intadd_23_B_10_), .B(intadd_23_B_9_), .CI(
        intadd_23_n10), .CO(intadd_23_n9), .S(intadd_23_SUM_9_) );
  fad1_hd intadd_23_U11 ( .A(intadd_23_B_9_), .B(intadd_23_B_8_), .CI(
        intadd_23_n11), .CO(intadd_23_n10), .S(intadd_23_SUM_8_) );
  fad1_hd intadd_23_U12 ( .A(intadd_23_B_8_), .B(intadd_23_B_7_), .CI(
        intadd_23_n12), .CO(intadd_23_n11), .S(intadd_23_SUM_7_) );
  fad1_hd intadd_23_U13 ( .A(intadd_23_B_7_), .B(intadd_23_B_6_), .CI(
        intadd_23_n13), .CO(intadd_23_n12), .S(intadd_23_SUM_6_) );
  fad1_hd intadd_23_U4 ( .A(intadd_23_B_16_), .B(intadd_23_B_15_), .CI(
        intadd_23_n4), .CO(intadd_23_n3), .S(intadd_23_SUM_15_) );
  fad1_hd intadd_23_U7 ( .A(intadd_23_B_13_), .B(intadd_23_B_12_), .CI(
        intadd_23_n7), .CO(intadd_23_n6), .S(intadd_23_SUM_12_) );
  fad1_hd intadd_20_U19 ( .A(intadd_20_A_19_), .B(intadd_20_B_19_), .CI(
        intadd_20_n19), .CO(intadd_20_n18), .S(N205) );
  fad1_hd intadd_20_U17 ( .A(intadd_20_A_21_), .B(intadd_20_B_21_), .CI(
        intadd_20_n17), .CO(intadd_20_n16), .S(N207) );
  fad1_hd intadd_20_U9 ( .A(intadd_20_A_29_), .B(intadd_31_n1), .CI(
        intadd_20_n9), .CO(intadd_20_n8), .S(N215) );
  fad1_hd intadd_20_U7 ( .A(intadd_20_A_31_), .B(intadd_20_B_31_), .CI(
        intadd_20_n7), .CO(intadd_20_n6), .S(N217) );
  fad4_hd intadd_20_U14 ( .A(intadd_20_A_24_), .B(intadd_20_B_24_), .CI(
        intadd_20_n14), .CO(intadd_20_n13), .S(N210) );
  fad4_hd intadd_20_U13 ( .A(intadd_28_SUM_8_), .B(intadd_20_B_25_), .CI(
        intadd_20_n13), .CO(intadd_20_n12), .S(N211) );
  fad1_hd intadd_20_U21 ( .A(intadd_20_A_17_), .B(intadd_20_B_17_), .CI(
        intadd_20_n21), .CO(intadd_20_n20), .S(N203) );
  fad1_hd intadd_20_U6 ( .A(intadd_33_SUM_2_), .B(intadd_20_B_32_), .CI(
        intadd_20_n6), .CO(intadd_20_n5), .S(N218) );
  fad1_hd intadd_20_U2 ( .A(intadd_20_A_36_), .B(intadd_20_B_36_), .CI(
        intadd_20_n2), .CO(intadd_20_n1), .S(N222) );
  fad1_hd intadd_22_U9 ( .A(intadd_22_A_11_), .B(intadd_22_B_11_), .CI(
        intadd_22_n9), .CO(intadd_22_n8), .S(intadd_21_B_14_) );
  fad1_hd intadd_22_U2 ( .A(intadd_22_A_18_), .B(intadd_22_B_18_), .CI(
        intadd_22_n2), .CO(intadd_22_n1), .S(intadd_21_B_21_) );
  fad2_hd intadd_20_U15 ( .A(intadd_20_A_23_), .B(intadd_27_n1), .CI(
        intadd_20_n15), .CO(intadd_20_n14), .S(N209) );
  fad2_hd intadd_20_U16 ( .A(intadd_27_SUM_10_), .B(intadd_20_B_22_), .CI(
        intadd_20_n16), .CO(intadd_20_n15), .S(N208) );
  fad2_hd intadd_20_U5 ( .A(intadd_20_A_33_), .B(intadd_33_n1), .CI(
        intadd_20_n5), .CO(intadd_20_n4), .S(N219) );
  oa22ad1_hd U367 ( .A(n606), .B(a_m[9]), .C(a_m[9]), .D(n608), .Y(n700) );
  nr3d2_hd U368 ( .A(n700), .B(n699), .C(n698), .Y(n967) );
  fad1_hd U369 ( .A(intadd_22_A_12_), .B(intadd_22_B_12_), .CI(intadd_22_n8), 
        .CO(intadd_22_n7), .S(intadd_21_B_15_) );
  fad2_hd U370 ( .A(intadd_20_A_35_), .B(intadd_20_B_35_), .CI(intadd_20_n3), 
        .CO(intadd_20_n2), .S(N221) );
  clknd2d1_hd U371 ( .A(n703), .B(n702), .Y(n713) );
  nid2_hd U372 ( .A(n967), .Y(n410) );
  ivd1_hd U373 ( .A(intadd_21_n1), .Y(intadd_20_A_17_) );
  fad2_hd U374 ( .A(intadd_22_A_17_), .B(intadd_22_B_17_), .CI(intadd_22_n3), 
        .CO(intadd_22_n2), .S(intadd_21_A_20_) );
  nid1_hd U375 ( .A(n419), .Y(n421) );
  clknd2d1_hd U376 ( .A(n746), .B(n747), .Y(n759) );
  nid1_hd U377 ( .A(n464), .Y(n463) );
  clknd2d1_hd U378 ( .A(n719), .B(n720), .Y(n730) );
  clknd2d1_hd U379 ( .A(n125), .B(n728), .Y(n714) );
  ivd1_hd U380 ( .A(n1065), .Y(n847) );
  ivd1_hd U381 ( .A(intadd_23_n1), .Y(n823) );
  scg2d1_hd U382 ( .A(n109), .B(n1065), .C(n847), .D(n126), .Y(n1055) );
  nid1_hd U383 ( .A(n383), .Y(n385) );
  nid1_hd U384 ( .A(n852), .Y(n387) );
  nid1_hd U385 ( .A(n1404), .Y(n472) );
  ivd1_hd U386 ( .A(n92), .Y(n1377) );
  clknd2d1_hd U387 ( .A(n634), .B(n633), .Y(n635) );
  clknd2d1_hd U388 ( .A(n1071), .B(n1074), .Y(n1070) );
  clknd2d1_hd U389 ( .A(n609), .B(b_m[0]), .Y(n858) );
  clknd2d1_hd U390 ( .A(n815), .B(n816), .Y(n833) );
  clknd2d1_hd U391 ( .A(n122), .B(n780), .Y(n778) );
  clknd2d1_hd U392 ( .A(n120), .B(n777), .Y(n779) );
  clknd2d1_hd U393 ( .A(n619), .B(intadd_23_B_5_), .Y(n941) );
  clknd2d1_hd U394 ( .A(n619), .B(intadd_23_B_3_), .Y(intadd_29_B_2_) );
  nid1_hd U395 ( .A(n446), .Y(n444) );
  clknd2d1_hd U396 ( .A(n619), .B(intadd_23_B_2_), .Y(intadd_29_CI) );
  clknd2d1_hd U397 ( .A(n619), .B(n503), .Y(n888) );
  clknd2d1_hd U398 ( .A(n124), .B(n811), .Y(n814) );
  clknd2d1_hd U399 ( .A(n792), .B(n791), .Y(n810) );
  nid1_hd U400 ( .A(n427), .Y(n429) );
  nid1_hd U401 ( .A(n458), .Y(n460) );
  clknd2d1_hd U402 ( .A(n609), .B(n535), .Y(intadd_31_A_0_) );
  nid1_hd U403 ( .A(n1042), .Y(n437) );
  nid1_hd U404 ( .A(n531), .Y(n533) );
  clknd2d1_hd U405 ( .A(b_m[0]), .B(n775), .Y(n777) );
  clknd2d1_hd U406 ( .A(n620), .B(intadd_23_B_11_), .Y(n1000) );
  nid1_hd U407 ( .A(n439), .Y(n441) );
  clknd2d1_hd U408 ( .A(n619), .B(intadd_23_B_9_), .Y(intadd_30_B_1_) );
  nid1_hd U409 ( .A(n1041), .Y(n432) );
  nid1_hd U410 ( .A(n437), .Y(n436) );
  nid1_hd U411 ( .A(b_m[12]), .Y(n552) );
  nid1_hd U412 ( .A(n423), .Y(n424) );
  nid1_hd U413 ( .A(n411), .Y(n412) );
  clknd2d1_hd U414 ( .A(n759), .B(n749), .Y(intadd_26_CI) );
  nid1_hd U415 ( .A(n410), .Y(n407) );
  clknd2d1_hd U416 ( .A(n620), .B(intadd_23_B_14_), .Y(n1027) );
  nid1_hd U417 ( .A(n439), .Y(n440) );
  nid1_hd U418 ( .A(n1064), .Y(n439) );
  nid1_hd U419 ( .A(n446), .Y(n445) );
  nid1_hd U420 ( .A(n431), .Y(n433) );
  nid1_hd U421 ( .A(n423), .Y(n425) );
  nid1_hd U422 ( .A(n418), .Y(n416) );
  nid1_hd U423 ( .A(n418), .Y(n415) );
  clknd2d1_hd U424 ( .A(n730), .B(n722), .Y(intadd_24_CI) );
  nid1_hd U425 ( .A(n403), .Y(n406) );
  clknd2d1_hd U426 ( .A(a_m[11]), .B(n693), .Y(n687) );
  clknd2d1_hd U427 ( .A(n84), .B(n690), .Y(n688) );
  clknd2d1_hd U428 ( .A(n605), .B(n669), .Y(n667) );
  clknd2d1_hd U429 ( .A(n604), .B(n666), .Y(n668) );
  nid1_hd U430 ( .A(n620), .Y(n619) );
  clknd2d1_hd U431 ( .A(n620), .B(intadd_23_B_17_), .Y(n1046) );
  nid1_hd U432 ( .A(n439), .Y(n442) );
  nid1_hd U433 ( .A(n1066), .Y(n446) );
  clknd2d1_hd U434 ( .A(n620), .B(intadd_23_B_15_), .Y(intadd_34_B_1_) );
  clknd2d1_hd U435 ( .A(intadd_33_A_0_), .B(n1027), .Y(n1035) );
  clknd2d1_hd U436 ( .A(n787), .B(n775), .Y(n786) );
  nid1_hd U437 ( .A(n1042), .Y(n438) );
  nid1_hd U438 ( .A(n427), .Y(n430) );
  clknd2d1_hd U439 ( .A(n726), .B(n728), .Y(n977) );
  nid1_hd U440 ( .A(n1022), .Y(n427) );
  nid1_hd U441 ( .A(n1377), .Y(n458) );
  ivd1_hd U442 ( .A(n847), .Y(n196) );
  nid1_hd U443 ( .A(n995), .Y(n419) );
  clknd2d1_hd U444 ( .A(n698), .B(n700), .Y(n697) );
  nid1_hd U445 ( .A(n419), .Y(n422) );
  nid1_hd U446 ( .A(b_m[18]), .Y(n578) );
  nid1_hd U447 ( .A(n411), .Y(n414) );
  nid1_hd U448 ( .A(n936), .Y(n403) );
  nid1_hd U449 ( .A(n968), .Y(n411) );
  nid1_hd U450 ( .A(n399), .Y(n402) );
  nid1_hd U451 ( .A(n935), .Y(n399) );
  clknd2d1_hd U452 ( .A(n674), .B(n676), .Y(n673) );
  clknd2d1_hd U453 ( .A(n643), .B(n653), .Y(n880) );
  scg2d1_hd U454 ( .A(n1068), .B(intadd_23_n1), .C(n823), .D(n804), .Y(n1039)
         );
  nid1_hd U455 ( .A(n573), .Y(n575) );
  nid1_hd U456 ( .A(n909), .Y(n398) );
  nid1_hd U457 ( .A(n560), .Y(n562) );
  nid1_hd U458 ( .A(n518), .Y(n520) );
  clknd2d1_hd U459 ( .A(n123), .B(n700), .Y(n693) );
  nid1_hd U460 ( .A(n522), .Y(n524) );
  nid1_hd U461 ( .A(n909), .Y(n397) );
  clknd2d1_hd U462 ( .A(n679), .B(n678), .Y(n692) );
  nid1_hd U463 ( .A(n518), .Y(n521) );
  nid1_hd U464 ( .A(n397), .Y(n396) );
  nid1_hd U465 ( .A(n394), .Y(n391) );
  nid1_hd U466 ( .A(n394), .Y(n392) );
  nid1_hd U467 ( .A(n469), .Y(n471) );
  nid1_hd U468 ( .A(n398), .Y(n395) );
  nid1_hd U469 ( .A(n1398), .Y(n469) );
  clknd2d1_hd U470 ( .A(n641), .B(a_m[5]), .Y(n645) );
  nid1_hd U471 ( .A(n465), .Y(n467) );
  nid1_hd U472 ( .A(n1387), .Y(n465) );
  nid1_hd U473 ( .A(n1382), .Y(n461) );
  nid1_hd U474 ( .A(n609), .Y(n620) );
  nid1_hd U475 ( .A(a_m[23]), .Y(n609) );
  nid1_hd U476 ( .A(n446), .Y(n443) );
  ad3d1_hd U477 ( .A(n830), .B(n829), .C(n828), .Y(n1064) );
  nid1_hd U478 ( .A(n1041), .Y(n434) );
  nid1_hd U479 ( .A(n438), .Y(n435) );
  nid1_hd U480 ( .A(n1041), .Y(n431) );
  nid1_hd U481 ( .A(n1021), .Y(n423) );
  ivd1_hd U482 ( .A(n1055), .Y(n62) );
  clknd2d1_hd U483 ( .A(n757), .B(n755), .Y(n1014) );
  nid1_hd U484 ( .A(n1022), .Y(n428) );
  nid1_hd U485 ( .A(n1021), .Y(n426) );
  clknd2d1_hd U486 ( .A(n716), .B(n727), .Y(n989) );
  nid1_hd U487 ( .A(n418), .Y(n417) );
  nid1_hd U488 ( .A(n995), .Y(n420) );
  clknd2d1_hd U489 ( .A(n685), .B(n699), .Y(n958) );
  nid1_hd U490 ( .A(n410), .Y(n409) );
  nid1_hd U491 ( .A(n935), .Y(n400) );
  clknd2d1_hd U492 ( .A(n664), .B(n675), .Y(n928) );
  nid1_hd U493 ( .A(n403), .Y(n404) );
  nid1_hd U494 ( .A(n394), .Y(n393) );
  nid1_hd U495 ( .A(n399), .Y(n401) );
  clknd2d1_hd U496 ( .A(intadd_23_A_17_), .B(intadd_23_n1), .Y(n822) );
  ivd1_hd U497 ( .A(n1055), .Y(n61) );
  nid1_hd U498 ( .A(b_m[20]), .Y(n587) );
  nid1_hd U499 ( .A(n586), .Y(n588) );
  nid1_hd U500 ( .A(n577), .Y(n579) );
  nid1_hd U501 ( .A(b_m[17]), .Y(n574) );
  nid1_hd U502 ( .A(b_m[14]), .Y(n561) );
  nid1_hd U503 ( .A(n551), .Y(n553) );
  clknd2d1_hd U504 ( .A(n106), .B(n1406), .Y(n631) );
  nid1_hd U505 ( .A(n472), .Y(n475) );
  nid1_hd U506 ( .A(n531), .Y(n532) );
  nid1_hd U507 ( .A(n390), .Y(n389) );
  nid1_hd U508 ( .A(b_m[6]), .Y(n523) );
  clknd2d1_hd U509 ( .A(n125), .B(n676), .Y(n666) );
  nid1_hd U510 ( .A(b_m[5]), .Y(n519) );
  nid1_hd U511 ( .A(n383), .Y(n386) );
  nid1_hd U512 ( .A(n475), .Y(n474) );
  clknd2d1_hd U513 ( .A(n124), .B(n654), .Y(n641) );
  nid1_hd U514 ( .A(n387), .Y(n390) );
  nid1_hd U515 ( .A(n851), .Y(n384) );
  clknd2d1_hd U516 ( .A(n1408), .B(a_m[1]), .Y(n849) );
  clknd2d1_hd U517 ( .A(a_m[0]), .B(n622), .Y(n629) );
  nid1_hd U518 ( .A(n852), .Y(n388) );
  clknd2d1_hd U519 ( .A(state[2]), .B(n1121), .Y(n621) );
  clknd2d1_hd U520 ( .A(n1415), .B(n1131), .Y(n1132) );
  clknd2d1_hd U521 ( .A(n1346), .B(n1133), .Y(n1130) );
  ivd1_hd U522 ( .A(a_m[8]), .Y(n607) );
  nid1_hd U523 ( .A(n465), .Y(n468) );
  clknd2d1_hd U524 ( .A(n1272), .B(n105), .Y(n1261) );
  clknd2d1_hd U525 ( .A(n1299), .B(n1426), .Y(n1271) );
  nid1_hd U526 ( .A(b_m[20]), .Y(n586) );
  nid1_hd U527 ( .A(b_m[8]), .Y(n531) );
  nid1_hd U528 ( .A(n513), .Y(n512) );
  ivd1_hd U529 ( .A(b_m[7]), .Y(n530) );
  nid1_hd U530 ( .A(b_m[6]), .Y(n522) );
  nid1_hd U531 ( .A(b_m[14]), .Y(n560) );
  nid1_hd U532 ( .A(b_m[12]), .Y(n551) );
  nid1_hd U533 ( .A(b_m[17]), .Y(n573) );
  nid1_hd U534 ( .A(b_m[18]), .Y(n577) );
  ivd1_hd U535 ( .A(b_m[21]), .Y(n595) );
  clknd2d1_hd U536 ( .A(n1126), .B(n1089), .Y(n1143) );
  nid1_hd U537 ( .A(n485), .Y(n483) );
  nid1_hd U538 ( .A(n609), .Y(n616) );
  clknd2d1_hd U539 ( .A(n1432), .B(state[3]), .Y(n1129) );
  clknd2d1_hd U540 ( .A(state[3]), .B(n1116), .Y(n1120) );
  nid1_hd U541 ( .A(n616), .Y(n617) );
  ivd1_hd U542 ( .A(n1117), .Y(n126) );
  clknd2d1_hd U543 ( .A(intadd_23_A_17_), .B(n128), .Y(n1076) );
  clknd2d1_hd U544 ( .A(n620), .B(n1068), .Y(n1071) );
  clknd2d1_hd U545 ( .A(n609), .B(n1069), .Y(n1072) );
  clknd2d1_hd U546 ( .A(n656), .B(n648), .Y(intadd_21_A_0_) );
  clknd2d1_hd U547 ( .A(n641), .B(n635), .Y(n640) );
  clknd2d1_hd U548 ( .A(n639), .B(n640), .Y(intadd_21_CI) );
  nid1_hd U549 ( .A(n498), .Y(n499) );
  clknd2d1_hd U550 ( .A(n107), .B(n626), .Y(n624) );
  clknd2d1_hd U551 ( .A(n107), .B(n628), .Y(n625) );
  clknd2d1_hd U553 ( .A(a_m[0]), .B(b_m[0]), .Y(n626) );
  nid1_hd U554 ( .A(n1398), .Y(n470) );
  nid1_hd U555 ( .A(n1404), .Y(n473) );
  nid1_hd U556 ( .A(n485), .Y(n484) );
  ivd1_hd U557 ( .A(n91), .Y(n92) );
  nid1_hd U558 ( .A(n1332), .Y(n486) );
  nid1_hd U559 ( .A(n1332), .Y(n487) );
  nid1_hd U560 ( .A(n487), .Y(n477) );
  clknd2d1_hd U561 ( .A(n1164), .B(n1161), .Y(n1160) );
  clknd2d1_hd U562 ( .A(n1179), .B(n1178), .Y(n1182) );
  clknd2d1_hd U563 ( .A(n1172), .B(n1168), .Y(n1167) );
  clknd2d1_hd U564 ( .A(n1131), .B(n1130), .Y(n1136) );
  clknd2d1_hd U565 ( .A(n1133), .B(n1132), .Y(n1134) );
  nid1_hd U566 ( .A(n607), .Y(n606) );
  nid1_hd U567 ( .A(n468), .Y(n466) );
  nid1_hd U568 ( .A(n464), .Y(n462) );
  nid1_hd U569 ( .A(n1377), .Y(n459) );
  clknd2d1_hd U570 ( .A(n118), .B(n222), .Y(n1392) );
  ivd1_hd U571 ( .A(n600), .Y(n596) );
  clknd2d1_hd U572 ( .A(n1157), .B(n1154), .Y(n1153) );
  clknd2d1_hd U573 ( .A(state[1]), .B(n1119), .Y(n1297) );
  nid1_hd U574 ( .A(n1308), .Y(n454) );
  clknd2d1_hd U575 ( .A(n1281), .B(n1263), .Y(n1267) );
  clknd2d1_hd U576 ( .A(n201), .B(n1245), .Y(n1249) );
  clknd2d1_hd U577 ( .A(n1281), .B(n1201), .Y(n1205) );
  clknd2d1_hd U578 ( .A(n200), .B(n1228), .Y(n1232) );
  clknd2d1_hd U579 ( .A(n201), .B(n1237), .Y(n1243) );
  clknd2d1_hd U580 ( .A(n200), .B(n1218), .Y(n1225) );
  clknd2d1_hd U581 ( .A(n201), .B(n1274), .Y(n1280) );
  clknd2d1_hd U582 ( .A(n1281), .B(n1192), .Y(n1199) );
  clknd2d1_hd U583 ( .A(n200), .B(n1254), .Y(n1260) );
  nid1_hd U584 ( .A(n1308), .Y(n456) );
  nid1_hd U585 ( .A(n454), .Y(n455) );
  nid1_hd U586 ( .A(n454), .Y(n457) );
  ivd1_hd U587 ( .A(n584), .Y(intadd_23_B_16_) );
  nid1_hd U588 ( .A(n586), .Y(n589) );
  nid1_hd U589 ( .A(n531), .Y(n534) );
  ivd1_hd U590 ( .A(n529), .Y(intadd_23_B_4_) );
  ivd1_hd U591 ( .A(n517), .Y(intadd_23_B_1_) );
  nid1_hd U592 ( .A(b_m[5]), .Y(n518) );
  nid1_hd U593 ( .A(b_m[14]), .Y(intadd_23_B_11_) );
  nid1_hd U594 ( .A(n568), .Y(n567) );
  ivd1_hd U595 ( .A(n512), .Y(intadd_23_B_0_) );
  nid1_hd U596 ( .A(n601), .Y(n600) );
  ivd1_hd U597 ( .A(n594), .Y(intadd_23_A_17_) );
  nid1_hd U598 ( .A(n485), .Y(n482) );
  nid1_hd U599 ( .A(b_m[6]), .Y(intadd_23_B_3_) );
  nid1_hd U600 ( .A(n530), .Y(n529) );
  nid1_hd U601 ( .A(b_m[5]), .Y(intadd_23_B_2_) );
  nid1_hd U602 ( .A(n522), .Y(n525) );
  ivd1_hd U603 ( .A(n539), .Y(intadd_23_B_6_) );
  ivd1_hd U604 ( .A(n544), .Y(intadd_23_B_7_) );
  nid1_hd U605 ( .A(n550), .Y(n549) );
  nid1_hd U606 ( .A(b_m[18]), .Y(intadd_23_B_15_) );
  nid1_hd U607 ( .A(n585), .Y(n584) );
  ivd1_hd U608 ( .A(n558), .Y(intadd_23_B_10_) );
  nid1_hd U609 ( .A(n560), .Y(n563) );
  ivd1_hd U610 ( .A(n507), .Y(n502) );
  nid1_hd U611 ( .A(b_m[8]), .Y(intadd_23_B_5_) );
  nid1_hd U612 ( .A(n540), .Y(n539) );
  nid1_hd U613 ( .A(n486), .Y(n479) );
  nid1_hd U614 ( .A(n551), .Y(n554) );
  ivd1_hd U615 ( .A(n549), .Y(intadd_23_B_8_) );
  nid1_hd U616 ( .A(n559), .Y(n558) );
  nid1_hd U617 ( .A(b_m[12]), .Y(intadd_23_B_9_) );
  nid1_hd U618 ( .A(n486), .Y(n480) );
  ivd1_hd U619 ( .A(n567), .Y(intadd_23_B_12_) );
  ivd1_hd U620 ( .A(n572), .Y(intadd_23_B_13_) );
  nid1_hd U621 ( .A(n573), .Y(n576) );
  nid1_hd U622 ( .A(b_m[17]), .Y(intadd_23_B_14_) );
  nid1_hd U623 ( .A(n577), .Y(n580) );
  nid1_hd U624 ( .A(n486), .Y(n481) );
  nid1_hd U625 ( .A(n508), .Y(n507) );
  nid1_hd U626 ( .A(n595), .Y(n594) );
  nid1_hd U627 ( .A(b_m[20]), .Y(intadd_23_B_17_) );
  nid1_hd U628 ( .A(n487), .Y(n478) );
  clknd2d1_hd U629 ( .A(n1119), .B(n77), .Y(n1416) );
  clknd2d1_hd U630 ( .A(n1121), .B(n1089), .Y(n1356) );
  clknd2d1_hd U631 ( .A(n1087), .B(n1086), .Y(n1146) );
  clknd2d1_hd U632 ( .A(z_e[7]), .B(z_e[8]), .Y(n1145) );
  clknd2d1_hd U633 ( .A(n78), .B(n1125), .Y(n1188) );
  nid1_hd U634 ( .A(n616), .Y(n618) );
  clknd2d1_hd U635 ( .A(state[1]), .B(n1125), .Y(n1148) );
  xo2d1_hd U636 ( .A(intadd_20_n1), .B(n1079), .Y(N223) );
  fad1_hd U637 ( .A(intadd_20_A_27_), .B(intadd_20_B_27_), .CI(intadd_20_n11), 
        .CO(intadd_20_n10), .S(N213) );
  clknd2d1_hd U638 ( .A(z_m[23]), .B(n1423), .Y(n1425) );
  clknd2d1_hd U639 ( .A(n1424), .B(n1297), .Y(n105) );
  nid1_hd U640 ( .A(n1), .Y(n15) );
  nid1_hd U641 ( .A(n1), .Y(n7) );
  nid1_hd U642 ( .A(n1), .Y(n16) );
  nid1_hd U643 ( .A(n1), .Y(n6) );
  nid1_hd U644 ( .A(n146), .Y(n2) );
  nid1_hd U645 ( .A(n146), .Y(n5) );
  nid1_hd U646 ( .A(n1), .Y(n17) );
  clknd2d1_hd U647 ( .A(n194), .B(n1163), .Y(n233) );
  clknd2d1_hd U648 ( .A(n194), .B(n1156), .Y(n231) );
  clknd2d1_hd U649 ( .A(n451), .B(z[23]), .Y(n1175) );
  clknd2d1_hd U650 ( .A(n451), .B(z[24]), .Y(n1173) );
  clknd2d1_hd U651 ( .A(n451), .B(z[26]), .Y(n1165) );
  clknd2d1_hd U652 ( .A(n451), .B(z[28]), .Y(n1158) );
  clknd2d1_hd U653 ( .A(n194), .B(n1171), .Y(n235) );
  clknd2d1_hd U654 ( .A(n453), .B(n1140), .Y(n1141) );
  clknd2d1_hd U655 ( .A(z_e[7]), .B(n1153), .Y(n1151) );
  clknd2d1_hd U656 ( .A(n1351), .B(n138), .Y(n311) );
  clknd2d1_hd U657 ( .A(n1368), .B(n148), .Y(n320) );
  clknd2d1_hd U658 ( .A(n1282), .B(n199), .Y(n1283) );
  clknd2d1_hd U659 ( .A(n1286), .B(n1285), .Y(n1284) );
  clknd2d1_hd U660 ( .A(n1307), .B(n1285), .Y(n1288) );
  clknd2d1_hd U661 ( .A(n1353), .B(n138), .Y(n317) );
  clknd2d1_hd U662 ( .A(n1369), .B(n148), .Y(n326) );
  clknd2d1_hd U663 ( .A(n1420), .B(n1419), .Y(n1417) );
  clknd2d1_hd U664 ( .A(n1360), .B(n1359), .Y(n1357) );
  clknd2d1_hd U665 ( .A(n1139), .B(n1370), .Y(n148) );
  clknd2d1_hd U666 ( .A(n1139), .B(n1363), .Y(n138) );
  nid1_hd U667 ( .A(n9), .Y(n476) );
  clknd2d1_hd U668 ( .A(n1121), .B(n78), .Y(n1122) );
  nid1_hd U669 ( .A(n501), .Y(n500) );
  clknd2d1_hd U670 ( .A(n1126), .B(n1116), .Y(n155) );
  ivd1_hd U671 ( .A(n83), .Y(n84) );
  fad1_hd U672 ( .A(b_m[23]), .B(n596), .CI(n846), .CO(n1065), .S(n1048) );
  ivd1_hd U673 ( .A(n119), .Y(n120) );
  ivd1_hd U674 ( .A(n85), .Y(n86) );
  ivd1_hd U675 ( .A(n84), .Y(n1387) );
  nid1_hd U676 ( .A(n146), .Y(n1) );
  scg12d1_hd U677 ( .A(o_AB_ACK), .B(i_AB_STB), .C(n155), .Y(n146) );
  ivd1_hd U678 ( .A(n1428), .Y(n3) );
  ivd1_hd U679 ( .A(n1428), .Y(n4) );
  nid1_hd U680 ( .A(n1430), .Y(n8) );
  or3d1_hd U681 ( .A(n77), .B(n1129), .C(n1431), .Y(n1428) );
  ivd1_hd U682 ( .A(n1428), .Y(n9) );
  ivd1_hd U683 ( .A(n1428), .Y(n11) );
  ivd1_hd U684 ( .A(n1428), .Y(n12) );
  nid1_hd U685 ( .A(n146), .Y(n13) );
  ivd1_hd U686 ( .A(n1048), .Y(n26) );
  ivd1_hd U687 ( .A(intadd_23_SUM_17_), .Y(n63) );
  ivd1_hd U688 ( .A(intadd_23_SUM_16_), .Y(n65) );
  ivd1_hd U689 ( .A(intadd_23_SUM_15_), .Y(n57) );
  ad2d1_hd U690 ( .A(n829), .B(n811), .Y(n1066) );
  ivd1_hd U691 ( .A(a_m[20]), .Y(n114) );
  ivd1_hd U692 ( .A(b_m[9]), .Y(n540) );
  ivd1_hd U693 ( .A(b_m[11]), .Y(n550) );
  fad1_hd U694 ( .A(n1007), .B(n1006), .CI(n1005), .CO(n1008), .S(n998) );
  fad1_hd U695 ( .A(n949), .B(n948), .CI(n947), .CO(n950), .S(n939) );
  fad1_hd U696 ( .A(n981), .B(n980), .CI(n979), .CO(n982), .S(n971) );
  xo2d1_hd U697 ( .A(a_m[14]), .B(n978), .Y(intadd_28_B_8_) );
  xo2d1_hd U698 ( .A(n472), .B(n824), .Y(intadd_21_A_19_) );
  ivd1_hd U699 ( .A(n26), .Y(n27) );
  xo2d1_hd U700 ( .A(n472), .B(n805), .Y(intadd_21_A_18_) );
  xo2d1_hd U701 ( .A(n470), .B(n845), .Y(intadd_22_B_17_) );
  xo2d1_hd U702 ( .A(n474), .B(n797), .Y(intadd_21_A_17_) );
  ivd1_hd U703 ( .A(n1039), .Y(n67) );
  ivd1_hd U704 ( .A(n1039), .Y(n68) );
  xo2d1_hd U705 ( .A(n475), .B(n769), .Y(intadd_21_A_15_) );
  ivd1_hd U706 ( .A(n63), .Y(n64) );
  ao22d1_hd U707 ( .A(n594), .B(n823), .C(n600), .D(n822), .Y(n846) );
  ivd1_hd U708 ( .A(n65), .Y(n66) );
  xo2d1_hd U709 ( .A(n83), .B(n869), .Y(intadd_26_A_10_) );
  ivd1_hd U710 ( .A(n57), .Y(n58) );
  xo2d1_hd U711 ( .A(n474), .B(n751), .Y(intadd_21_B_12_) );
  ivd1_hd U712 ( .A(intadd_23_SUM_14_), .Y(n59) );
  ivd1_hd U713 ( .A(intadd_23_SUM_13_), .Y(n55) );
  ivd1_hd U714 ( .A(intadd_23_SUM_12_), .Y(n51) );
  xo2d1_hd U715 ( .A(n467), .B(n820), .Y(intadd_24_B_9_) );
  xo2d1_hd U716 ( .A(n91), .B(n884), .Y(intadd_25_A_8_) );
  ivd1_hd U717 ( .A(intadd_23_SUM_11_), .Y(n53) );
  xo2d1_hd U718 ( .A(n85), .B(n807), .Y(intadd_26_A_6_) );
  xo2d1_hd U719 ( .A(n85), .B(n799), .Y(intadd_26_A_5_) );
  xo2d1_hd U720 ( .A(n91), .B(n840), .Y(intadd_25_A_5_) );
  xo2d1_hd U721 ( .A(n85), .B(n793), .Y(intadd_26_B_4_) );
  xo2d1_hd U722 ( .A(DP_OP_116J2_127_7148_n3), .B(n1364), .Y(n1118) );
  xo2d1_hd U723 ( .A(n460), .B(n827), .Y(intadd_25_A_4_) );
  xo2d1_hd U724 ( .A(n463), .B(n771), .Y(intadd_26_A_3_) );
  xo2d1_hd U725 ( .A(n471), .B(n683), .Y(intadd_22_B_2_) );
  or2d1_hd U726 ( .A(n756), .B(n757), .Y(n1003) );
  or2d1_hd U727 ( .A(n829), .B(n828), .Y(n1049) );
  or2d1_hd U728 ( .A(n775), .B(n788), .Y(n1029) );
  or2d1_hd U729 ( .A(n811), .B(n830), .Y(n1050) );
  nid1_hd U730 ( .A(n461), .Y(n464) );
  oa22d1_hd U731 ( .A(n114), .B(a_m[21]), .C(n1411), .D(n122), .Y(n811) );
  ivd1_hd U732 ( .A(n86), .Y(n1382) );
  ivd1_hd U733 ( .A(a_m[20]), .Y(n119) );
  ivd1_hd U734 ( .A(a_m[14]), .Y(n85) );
  ivd1_hd U735 ( .A(b_m[13]), .Y(n559) );
  ivd1_hd U736 ( .A(b_m[10]), .Y(n544) );
  ivd1_hd U737 ( .A(b_m[16]), .Y(n572) );
  ivd1_hd U738 ( .A(b_m[15]), .Y(n568) );
  ivd1_hd U739 ( .A(b_m[19]), .Y(n585) );
  xo2d1_hd U740 ( .A(n1078), .B(n1077), .Y(n1079) );
  ivd1_hd U741 ( .A(intadd_36_n1), .Y(intadd_20_B_27_) );
  ivd1_hd U742 ( .A(n998), .Y(intadd_20_A_27_) );
  xo2d1_hd U743 ( .A(n462), .B(n990), .Y(intadd_36_B_2_) );
  xo2d1_hd U744 ( .A(n121), .B(n1038), .Y(intadd_33_B_2_) );
  xo2d1_hd U745 ( .A(n1404), .B(n850), .Y(intadd_21_B_20_) );
  xo2d1_hd U746 ( .A(n468), .B(n959), .Y(intadd_37_B_2_) );
  xo2d1_hd U747 ( .A(n1377), .B(n1015), .Y(intadd_35_B_2_) );
  xo2d1_hd U748 ( .A(n610), .B(n1057), .Y(n1062) );
  xo2d1_hd U749 ( .A(n607), .B(n929), .Y(intadd_39_B_2_) );
  xo2d1_hd U750 ( .A(n470), .B(n881), .Y(n894) );
  xo2d1_hd U751 ( .A(n1024), .B(n459), .Y(n1031) );
  xo2d1_hd U752 ( .A(n970), .B(n466), .Y(n979) );
  xo2d1_hd U753 ( .A(n1044), .B(n115), .Y(n1052) );
  xo2d1_hd U754 ( .A(n997), .B(n462), .Y(n1005) );
  xo2d1_hd U755 ( .A(n84), .B(n946), .Y(intadd_27_B_10_) );
  xo2d1_hd U756 ( .A(n114), .B(n1030), .Y(intadd_30_B_5_) );
  xo2d1_hd U757 ( .A(n82), .B(n867), .Y(intadd_20_A_16_) );
  xo2d1_hd U758 ( .A(n607), .B(n921), .Y(intadd_24_B_16_) );
  xo2d1_hd U759 ( .A(n92), .B(n1004), .Y(intadd_31_B_4_) );
  xo2d1_hd U760 ( .A(n611), .B(n1051), .Y(intadd_34_B_2_) );
  xo2d1_hd U761 ( .A(a_m[5]), .B(n911), .Y(n914) );
  xo2d1_hd U762 ( .A(n938), .B(n608), .Y(n947) );
  xo2d1_hd U763 ( .A(n854), .B(n473), .Y(intadd_21_A_21_) );
  xo2d1_hd U764 ( .A(n468), .B(n930), .Y(n949) );
  xo2d1_hd U765 ( .A(n462), .B(n960), .Y(n981) );
  xo2d1_hd U766 ( .A(n610), .B(n1040), .Y(n1053) );
  xo2d1_hd U767 ( .A(n1377), .B(n991), .Y(n1007) );
  xo2d1_hd U768 ( .A(a_m[8]), .B(n912), .Y(n913) );
  xo2d1_hd U769 ( .A(n1398), .B(n865), .Y(intadd_22_B_18_) );
  xo2d1_hd U770 ( .A(n113), .B(n1016), .Y(n1032) );
  xo2d1_hd U771 ( .A(n458), .B(n987), .Y(intadd_29_B_7_) );
  xo2d1_hd U772 ( .A(n115), .B(n1012), .Y(intadd_30_B_3_) );
  xo2d1_hd U773 ( .A(n465), .B(n926), .Y(intadd_25_B_11_) );
  xo2d1_hd U774 ( .A(n612), .B(n1036), .Y(intadd_34_CI) );
  xo2d1_hd U775 ( .A(a_m[14]), .B(n956), .Y(intadd_28_B_6_) );
  xo2d1_hd U776 ( .A(n606), .B(n878), .Y(n895) );
  xo2d1_hd U777 ( .A(n470), .B(n837), .Y(intadd_22_B_16_) );
  xo2d1_hd U778 ( .A(n472), .B(n796), .Y(intadd_21_B_16_) );
  xo2d1_hd U779 ( .A(n607), .B(n868), .Y(intadd_24_A_13_) );
  xo2d1_hd U780 ( .A(n464), .B(n945), .Y(intadd_37_B_1_) );
  xo2d1_hd U781 ( .A(a_m[23]), .B(n1026), .Y(intadd_33_A_1_) );
  xo2d1_hd U782 ( .A(n114), .B(n1002), .Y(intadd_35_B_1_) );
  xo2d1_hd U783 ( .A(n465), .B(n916), .Y(intadd_39_A_1_) );
  xo2d1_hd U784 ( .A(n458), .B(n976), .Y(intadd_36_B_1_) );
  xo2d1_hd U785 ( .A(n458), .B(n966), .Y(intadd_36_CI) );
  xo2d1_hd U786 ( .A(n602), .B(n855), .Y(intadd_20_A_15_) );
  xo2d1_hd U787 ( .A(a_m[23]), .B(n1020), .Y(intadd_33_CI) );
  xo2d1_hd U788 ( .A(n470), .B(n821), .Y(intadd_22_B_15_) );
  xo2d1_hd U789 ( .A(n113), .B(n993), .Y(intadd_35_B_0_) );
  xo2d1_hd U790 ( .A(n1382), .B(n934), .Y(intadd_37_CI) );
  xo2d1_hd U791 ( .A(n83), .B(n905), .Y(intadd_39_CI) );
  xo2d1_hd U792 ( .A(n1398), .B(n803), .Y(intadd_22_B_14_) );
  xo2d1_hd U793 ( .A(n611), .B(n1011), .Y(n1017) );
  xo2d1_hd U794 ( .A(n86), .B(n925), .Y(intadd_27_B_8_) );
  xo2d1_hd U795 ( .A(n458), .B(n955), .Y(intadd_38_B_2_) );
  xo2d1_hd U796 ( .A(n475), .B(n763), .Y(intadd_21_A_14_) );
  xo2d1_hd U797 ( .A(n83), .B(n883), .Y(n906) );
  xo2d1_hd U798 ( .A(a_m[8]), .B(n838), .Y(intadd_20_A_14_) );
  xo2d1_hd U799 ( .A(a_m[20]), .B(n986), .Y(intadd_31_B_2_) );
  xo2d1_hd U800 ( .A(n611), .B(n999), .Y(intadd_30_A_2_) );
  xo2d1_hd U801 ( .A(n464), .B(n917), .Y(intadd_25_A_10_) );
  xo2d1_hd U802 ( .A(a_m[17]), .B(n944), .Y(intadd_28_B_5_) );
  xo2d1_hd U803 ( .A(n115), .B(n975), .Y(intadd_29_B_6_) );
  xo2d1_hd U804 ( .A(n1398), .B(n795), .Y(intadd_22_B_13_) );
  xo2d1_hd U805 ( .A(n475), .B(n752), .Y(intadd_21_A_13_) );
  xo2d1_hd U806 ( .A(n603), .B(n825), .Y(intadd_20_A_13_) );
  ivd1_hd U807 ( .A(n59), .Y(n60) );
  xo2d1_hd U808 ( .A(n469), .B(n783), .Y(intadd_22_B_12_) );
  xo2d1_hd U809 ( .A(n461), .B(n897), .Y(intadd_39_A_0_) );
  xo2d1_hd U810 ( .A(n611), .B(n992), .Y(intadd_35_A_0_) );
  xo2d1_hd U811 ( .A(n605), .B(n806), .Y(intadd_20_A_12_) );
  xo2d1_hd U812 ( .A(n114), .B(n965), .Y(intadd_36_B_0_) );
  xo2d1_hd U813 ( .A(n1377), .B(n933), .Y(intadd_37_B_0_) );
  xo2d1_hd U814 ( .A(n1387), .B(n864), .Y(intadd_24_B_12_) );
  xo2d1_hd U815 ( .A(n461), .B(n882), .Y(n907) );
  xo2d1_hd U816 ( .A(n92), .B(n924), .Y(intadd_28_B_3_) );
  xo2d1_hd U817 ( .A(n605), .B(n798), .Y(intadd_20_A_11_) );
  xo2d1_hd U818 ( .A(n113), .B(n954), .Y(intadd_29_B_4_) );
  xo2d1_hd U819 ( .A(n475), .B(n738), .Y(intadd_21_B_11_) );
  xo2d1_hd U820 ( .A(n469), .B(n768), .Y(intadd_22_B_11_) );
  xo2d1_hd U821 ( .A(n468), .B(n844), .Y(intadd_24_B_11_) );
  xo2d1_hd U822 ( .A(n611), .B(n985), .Y(intadd_30_CI) );
  xo2d1_hd U823 ( .A(n469), .B(n762), .Y(intadd_22_B_10_) );
  xo2d1_hd U824 ( .A(n1404), .B(n733), .Y(intadd_21_B_10_) );
  xo2d1_hd U825 ( .A(n115), .B(n943), .Y(intadd_38_B_1_) );
  xo2d1_hd U826 ( .A(n465), .B(n836), .Y(intadd_24_B_10_) );
  xo2d1_hd U827 ( .A(n461), .B(n870), .Y(intadd_25_A_7_) );
  xo2d1_hd U828 ( .A(a_m[17]), .B(n920), .Y(intadd_27_B_7_) );
  xo2d1_hd U829 ( .A(a_m[23]), .B(n972), .Y(intadd_31_A_1_) );
  xo2d1_hd U830 ( .A(n605), .B(n784), .Y(intadd_20_A_10_) );
  xo2d1_hd U831 ( .A(n461), .B(n863), .Y(intadd_26_B_9_) );
  xo2d1_hd U832 ( .A(n469), .B(n739), .Y(intadd_22_A_9_) );
  xo2d1_hd U833 ( .A(n609), .B(n964), .Y(intadd_31_CI) );
  xo2d1_hd U834 ( .A(n605), .B(n770), .Y(intadd_20_A_9_) );
  xo2d1_hd U835 ( .A(n1377), .B(n904), .Y(intadd_25_B_9_) );
  xo2d1_hd U836 ( .A(n114), .B(n932), .Y(intadd_38_CI) );
  xo2d1_hd U837 ( .A(n1404), .B(n723), .Y(intadd_21_B_9_) );
  xo2d1_hd U838 ( .A(n1387), .B(n802), .Y(intadd_24_B_8_) );
  xo2d1_hd U839 ( .A(n122), .B(n923), .Y(intadd_32_B_2_) );
  xo2d1_hd U840 ( .A(n81), .B(n734), .Y(intadd_22_A_8_) );
  xo2d1_hd U841 ( .A(n1084), .B(n1433), .Y(N475) );
  xo2d1_hd U842 ( .A(n103), .B(n709), .Y(intadd_21_B_8_) );
  xo2d1_hd U843 ( .A(n603), .B(n764), .Y(intadd_20_A_8_) );
  xo2d1_hd U844 ( .A(n1382), .B(n839), .Y(intadd_26_A_8_) );
  xo2d1_hd U845 ( .A(n611), .B(n953), .Y(n961) );
  xo2d1_hd U846 ( .A(n103), .B(n705), .Y(intadd_21_B_7_) );
  xo2d1_hd U847 ( .A(n81), .B(n724), .Y(intadd_22_A_7_) );
  xo2d1_hd U848 ( .A(n92), .B(n871), .Y(intadd_27_A_4_) );
  xo2d1_hd U849 ( .A(n612), .B(n940), .Y(intadd_29_A_3_) );
  xo2d1_hd U850 ( .A(DP_OP_125J2_130_6300_n2), .B(n1083), .Y(n1084) );
  xo2d1_hd U851 ( .A(n121), .B(n919), .Y(intadd_28_B_2_) );
  xo2d1_hd U852 ( .A(n603), .B(n753), .Y(intadd_20_A_7_) );
  xo2d1_hd U853 ( .A(n1382), .B(n826), .Y(intadd_26_A_7_) );
  xo2d1_hd U854 ( .A(n103), .B(n695), .Y(intadd_21_B_6_) );
  xo2d1_hd U855 ( .A(n81), .B(n710), .Y(intadd_22_A_6_) );
  fad1_hd U856 ( .A(intadd_22_A_2_), .B(intadd_22_B_2_), .CI(intadd_22_n18), 
        .CO(intadd_22_n17), .S(intadd_21_B_5_) );
  xo2d1_hd U857 ( .A(n612), .B(n931), .Y(intadd_38_B_0_) );
  xo2d1_hd U858 ( .A(n120), .B(n903), .Y(intadd_27_B_6_) );
  xo2d1_hd U859 ( .A(n603), .B(n740), .Y(intadd_20_A_6_) );
  xo2d1_hd U860 ( .A(n91), .B(n862), .Y(intadd_25_B_6_) );
  xo2d1_hd U861 ( .A(n81), .B(n706), .Y(intadd_22_A_5_) );
  xo2d1_hd U862 ( .A(n612), .B(n922), .Y(intadd_29_B_1_) );
  xo2d1_hd U863 ( .A(n113), .B(n890), .Y(n899) );
  xo2d1_hd U864 ( .A(n475), .B(n681), .Y(intadd_21_A_5_) );
  xo2d1_hd U865 ( .A(n603), .B(n735), .Y(intadd_20_A_5_) );
  xo2d1_hd U866 ( .A(a_m[20]), .B(n877), .Y(n885) );
  xo2d1_hd U867 ( .A(n467), .B(n761), .Y(intadd_24_B_4_) );
  xo2d1_hd U868 ( .A(n474), .B(n680), .Y(intadd_21_B_4_) );
  xo2d1_hd U869 ( .A(n603), .B(n732), .Y(intadd_20_B_4_) );
  xo2d1_hd U870 ( .A(n618), .B(n918), .Y(intadd_32_A_1_) );
  xo2d1_hd U871 ( .A(n1398), .B(n704), .Y(intadd_22_B_4_) );
  xo2d1_hd U872 ( .A(n467), .B(n750), .Y(intadd_24_B_3_) );
  xo2d1_hd U873 ( .A(n460), .B(n808), .Y(intadd_25_A_3_) );
  xo2d1_hd U874 ( .A(n471), .B(n684), .Y(intadd_22_A_3_) );
  xo2d1_hd U875 ( .A(n618), .B(n902), .Y(intadd_32_CI) );
  xo2d1_hd U876 ( .A(n474), .B(n671), .Y(intadd_21_B_3_) );
  xo2d1_hd U877 ( .A(n604), .B(n711), .Y(intadd_20_A_3_) );
  xo2d1_hd U878 ( .A(n122), .B(n861), .Y(intadd_27_B_3_) );
  xo2d1_hd U879 ( .A(n618), .B(n891), .Y(intadd_28_CI) );
  xo2d1_hd U880 ( .A(n121), .B(n843), .Y(intadd_27_B_2_) );
  xo2d1_hd U881 ( .A(n463), .B(n766), .Y(intadd_26_B_2_) );
  xo2d1_hd U882 ( .A(n604), .B(n708), .Y(intadd_20_B_2_) );
  xo2d1_hd U883 ( .A(n474), .B(n660), .Y(intadd_21_B_2_) );
  xo2d1_hd U884 ( .A(n467), .B(n737), .Y(intadd_24_B_2_) );
  xo2d1_hd U885 ( .A(n460), .B(n801), .Y(intadd_25_B_2_) );
  xo2d1_hd U886 ( .A(n463), .B(n729), .Y(n731) );
  xo2d1_hd U887 ( .A(n460), .B(n785), .Y(intadd_25_A_1_) );
  xo2d1_hd U888 ( .A(n474), .B(n658), .Y(intadd_21_B_1_) );
  xo2d1_hd U889 ( .A(n604), .B(n696), .Y(intadd_20_A_1_) );
  xo2d1_hd U890 ( .A(n468), .B(n725), .Y(intadd_24_A_1_) );
  xo2d1_hd U891 ( .A(n463), .B(n754), .Y(intadd_26_A_1_) );
  xo2d1_hd U892 ( .A(n612), .B(n875), .Y(n889) );
  xo2d1_hd U893 ( .A(n463), .B(n743), .Y(intadd_26_B_0_) );
  xo2d1_hd U894 ( .A(n471), .B(n672), .Y(intadd_22_A_1_) );
  xo2d1_hd U895 ( .A(n467), .B(n715), .Y(intadd_24_B_0_) );
  xo2d1_hd U896 ( .A(n618), .B(n860), .Y(n872) );
  xo2d1_hd U897 ( .A(n91), .B(n774), .Y(intadd_25_B_0_) );
  xo2d1_hd U898 ( .A(a_m[11]), .B(n701), .Y(n702) );
  xo2d1_hd U899 ( .A(n604), .B(n694), .Y(intadd_20_CI) );
  scg6d1_hd U900 ( .A(n1346), .B(n1344), .C(n110), .Y(n1370) );
  xo2d1_hd U901 ( .A(n121), .B(n819), .Y(intadd_27_CI) );
  xo2d1_hd U902 ( .A(n472), .B(n651), .Y(intadd_21_B_0_) );
  xo2d1_hd U903 ( .A(n471), .B(n663), .Y(intadd_22_B_0_) );
  xo2d1_hd U904 ( .A(n460), .B(n758), .Y(n760) );
  xo2d1_hd U905 ( .A(n82), .B(n659), .Y(n661) );
  xo2d1_hd U906 ( .A(n115), .B(n800), .Y(n809) );
  xo2d1_hd U907 ( .A(n607), .B(n682), .Y(n691) );
  xo2d1_hd U908 ( .A(n612), .B(n842), .Y(n857) );
  xo2d1_hd U909 ( .A(n604), .B(n677), .Y(n678) );
  xo2d1_hd U910 ( .A(n613), .B(n832), .Y(n834) );
  xo2d1_hd U911 ( .A(n121), .B(n790), .Y(n791) );
  xo2d1_hd U912 ( .A(n471), .B(n655), .Y(n657) );
  nid1_hd U913 ( .A(n1340), .Y(n1343) );
  nid1_hd U914 ( .A(n994), .Y(n418) );
  nid1_hd U915 ( .A(n406), .Y(n405) );
  xo2d1_hd U916 ( .A(n602), .B(n942), .Y(intadd_29_B_3_) );
  nid1_hd U917 ( .A(n908), .Y(n394) );
  ad2d1_hd U918 ( .A(n1116), .B(n1121), .Y(n1434) );
  nid1_hd U919 ( .A(n109), .Y(n1117) );
  ivd1_hd U920 ( .A(b_m[23]), .Y(n108) );
  ivd1_hd U921 ( .A(b_m[22]), .Y(n601) );
  oa22ad1_hd U922 ( .A(a_m[21]), .B(a_m[22]), .C(a_m[22]), .D(a_m[21]), .Y(
        n830) );
  xo2d1_hd U923 ( .A(a_s), .B(b_s), .Y(N35) );
  xo2d1_hd U924 ( .A(n1387), .B(n794), .Y(intadd_24_B_7_) );
  xo2d1_hd U925 ( .A(n1387), .B(n782), .Y(intadd_24_B_6_) );
  scg2d1_hd U926 ( .A(n376), .B(n1371), .C(b_e[0]), .D(n80), .Y(n327) );
  scg2d1_hd U927 ( .A(b_e[2]), .B(n79), .C(C82_DATA2_2), .D(n376), .Y(n325) );
  xo2d1_hd U928 ( .A(n1387), .B(n767), .Y(intadd_24_B_5_) );
  scg2d1_hd U929 ( .A(b_e[4]), .B(n80), .C(C82_DATA2_4), .D(n376), .Y(n323) );
  scg2d1_hd U930 ( .A(b_e[5]), .B(n79), .C(C82_DATA2_5), .D(n376), .Y(n322) );
  scg2d1_hd U931 ( .A(b_e[6]), .B(n80), .C(C82_DATA2_6), .D(n376), .Y(n321) );
  scg2d1_hd U932 ( .A(b_e[3]), .B(n80), .C(C82_DATA2_3), .D(n1418), .Y(n324)
         );
  scg9d1_hd U933 ( .A(n640), .B(n639), .C(intadd_21_CI), .Y(N179) );
  xo2d1_hd U934 ( .A(n120), .B(n835), .Y(intadd_27_B_1_) );
  scg9d1_hd U935 ( .A(n634), .B(n633), .C(n635), .Y(N178) );
  scg9d1_hd U936 ( .A(n703), .B(n702), .C(n713), .Y(intadd_20_B_1_) );
  nid1_hd U937 ( .A(n200), .Y(n1281) );
  scg8d1_hd U938 ( .A(n1382), .B(n721), .C(n720), .D(n719), .Y(n722) );
  xo2d1_hd U939 ( .A(a_m[14]), .B(n736), .Y(n741) );
  scg8d1_hd U940 ( .A(n91), .B(n748), .C(n747), .D(n746), .Y(n749) );
  xo2d1_hd U941 ( .A(a_m[17]), .B(n765), .Y(n772) );
  scg10d1_hd U942 ( .A(n1180), .B(n1141), .C(z[31]), .D(n453), .Y(n229) );
  or2d1_hd U943 ( .A(n1433), .B(n94), .Y(n1307) );
  scg6d1_hd U944 ( .A(n1415), .B(n1344), .C(n1392), .Y(n1352) );
  xo2d1_hd U945 ( .A(n465), .B(n707), .Y(n712) );
  nid1_hd U946 ( .A(n453), .Y(n452) );
  or2d1_hd U947 ( .A(n1340), .B(n1416), .Y(n1341) );
  xo2d1_hd U948 ( .A(n107), .B(n638), .Y(n639) );
  scg2d1_hd U949 ( .A(z_e[6]), .B(n89), .C(n496), .D(DP_OP_125J2_130_6300_n40), 
        .Y(DP_OP_125J2_130_6300_n30) );
  scg2d1_hd U950 ( .A(z_e[2]), .B(n89), .C(n497), .D(DP_OP_125J2_130_6300_n36), 
        .Y(DP_OP_125J2_130_6300_n26) );
  scg2d1_hd U951 ( .A(z_e[5]), .B(n90), .C(n496), .D(DP_OP_125J2_130_6300_n39), 
        .Y(DP_OP_125J2_130_6300_n29) );
  scg2d1_hd U952 ( .A(n482), .B(b[29]), .C(b_e[6]), .D(n102), .Y(n1213) );
  scg2d1_hd U953 ( .A(z_e[7]), .B(n90), .C(n496), .D(DP_OP_125J2_130_6300_n41), 
        .Y(DP_OP_125J2_130_6300_n31) );
  scg2d1_hd U954 ( .A(z_e[3]), .B(n90), .C(n497), .D(DP_OP_125J2_130_6300_n37), 
        .Y(DP_OP_125J2_130_6300_n27) );
  xo2d1_hd U955 ( .A(n106), .B(n632), .Y(n633) );
  scg2d1_hd U956 ( .A(z_e[4]), .B(n89), .C(n497), .D(DP_OP_125J2_130_6300_n38), 
        .Y(DP_OP_125J2_130_6300_n28) );
  scg2d1_hd U957 ( .A(z_e[1]), .B(n90), .C(n497), .D(DP_OP_125J2_130_6300_n35), 
        .Y(DP_OP_125J2_130_6300_n25) );
  scg2d1_hd U958 ( .A(n483), .B(b[24]), .C(b_e[1]), .D(n101), .Y(n1208) );
  scg2d1_hd U959 ( .A(z_e[8]), .B(n89), .C(n496), .D(DP_OP_125J2_130_6300_n42), 
        .Y(DP_OP_125J2_130_6300_n32) );
  scg2d1_hd U960 ( .A(n483), .B(b[25]), .C(b_e[2]), .D(n101), .Y(n1209) );
  scg2d1_hd U961 ( .A(n483), .B(b[26]), .C(b_e[3]), .D(n102), .Y(n1210) );
  scg2d1_hd U962 ( .A(n483), .B(b[27]), .C(b_e[4]), .D(n102), .Y(n1211) );
  scg2d1_hd U963 ( .A(n483), .B(b[28]), .C(b_e[5]), .D(n101), .Y(n1212) );
  scg2d1_hd U964 ( .A(n483), .B(a[29]), .C(n99), .D(a_e[6]), .Y(C1_Z_6) );
  scg2d1_hd U965 ( .A(n484), .B(a[28]), .C(n100), .D(a_e[5]), .Y(C1_Z_5) );
  scg2d1_hd U966 ( .A(n484), .B(a[24]), .C(n99), .D(a_e[1]), .Y(C1_Z_1) );
  scg2d1_hd U967 ( .A(n484), .B(a[27]), .C(n99), .D(a_e[4]), .Y(C1_Z_4) );
  scg2d1_hd U968 ( .A(n484), .B(a[25]), .C(n99), .D(a_e[2]), .Y(C1_Z_2) );
  scg2d1_hd U969 ( .A(n484), .B(a[26]), .C(n100), .D(a_e[3]), .Y(C1_Z_3) );
  ad2d1_hd U970 ( .A(n100), .B(n614), .Y(n1412) );
  xo2d1_hd U971 ( .A(n459), .B(n1028), .Y(intadd_33_B_1_) );
  nid1_hd U972 ( .A(n1332), .Y(n485) );
  or2d1_hd U973 ( .A(n1108), .B(n649), .Y(n812) );
  or2d1_hd U974 ( .A(n1424), .B(n1188), .Y(n1301) );
  ad2d1_hd U975 ( .A(n1120), .B(n1433), .Y(n1128) );
  nid1_hd U976 ( .A(n381), .Y(n498) );
  xn2d1_hd U977 ( .A(n637), .B(n512), .Y(n841) );
  xo2d1_hd U978 ( .A(n122), .B(n1047), .Y(intadd_34_A_2_) );
  xo2d1_hd U979 ( .A(n86), .B(n1001), .Y(intadd_30_B_2_) );
  scg2d1_hd U980 ( .A(n1427), .B(z_m[0]), .C(round_bit), .D(n379), .Y(n1085)
         );
  xo2d1_hd U981 ( .A(n468), .B(n974), .Y(intadd_31_B_1_) );
  xn2d1_hd U982 ( .A(n502), .B(n630), .Y(n831) );
  nid1_hd U983 ( .A(n851), .Y(n383) );
  nid1_hd U984 ( .A(n13), .Y(n501) );
  or2d1_hd U985 ( .A(state[1]), .B(n621), .Y(n381) );
  ad4d1_hd U986 ( .A(n1091), .B(a_e[0]), .C(a_e[9]), .D(a_e[8]), .Y(n1415) );
  ad4d1_hd U987 ( .A(b_e[8]), .B(b_e[9]), .C(n1106), .D(b_e[0]), .Y(n1346) );
  or4d1_hd U988 ( .A(product[3]), .B(product[10]), .C(product[11]), .D(
        product[6]), .Y(n1294) );
  ivd1_hd U989 ( .A(b_m[1]), .Y(n380) );
  ivd1_hd U990 ( .A(b_m[0]), .Y(n382) );
  or4d1_hd U991 ( .A(n14), .B(b_e[6]), .C(b_e[1]), .D(b_e[3]), .Y(n1093) );
  or4d1_hd U992 ( .A(a_e[5]), .B(a_e[4]), .C(a_e[1]), .D(a_e[3]), .Y(n1090) );
  ad2d1_hd U993 ( .A(o_Z_STB), .B(i_Z_ACK), .Y(n177) );
  ivd1_hd U994 ( .A(b_m[4]), .Y(n517) );
  ivd1_hd U995 ( .A(b_m[3]), .Y(n513) );
  ivd1_hd U996 ( .A(b_m[2]), .Y(n508) );
  ivd1_hd U997 ( .A(z_m[11]), .Y(n18) );
  ivd1_hd U998 ( .A(n18), .Y(n19) );
  ivd1_hd U999 ( .A(z_m[15]), .Y(n20) );
  ivd1_hd U1000 ( .A(n20), .Y(n21) );
  ivd1_hd U1001 ( .A(z_m[19]), .Y(n22) );
  ivd1_hd U1002 ( .A(n22), .Y(n23) );
  ivd1_hd U1003 ( .A(z_m[0]), .Y(n24) );
  ivd1_hd U1004 ( .A(n24), .Y(n25) );
  ivd1_hd U1005 ( .A(intadd_23_SUM_0_), .Y(n28) );
  ivd1_hd U1006 ( .A(n28), .Y(n29) );
  ivd1_hd U1007 ( .A(intadd_23_SUM_2_), .Y(n30) );
  ivd1_hd U1008 ( .A(n30), .Y(n31) );
  ivd1_hd U1009 ( .A(intadd_23_SUM_1_), .Y(n32) );
  ivd1_hd U1010 ( .A(n32), .Y(n33) );
  ivd1_hd U1011 ( .A(intadd_23_SUM_3_), .Y(n34) );
  ivd1_hd U1012 ( .A(n34), .Y(n35) );
  ivd1_hd U1013 ( .A(intadd_23_SUM_4_), .Y(n37) );
  ivd1_hd U1014 ( .A(n37), .Y(n38) );
  ivd1_hd U1015 ( .A(intadd_23_SUM_6_), .Y(n39) );
  ivd1_hd U1016 ( .A(n39), .Y(n40) );
  ivd1_hd U1017 ( .A(intadd_23_SUM_5_), .Y(n41) );
  ivd1_hd U1018 ( .A(n41), .Y(n42) );
  ivd1_hd U1019 ( .A(intadd_23_SUM_7_), .Y(n43) );
  ivd1_hd U1020 ( .A(n43), .Y(n44) );
  ivd1_hd U1021 ( .A(intadd_23_SUM_8_), .Y(n45) );
  ivd1_hd U1022 ( .A(n45), .Y(n46) );
  ivd1_hd U1023 ( .A(intadd_23_SUM_9_), .Y(n47) );
  ivd1_hd U1024 ( .A(n47), .Y(n48) );
  ivd1_hd U1025 ( .A(intadd_23_SUM_10_), .Y(n49) );
  ivd1_hd U1026 ( .A(n49), .Y(n50) );
  ivd1_hd U1027 ( .A(n51), .Y(n52) );
  ivd1_hd U1028 ( .A(n53), .Y(n54) );
  ivd1_hd U1029 ( .A(n55), .Y(n56) );
  ivd1_hd U1030 ( .A(n1352), .Y(n69) );
  ivd1_hd U1031 ( .A(n1352), .Y(n70) );
  ivd1_hd U1032 ( .A(n812), .Y(n71) );
  ivd1_hd U1033 ( .A(n812), .Y(n72) );
  ivd1_hd U1034 ( .A(n841), .Y(n73) );
  ivd1_hd U1035 ( .A(n841), .Y(n74) );
  ivd1_hd U1036 ( .A(n831), .Y(n75) );
  ivd1_hd U1037 ( .A(n831), .Y(n76) );
  ivd1_hd U1038 ( .A(state[1]), .Y(n77) );
  ivd1_hd U1039 ( .A(state[1]), .Y(n78) );
  ivd1_hd U1040 ( .A(n1370), .Y(n79) );
  ivd1_hd U1041 ( .A(n1370), .Y(n80) );
  ivd1_hd U1042 ( .A(a_m[5]), .Y(n81) );
  ivd1_hd U1043 ( .A(n81), .Y(n82) );
  ivd1_hd U1044 ( .A(a_m[11]), .Y(n83) );
  ivd1_hd U1045 ( .A(n123), .Y(n87) );
  ivd1_hd U1046 ( .A(b_m[0]), .Y(n88) );
  ivd1_hd U1047 ( .A(n1128), .Y(n89) );
  ivd1_hd U1048 ( .A(n1128), .Y(n90) );
  ivd1_hd U1049 ( .A(a_m[17]), .Y(n91) );
  ivd1_hd U1050 ( .A(n1271), .Y(n93) );
  ivd1_hd U1051 ( .A(n1271), .Y(n94) );
  ivd1_hd U1052 ( .A(n1281), .Y(n95) );
  ivd1_hd U1053 ( .A(n1281), .Y(n96) );
  ivd1_hd U1054 ( .A(n1307), .Y(n97) );
  ivd1_hd U1055 ( .A(n1307), .Y(n98) );
  ivd1_hd U1056 ( .A(n1356), .Y(n99) );
  ivd1_hd U1057 ( .A(n1356), .Y(n100) );
  ivd1_hd U1058 ( .A(n1416), .Y(n101) );
  ivd1_hd U1059 ( .A(n1416), .Y(n102) );
  ivd1_hd U1060 ( .A(a_m[2]), .Y(n103) );
  ivd1_hd U1061 ( .A(n103), .Y(n106) );
  ivd1_hd U1062 ( .A(n103), .Y(n107) );
  ivd1_hd U1063 ( .A(n108), .Y(n109) );
  ivd1_hd U1064 ( .A(n1343), .Y(n110) );
  ivd1_hd U1065 ( .A(n1343), .Y(n111) );
  ivd1_hd U1066 ( .A(n1343), .Y(n112) );
  ivd1_hd U1067 ( .A(n120), .Y(n113) );
  ivd1_hd U1068 ( .A(a_m[20]), .Y(n115) );
  ivd1_hd U1069 ( .A(n1434), .Y(n116) );
  ivd1_hd U1070 ( .A(n1434), .Y(n117) );
  ivd1_hd U1071 ( .A(n1434), .Y(n118) );
  ivd1_hd U1072 ( .A(n119), .Y(n121) );
  ivd1_hd U1073 ( .A(n119), .Y(n122) );
  ivd1_hd U1074 ( .A(n382), .Y(n123) );
  ivd1_hd U1075 ( .A(n382), .Y(n124) );
  ivd1_hd U1076 ( .A(n382), .Y(n125) );
  ivd1_hd U1077 ( .A(n1117), .Y(n127) );
  ivd1_hd U1078 ( .A(n1117), .Y(n128) );
  ivd1_hd U1079 ( .A(n1341), .Y(n129) );
  ivd1_hd U1080 ( .A(n1341), .Y(n130) );
  ivd1_hd U1081 ( .A(n1341), .Y(n131) );
  ivd1_hd U1082 ( .A(n1341), .Y(n132) );
  ivd1_hd U1083 ( .A(n849), .Y(n133) );
  ivd1_hd U1084 ( .A(n849), .Y(n134) );
  ivd1_hd U1085 ( .A(n849), .Y(n135) );
  ivd1_hd U1086 ( .A(n849), .Y(n136) );
  ivd1_hd U1087 ( .A(n880), .Y(n137) );
  ivd1_hd U1088 ( .A(n880), .Y(n139) );
  ivd1_hd U1089 ( .A(n880), .Y(n140) );
  ivd1_hd U1090 ( .A(n880), .Y(n142) );
  ivd1_hd U1091 ( .A(n928), .Y(n143) );
  ivd1_hd U1092 ( .A(n928), .Y(n144) );
  ivd1_hd U1093 ( .A(n928), .Y(n145) );
  ivd1_hd U1094 ( .A(n928), .Y(n147) );
  ivd1_hd U1095 ( .A(n958), .Y(n149) );
  ivd1_hd U1096 ( .A(n958), .Y(n150) );
  ivd1_hd U1097 ( .A(n958), .Y(n152) );
  ivd1_hd U1098 ( .A(n958), .Y(n153) );
  ivd1_hd U1099 ( .A(n989), .Y(n154) );
  ivd1_hd U1100 ( .A(n989), .Y(n159) );
  ivd1_hd U1101 ( .A(n989), .Y(n162) );
  ivd1_hd U1102 ( .A(n989), .Y(n163) );
  ivd1_hd U1103 ( .A(n1014), .Y(n164) );
  ivd1_hd U1104 ( .A(n1014), .Y(n165) );
  ivd1_hd U1105 ( .A(n1014), .Y(n166) );
  ivd1_hd U1106 ( .A(n1014), .Y(n167) );
  ivd1_hd U1107 ( .A(n786), .Y(n168) );
  ivd1_hd U1108 ( .A(n786), .Y(n169) );
  ivd1_hd U1109 ( .A(n786), .Y(n170) );
  ivd1_hd U1110 ( .A(n786), .Y(n175) );
  ivd1_hd U1111 ( .A(n380), .Y(n176) );
  ivd1_hd U1112 ( .A(n380), .Y(n178) );
  ivd1_hd U1113 ( .A(n380), .Y(n180) );
  ivd1_hd U1114 ( .A(n380), .Y(n181) );
  ivd1_hd U1115 ( .A(n1049), .Y(n182) );
  ivd1_hd U1116 ( .A(n1049), .Y(n183) );
  ivd1_hd U1117 ( .A(n1049), .Y(n184) );
  ivd1_hd U1118 ( .A(n1049), .Y(n185) );
  ivd1_hd U1119 ( .A(n1301), .Y(n186) );
  ivd1_hd U1120 ( .A(n1301), .Y(n187) );
  ivd1_hd U1121 ( .A(n1301), .Y(n188) );
  ivd1_hd U1122 ( .A(n1301), .Y(n189) );
  nid1_hd U1123 ( .A(z_m[7]), .Y(n190) );
  nid1_hd U1124 ( .A(z_m[3]), .Y(n191) );
  ivd1_hd U1125 ( .A(n1231), .Y(n192) );
  ivd1_hd U1126 ( .A(n1204), .Y(n193) );
  nid1_hd U1127 ( .A(n1176), .Y(n194) );
  scg10d1_hd U1128 ( .A(n1144), .B(n1143), .C(n1178), .D(n1148), .Y(n1176) );
  ivd1_hd U1129 ( .A(n1355), .Y(n195) );
  scg2d1_hd U1130 ( .A(a_e[2]), .B(n70), .C(C81_DATA2_2), .D(n195), .Y(n316)
         );
  scg2d1_hd U1131 ( .A(a_e[3]), .B(n69), .C(C81_DATA2_3), .D(n1358), .Y(n315)
         );
  scg2d1_hd U1132 ( .A(a_e[4]), .B(n70), .C(C81_DATA2_4), .D(n1358), .Y(n314)
         );
  scg2d1_hd U1133 ( .A(a_e[5]), .B(n69), .C(C81_DATA2_5), .D(n1358), .Y(n313)
         );
  scg2d1_hd U1134 ( .A(a_e[6]), .B(n70), .C(C81_DATA2_6), .D(n1358), .Y(n312)
         );
  ivd1_hd U1135 ( .A(b_m[1]), .Y(n197) );
  ivd1_hd U1136 ( .A(n176), .Y(n1339) );
  nid1_hd U1137 ( .A(n97), .Y(n1305) );
  ivd1_hd U1138 ( .A(n1305), .Y(n198) );
  ivd1_hd U1139 ( .A(n1305), .Y(n199) );
  or2d1_hd U1140 ( .A(n1272), .B(n93), .Y(n1312) );
  ivd1_hd U1141 ( .A(n1312), .Y(n200) );
  ivd1_hd U1142 ( .A(n1312), .Y(n201) );
  nid1_hd U1143 ( .A(n1392), .Y(n1409) );
  ivd1_hd U1144 ( .A(n1409), .Y(n202) );
  ivd1_hd U1145 ( .A(n1409), .Y(n203) );
  ivd1_hd U1146 ( .A(n1409), .Y(n204) );
  ivd1_hd U1147 ( .A(n1409), .Y(n205) );
  scg2d1_hd U1148 ( .A(n484), .B(a[0]), .C(n204), .D(a_m[0]), .Y(n349) );
  ivd1_hd U1149 ( .A(n1182), .Y(n206) );
  ivd1_hd U1150 ( .A(n1182), .Y(n207) );
  ivd1_hd U1151 ( .A(n1182), .Y(n208) );
  ivd1_hd U1152 ( .A(n1182), .Y(n209) );
  scg2d1_hd U1153 ( .A(n25), .B(n207), .C(n449), .D(z[0]), .Y(n260) );
  scg2d1_hd U1154 ( .A(z_m[1]), .B(n206), .C(n447), .D(z[1]), .Y(n259) );
  scg2d1_hd U1155 ( .A(z_m[2]), .B(n209), .C(n447), .D(z[2]), .Y(n258) );
  scg2d1_hd U1156 ( .A(n191), .B(n208), .C(n447), .D(z[3]), .Y(n257) );
  scg2d1_hd U1157 ( .A(z_m[4]), .B(n207), .C(n447), .D(z[4]), .Y(n256) );
  scg2d1_hd U1158 ( .A(z_m[5]), .B(n206), .C(n447), .D(z[5]), .Y(n255) );
  scg2d1_hd U1159 ( .A(z_m[6]), .B(n209), .C(n447), .D(z[6]), .Y(n254) );
  scg2d1_hd U1160 ( .A(n190), .B(n208), .C(n448), .D(z[7]), .Y(n253) );
  scg2d1_hd U1161 ( .A(z_m[8]), .B(n207), .C(n448), .D(z[8]), .Y(n252) );
  scg2d1_hd U1162 ( .A(z_m[9]), .B(n206), .C(n448), .D(z[9]), .Y(n251) );
  scg2d1_hd U1163 ( .A(z_m[10]), .B(n209), .C(n448), .D(z[10]), .Y(n250) );
  scg2d1_hd U1164 ( .A(z_m[11]), .B(n208), .C(n448), .D(z[11]), .Y(n249) );
  scg2d1_hd U1165 ( .A(z_m[12]), .B(n207), .C(n448), .D(z[12]), .Y(n248) );
  scg2d1_hd U1166 ( .A(n192), .B(n206), .C(n449), .D(z[13]), .Y(n247) );
  scg2d1_hd U1167 ( .A(z_m[14]), .B(n209), .C(n449), .D(z[14]), .Y(n246) );
  scg2d1_hd U1168 ( .A(z_m[15]), .B(n208), .C(n449), .D(z[15]), .Y(n245) );
  scg2d1_hd U1169 ( .A(z_m[16]), .B(n207), .C(n449), .D(z[16]), .Y(n244) );
  scg2d1_hd U1170 ( .A(n193), .B(n206), .C(n449), .D(z[17]), .Y(n243) );
  scg2d1_hd U1171 ( .A(z_m[18]), .B(n209), .C(n450), .D(z[18]), .Y(n242) );
  scg2d1_hd U1172 ( .A(z_m[19]), .B(n208), .C(n450), .D(z[19]), .Y(n241) );
  scg2d1_hd U1173 ( .A(z_m[20]), .B(n207), .C(n450), .D(z[20]), .Y(n240) );
  scg2d1_hd U1174 ( .A(z_m[21]), .B(n206), .C(n450), .D(z[21]), .Y(n239) );
  ivd1_hd U1175 ( .A(n629), .Y(n210) );
  ivd1_hd U1176 ( .A(n629), .Y(n211) );
  ivd1_hd U1177 ( .A(n629), .Y(n212) );
  ivd1_hd U1178 ( .A(n629), .Y(n213) );
  ivd1_hd U1179 ( .A(n673), .Y(n214) );
  ivd1_hd U1180 ( .A(n673), .Y(n215) );
  ivd1_hd U1181 ( .A(n673), .Y(n216) );
  ivd1_hd U1182 ( .A(n673), .Y(n217) );
  ivd1_hd U1183 ( .A(n697), .Y(n218) );
  ivd1_hd U1184 ( .A(n697), .Y(n219) );
  ivd1_hd U1185 ( .A(n697), .Y(n220) );
  ivd1_hd U1186 ( .A(n697), .Y(n221) );
  ivd1_hd U1187 ( .A(n1412), .Y(n222) );
  ivd1_hd U1188 ( .A(n1412), .Y(n223) );
  ivd1_hd U1189 ( .A(n1412), .Y(n224) );
  ivd1_hd U1190 ( .A(n1412), .Y(n225) );
  ivd1_hd U1191 ( .A(n977), .Y(n226) );
  ivd1_hd U1192 ( .A(n977), .Y(n227) );
  ivd1_hd U1193 ( .A(n977), .Y(n228) );
  ivd1_hd U1194 ( .A(n977), .Y(n359) );
  or2d1_hd U1195 ( .A(n642), .B(n643), .Y(n866) );
  ivd1_hd U1196 ( .A(n866), .Y(n360) );
  ivd1_hd U1197 ( .A(n866), .Y(n361) );
  ivd1_hd U1198 ( .A(n866), .Y(n362) );
  ivd1_hd U1199 ( .A(n866), .Y(n363) );
  ivd1_hd U1200 ( .A(n1003), .Y(n364) );
  ivd1_hd U1201 ( .A(n1003), .Y(n365) );
  ivd1_hd U1202 ( .A(n1003), .Y(n366) );
  ivd1_hd U1203 ( .A(n1003), .Y(n367) );
  ivd1_hd U1204 ( .A(n1029), .Y(n368) );
  ivd1_hd U1205 ( .A(n1029), .Y(n369) );
  ivd1_hd U1206 ( .A(n1029), .Y(n370) );
  ivd1_hd U1207 ( .A(n1029), .Y(n371) );
  ivd1_hd U1208 ( .A(n1050), .Y(n372) );
  ivd1_hd U1209 ( .A(n1050), .Y(n373) );
  ivd1_hd U1210 ( .A(n1050), .Y(n374) );
  ivd1_hd U1211 ( .A(n1050), .Y(n375) );
  nid1_hd U1212 ( .A(n1418), .Y(n376) );
  nid1_hd U1213 ( .A(n1340), .Y(n377) );
  scg2d1_hd U1214 ( .A(n482), .B(b[0]), .C(b_m[0]), .D(n1340), .Y(n308) );
  or2d1_hd U1215 ( .A(n77), .B(n621), .Y(n1433) );
  ivd1_hd U1216 ( .A(n1433), .Y(n378) );
  ivd1_hd U1217 ( .A(n1433), .Y(n379) );
  ao21d1_hd U1218 ( .A(n128), .B(n101), .C(n482), .Y(n1340) );
  ivd1_hd U1219 ( .A(n116), .Y(n1332) );
  oa211d1_hd U1220 ( .A(n1426), .B(n1425), .C(n1424), .D(n499), .Y(n1430) );
  scg12d1_hd U1221 ( .A(n757), .B(n756), .C(n755), .Y(n1021) );
  nr2bd1_hd U1222 ( .AN(n756), .B(n757), .Y(n1022) );
  scg4d1_hd U1223 ( .A(n590), .B(n182), .C(n581), .D(n439), .E(n372), .F(n589), 
        .G(n446), .H(n64), .Y(n1036) );
  ivd1_hd U1224 ( .A(n616), .Y(n614) );
  ivd1_hd U1225 ( .A(n811), .Y(n828) );
  ivd1_hd U1226 ( .A(n1183), .Y(n453) );
  ivd1_hd U1227 ( .A(n1355), .Y(n1358) );
  ivd1_hd U1228 ( .A(n606), .Y(n602) );
  ivd1_hd U1229 ( .A(n789), .Y(n775) );
  scg12d1_hd U1230 ( .A(n789), .B(n788), .C(n787), .Y(n1041) );
  ivd1_hd U1231 ( .A(n617), .Y(n612) );
  ivd1_hd U1232 ( .A(n617), .Y(n611) );
  ivd1_hd U1233 ( .A(n453), .Y(n450) );
  ivd1_hd U1234 ( .A(n452), .Y(n449) );
  ivd1_hd U1235 ( .A(n452), .Y(n448) );
  ivd1_hd U1236 ( .A(n452), .Y(n447) );
  ivd1_hd U1237 ( .A(n452), .Y(n451) );
  ivd1_hd U1238 ( .A(n1148), .Y(n1179) );
  ivd1_hd U1239 ( .A(n69), .Y(n1363) );
  oa21d1_hd U1240 ( .A(n79), .B(n1416), .C(n118), .Y(n1418) );
  ivd1_hd U1241 ( .A(n1143), .Y(n1139) );
  ivd1_hd U1242 ( .A(n1297), .Y(n1308) );
  ivd1_hd U1243 ( .A(n105), .Y(n1299) );
  ivd1_hd U1244 ( .A(n1227), .Y(n1272) );
  scg17d1_hd U1245 ( .A(n1184), .B(n24), .C(net908), .D(n1227), .Y(n1426) );
  ivd1_hd U1246 ( .A(n498), .Y(n496) );
  ivd1_hd U1247 ( .A(n654), .Y(n643) );
  ivd1_hd U1248 ( .A(n950), .Y(intadd_20_B_22_) );
  ivd1_hd U1249 ( .A(a_m[5]), .Y(n1398) );
  ivd1_hd U1250 ( .A(n982), .Y(intadd_20_B_25_) );
  ivd1_hd U1251 ( .A(intadd_36_SUM_2_), .Y(intadd_20_A_26_) );
  ivd1_hd U1252 ( .A(n1008), .Y(intadd_20_B_28_) );
  ivd1_hd U1253 ( .A(intadd_35_SUM_2_), .Y(intadd_20_A_29_) );
  ivd1_hd U1254 ( .A(intadd_30_n1), .Y(intadd_20_B_32_) );
  ivd1_hd U1255 ( .A(n1045), .Y(intadd_20_A_33_) );
  ivd1_hd U1256 ( .A(n1063), .Y(intadd_20_A_36_) );
  ivd1_hd U1257 ( .A(n617), .Y(n610) );
  ivd1_hd U1258 ( .A(n381), .Y(n491) );
  ivd1_hd U1259 ( .A(n381), .Y(n490) );
  ivd1_hd U1260 ( .A(n498), .Y(n495) );
  ivd1_hd U1261 ( .A(n499), .Y(n494) );
  ivd1_hd U1262 ( .A(n499), .Y(n493) );
  ivd1_hd U1263 ( .A(n499), .Y(n492) );
  ivd1_hd U1264 ( .A(n499), .Y(n488) );
  ivd1_hd U1265 ( .A(n499), .Y(n489) );
  ivd1_hd U1266 ( .A(n1170), .Y(n1177) );
  ao21d1_hd U1267 ( .A(n1139), .B(n1127), .C(n1179), .Y(n1183) );
  nr2d1_hd U1268 ( .A(n1127), .B(n1143), .Y(n1344) );
  nd3d1_hd U1269 ( .A(n1144), .B(n1132), .C(n1130), .Y(n1127) );
  nr2d1_hd U1270 ( .A(n1432), .B(n1123), .Y(n1119) );
  ao21d1_hd U1271 ( .A(n379), .B(n1315), .C(n1295), .Y(n1424) );
  nr2d1_hd U1272 ( .A(n1431), .B(n1120), .Y(n1227) );
  ivd1_hd U1273 ( .A(n498), .Y(n497) );
  nr2d1_hd U1274 ( .A(state[3]), .B(n1431), .Y(n1121) );
  ivd1_hd U1275 ( .A(state[0]), .Y(n1431) );
  ivd1_hd U1276 ( .A(n896), .Y(intadd_20_A_18_) );
  ivd1_hd U1277 ( .A(intadd_24_SUM_16_), .Y(intadd_20_B_19_) );
  ivd1_hd U1278 ( .A(intadd_37_SUM_2_), .Y(intadd_20_A_23_) );
  ivd1_hd U1279 ( .A(intadd_37_n1), .Y(intadd_20_B_24_) );
  ivd1_hd U1280 ( .A(n971), .Y(intadd_20_A_24_) );
  ivd1_hd U1281 ( .A(n106), .Y(n1404) );
  ivd1_hd U1282 ( .A(n728), .Y(n716) );
  ivd1_hd U1283 ( .A(n600), .Y(n597) );
  ivd1_hd U1284 ( .A(n1033), .Y(intadd_20_B_31_) );
  ivd1_hd U1285 ( .A(intadd_30_SUM_5_), .Y(intadd_20_A_31_) );
  ivd1_hd U1286 ( .A(n616), .Y(n613) );
  fad1_hd U1287 ( .A(n1053), .B(intadd_34_SUM_1_), .CI(n1052), .CO(n1054), .S(
        n1045) );
  ivd1_hd U1288 ( .A(a_m[18]), .Y(n1376) );
  ivd1_hd U1289 ( .A(intadd_34_n1), .Y(intadd_20_B_35_) );
  ivd1_hd U1290 ( .A(n584), .Y(n581) );
  ivd1_hd U1291 ( .A(n600), .Y(n598) );
  ivd1_hd U1292 ( .A(n594), .Y(n590) );
  ivd1_hd U1293 ( .A(n1060), .Y(intadd_20_A_35_) );
  scg14d1_hd U1294 ( .A(n589), .B(n1340), .C(n1318), .Y(n288) );
  scg14d1_hd U1295 ( .A(n576), .B(n1340), .C(n1321), .Y(n291) );
  scg14d1_hd U1296 ( .A(n554), .B(n377), .C(n1326), .Y(n296) );
  scg14d1_hd U1297 ( .A(n534), .B(n377), .C(n1330), .Y(n300) );
  scg14d1_hd U1298 ( .A(n525), .B(n377), .C(n1333), .Y(n302) );
  scg14d1_hd U1299 ( .A(n580), .B(n377), .C(n1320), .Y(n290) );
  scg14d1_hd U1300 ( .A(n518), .B(n377), .C(n1334), .Y(n303) );
  scg14d1_hd U1301 ( .A(n563), .B(n377), .C(n1324), .Y(n294) );
  scg17d1_hd U1302 ( .A(z_m[8]), .B(n98), .C(n1252), .D(n1251), .Y(n274) );
  scg17d1_hd U1303 ( .A(z_m[4]), .B(n97), .C(n1270), .D(n1269), .Y(n278) );
  scg17d1_hd U1304 ( .A(z_m[12]), .B(n98), .C(n1235), .D(n1234), .Y(n270) );
  scg17d1_hd U1305 ( .A(z_m[16]), .B(n97), .C(n1216), .D(n1215), .Y(n266) );
  oa21d1_hd U1306 ( .A(z_e[7]), .B(z_e[8]), .C(n1142), .Y(n1178) );
  ivd1_hd U1307 ( .A(z_e[9]), .Y(n1142) );
  scg17d1_hd U1308 ( .A(z_m[20]), .B(n98), .C(n1190), .D(n1189), .Y(n262) );
  ivd1_hd U1309 ( .A(n1126), .Y(n1123) );
  nr2d1_hd U1310 ( .A(state[3]), .B(state[0]), .Y(n1126) );
  ivd1_hd U1311 ( .A(state[2]), .Y(n1432) );
  ivd1_hd U1312 ( .A(z_m[23]), .Y(n1315) );
  scg12d1_hd U1313 ( .A(n1245), .B(z_m[10]), .C(n1248), .Y(n1237) );
  scg12d1_hd U1314 ( .A(n1263), .B(z_m[6]), .C(n1266), .Y(n1254) );
  scg12d1_hd U1315 ( .A(z_m[1]), .B(z_m[2]), .C(n24), .Y(n1274) );
  ivd1_hd U1316 ( .A(z_m[22]), .Y(n1311) );
  nr2d1_hd U1317 ( .A(state[1]), .B(state[2]), .Y(n1116) );
  fad1_hd U1318 ( .A(n895), .B(n894), .CI(intadd_24_SUM_14_), .CO(n896), .S(
        n893) );
  nr2d1_hd U1319 ( .A(n625), .B(n624), .Y(n634) );
  ivd1_hd U1320 ( .A(a_m[0]), .Y(n1408) );
  ivd1_hd U1321 ( .A(a_m[1]), .Y(n1406) );
  ivd1_hd U1322 ( .A(n608), .Y(n604) );
  ivd1_hd U1323 ( .A(n608), .Y(n603) );
  fad1_hd U1324 ( .A(n915), .B(n914), .CI(n913), .CO(intadd_20_A_19_), .S(
        intadd_20_B_18_) );
  ivd1_hd U1325 ( .A(a_m[4]), .Y(n1400) );
  ivd1_hd U1326 ( .A(a_m[3]), .Y(n1402) );
  ivd1_hd U1327 ( .A(a_m[7]), .Y(n1394) );
  ivd1_hd U1328 ( .A(a_m[6]), .Y(n1396) );
  ivd1_hd U1329 ( .A(n507), .Y(n504) );
  ivd1_hd U1330 ( .A(a_m[9]), .Y(n1391) );
  ivd1_hd U1331 ( .A(a_m[10]), .Y(n1389) );
  ivd1_hd U1332 ( .A(a_m[13]), .Y(n1384) );
  ivd1_hd U1333 ( .A(a_m[12]), .Y(n1386) );
  ivd1_hd U1334 ( .A(a_m[8]), .Y(n608) );
  ivd1_hd U1335 ( .A(a_m[15]), .Y(n1381) );
  ivd1_hd U1336 ( .A(a_m[16]), .Y(n1379) );
  ivd1_hd U1337 ( .A(n539), .Y(n535) );
  ivd1_hd U1338 ( .A(a_m[19]), .Y(n1374) );
  ivd1_hd U1339 ( .A(a_m[21]), .Y(n1411) );
  nr2d1_hd U1340 ( .A(state[2]), .B(n78), .Y(n1089) );
  nr2d1_hd U1341 ( .A(n1129), .B(state[0]), .Y(n1125) );
  nr2d1_hd U1342 ( .A(n36), .B(n1188), .Y(n1295) );
  ivd1_hd U1343 ( .A(n517), .Y(n516) );
  ivd1_hd U1344 ( .A(n529), .Y(n528) );
  ivd1_hd U1345 ( .A(n544), .Y(n543) );
  ivd1_hd U1346 ( .A(n558), .Y(n557) );
  ivd1_hd U1347 ( .A(n567), .Y(n566) );
  ivd1_hd U1348 ( .A(n595), .Y(n593) );
  ivd1_hd U1349 ( .A(n517), .Y(n515) );
  ivd1_hd U1350 ( .A(n529), .Y(n527) );
  nid2_hd U1351 ( .A(n411), .Y(n413) );
  ivd1_hd U1352 ( .A(n544), .Y(n542) );
  ivd1_hd U1353 ( .A(n558), .Y(n556) );
  ivd1_hd U1354 ( .A(n567), .Y(n565) );
  ivd1_hd U1355 ( .A(n539), .Y(n536) );
  nid2_hd U1356 ( .A(n410), .Y(n408) );
  ivd1_hd U1357 ( .A(n508), .Y(n505) );
  ivd1_hd U1358 ( .A(n549), .Y(n545) );
  ivd1_hd U1359 ( .A(n512), .Y(n511) );
  ivd1_hd U1360 ( .A(n517), .Y(n514) );
  ivd1_hd U1361 ( .A(n512), .Y(n509) );
  ivd1_hd U1362 ( .A(n616), .Y(n615) );
  ivd1_hd U1363 ( .A(n507), .Y(n503) );
  ivd1_hd U1364 ( .A(n512), .Y(n510) );
  ivd1_hd U1365 ( .A(n529), .Y(n526) );
  ivd1_hd U1366 ( .A(n595), .Y(n592) );
  ivd1_hd U1367 ( .A(n544), .Y(n541) );
  ivd1_hd U1368 ( .A(n572), .Y(n570) );
  ivd1_hd U1369 ( .A(n539), .Y(n537) );
  ivd1_hd U1370 ( .A(n539), .Y(n538) );
  ivd1_hd U1371 ( .A(n549), .Y(n546) );
  ivd1_hd U1372 ( .A(n549), .Y(n548) );
  ivd1_hd U1373 ( .A(n608), .Y(n605) );
  ivd1_hd U1374 ( .A(n550), .Y(n547) );
  ivd1_hd U1375 ( .A(n558), .Y(n555) );
  ivd1_hd U1376 ( .A(n584), .Y(n582) );
  ivd1_hd U1377 ( .A(n572), .Y(n571) );
  ivd1_hd U1378 ( .A(n567), .Y(n564) );
  ivd1_hd U1379 ( .A(n572), .Y(n569) );
  ivd1_hd U1380 ( .A(n595), .Y(n591) );
  ivd1_hd U1381 ( .A(n584), .Y(n583) );
  ivd1_hd U1382 ( .A(n600), .Y(n599) );
  ivd1_hd U1383 ( .A(n507), .Y(n506) );
  ivd1_hd U1384 ( .A(a_e[0]), .Y(n1354) );
  nr2d1_hd U1385 ( .A(n1356), .B(n1354), .Y(n1206) );
  ao22d1_hd U1386 ( .A(n497), .B(DP_OP_125J2_130_6300_n34), .C(z_e[0]), .D(n89), .Y(n1429) );
  ivd1_hd U1387 ( .A(n626), .Y(N176) );
  nr2d1_hd U1388 ( .A(n124), .B(n178), .Y(n1108) );
  nr2d1_hd U1389 ( .A(n87), .B(n1339), .Y(n649) );
  oa22d1_hd U1390 ( .A(n472), .B(n1406), .C(a_m[1]), .D(n107), .Y(n622) );
  nr2d1_hd U1391 ( .A(n622), .B(n1408), .Y(n852) );
  oa22d1_hd U1392 ( .A(n87), .B(n849), .C(n197), .D(n629), .Y(n623) );
  ao21d1_hd U1393 ( .A(n71), .B(n388), .C(n623), .Y(n628) );
  nr3d1_hd U1394 ( .A(n628), .B(n626), .C(n473), .Y(n627) );
  ao211d1_hd U1395 ( .A(n628), .B(n473), .C(n634), .D(n627), .Y(N177) );
  nr2d1_hd U1396 ( .A(n125), .B(n1339), .Y(n630) );
  nr2d1_hd U1397 ( .A(a_m[0]), .B(n631), .Y(n851) );
  scg4d1_hd U1398 ( .A(n504), .B(n210), .C(n181), .D(n133), .E(n852), .F(n75), 
        .G(n384), .H(n124), .Y(n632) );
  oa22d1_hd U1399 ( .A(n1402), .B(n107), .C(n473), .D(a_m[3]), .Y(n654) );
  nr2d1_hd U1400 ( .A(n502), .B(n1339), .Y(n636) );
  ao22d1_hd U1401 ( .A(n124), .B(n636), .C(n502), .D(n1339), .Y(n637) );
  scg4d1_hd U1402 ( .A(intadd_23_B_0_), .B(n212), .C(n178), .D(n384), .E(n390), 
        .F(n74), .G(n135), .H(n503), .Y(n638) );
  oa22d1_hd U1403 ( .A(n1402), .B(a_m[4]), .C(n1400), .D(a_m[3]), .Y(n653) );
  nr2d1_hd U1404 ( .A(a_m[4]), .B(n82), .Y(n1098) );
  ao21d1_hd U1405 ( .A(a_m[5]), .B(a_m[4]), .C(n1098), .Y(n642) );
  ivd1_hd U1406 ( .A(n642), .Y(n652) );
  nr2d1_hd U1407 ( .A(n643), .B(n652), .Y(n909) );
  ao22d1_hd U1408 ( .A(n180), .B(n360), .C(n395), .D(n71), .Y(n644) );
  oa21d1_hd U1409 ( .A(n88), .B(n880), .C(n644), .Y(n647) );
  nr2d1_hd U1410 ( .A(n471), .B(n647), .Y(n646) );
  nd2bd1_hd U1411 ( .AN(n645), .B(n646), .Y(n656) );
  scg17d1_hd U1412 ( .A(n469), .B(n647), .C(n646), .D(n645), .Y(n648) );
  nr2d1_hd U1413 ( .A(n502), .B(n649), .Y(n650) );
  oa22d1_hd U1414 ( .A(n512), .B(n650), .C(n1339), .D(n507), .Y(intadd_23_CI)
         );
  scg4d1_hd U1415 ( .A(n514), .B(n211), .C(n506), .D(n385), .E(n387), .F(n29), 
        .G(intadd_23_B_0_), .H(n134), .Y(n651) );
  ivd1_hd U1416 ( .A(intadd_21_SUM_0_), .Y(N180) );
  nr3d1_hd U1417 ( .A(n654), .B(n653), .C(n652), .Y(n908) );
  scg4d1_hd U1418 ( .A(n504), .B(n361), .C(n181), .D(n137), .E(n393), .F(n123), 
        .G(n395), .H(n75), .Y(n655) );
  nr2d1_hd U1419 ( .A(n657), .B(n656), .Y(n662) );
  scg6d1_hd U1420 ( .A(n657), .B(n656), .C(n662), .Y(intadd_21_A_1_) );
  scg4d1_hd U1421 ( .A(n516), .B(n136), .C(n510), .D(n386), .E(n387), .F(
        intadd_23_SUM_1_), .G(n213), .H(intadd_23_B_2_), .Y(n658) );
  ivd1_hd U1422 ( .A(intadd_21_SUM_1_), .Y(N181) );
  scg4d1_hd U1423 ( .A(n509), .B(n362), .C(n178), .D(n392), .E(n139), .F(n506), 
        .G(n73), .H(n395), .Y(n659) );
  oa22d1_hd U1424 ( .A(n470), .B(n1396), .C(a_m[6]), .D(n82), .Y(n664) );
  ivd1_hd U1425 ( .A(n664), .Y(n676) );
  xo3d1_hd U1426 ( .A(n662), .B(n661), .C(n666), .Y(intadd_21_A_2_) );
  scg4d1_hd U1427 ( .A(n516), .B(n383), .C(n519), .D(n133), .E(n522), .F(n210), 
        .G(n388), .H(intadd_23_SUM_2_), .Y(n660) );
  ivd1_hd U1428 ( .A(intadd_21_SUM_2_), .Y(N182) );
  scg16d1_hd U1429 ( .A(n666), .B(n662), .C(n661), .Y(intadd_22_A_0_) );
  scg4d1_hd U1430 ( .A(n516), .B(n363), .C(n505), .D(n392), .E(n140), .F(n511), 
        .G(n396), .H(n29), .Y(n663) );
  oa22d1_hd U1431 ( .A(n606), .B(n1394), .C(a_m[7]), .D(n602), .Y(n674) );
  nr2d1_hd U1432 ( .A(n664), .B(n674), .Y(n936) );
  nr2d1_hd U1433 ( .A(a_m[7]), .B(a_m[6]), .Y(n1097) );
  ao21d1_hd U1434 ( .A(a_m[6]), .B(a_m[7]), .C(n1097), .Y(n675) );
  oa22d1_hd U1435 ( .A(n87), .B(n928), .C(n1339), .D(n673), .Y(n665) );
  ao21d1_hd U1436 ( .A(n72), .B(n404), .C(n665), .Y(n669) );
  nr2d1_hd U1437 ( .A(n667), .B(n668), .Y(n679) );
  oa211d1_hd U1438 ( .A(n602), .B(n669), .C(n668), .D(n667), .Y(n670) );
  nd2bd1_hd U1439 ( .AN(n679), .B(n670), .Y(intadd_22_CI) );
  scg4d1_hd U1440 ( .A(n526), .B(n211), .C(n519), .D(n386), .E(n387), .F(
        intadd_23_SUM_3_), .G(n523), .H(n134), .Y(n671) );
  ivd1_hd U1441 ( .A(intadd_21_SUM_3_), .Y(N183) );
  scg4d1_hd U1442 ( .A(n516), .B(n142), .C(n510), .D(n391), .E(n521), .F(n360), 
        .G(n396), .H(n33), .Y(n672) );
  nr3d1_hd U1443 ( .A(n676), .B(n675), .C(n674), .Y(n935) );
  scg4d1_hd U1444 ( .A(n504), .B(n214), .C(n176), .D(n143), .E(n76), .F(n405), 
        .G(n125), .H(n400), .Y(n677) );
  oa21d1_hd U1445 ( .A(n679), .B(n678), .C(n692), .Y(intadd_22_B_1_) );
  scg4d1_hd U1446 ( .A(n528), .B(n135), .C(n523), .D(n386), .E(n387), .F(
        intadd_23_SUM_4_), .G(n212), .H(intadd_23_B_5_), .Y(n680) );
  ivd1_hd U1447 ( .A(intadd_21_SUM_4_), .Y(N184) );
  scg4d1_hd U1448 ( .A(n528), .B(n386), .C(n532), .D(n136), .E(n537), .F(n213), 
        .G(n389), .H(intadd_23_SUM_5_), .Y(n681) );
  scg4d1_hd U1449 ( .A(n509), .B(n215), .C(n181), .D(n401), .E(n144), .F(n505), 
        .G(n404), .H(n74), .Y(n682) );
  xo3d1_hd U1450 ( .A(n691), .B(n693), .C(n692), .Y(intadd_22_A_2_) );
  scg4d1_hd U1451 ( .A(n515), .B(n392), .C(n519), .D(n137), .E(n524), .F(n361), 
        .G(n397), .H(n31), .Y(n683) );
  ivd1_hd U1452 ( .A(intadd_21_SUM_5_), .Y(N185) );
  scg4d1_hd U1453 ( .A(n528), .B(n362), .C(n520), .D(n391), .E(n139), .F(n525), 
        .G(n396), .H(n35), .Y(n684) );
  oa22d1_hd U1454 ( .A(n466), .B(n1389), .C(a_m[10]), .D(n84), .Y(n698) );
  ivd1_hd U1455 ( .A(n700), .Y(n685) );
  nr2d1_hd U1456 ( .A(n698), .B(n685), .Y(n968) );
  nr2d1_hd U1457 ( .A(a_m[10]), .B(a_m[9]), .Y(n1096) );
  ao21d1_hd U1458 ( .A(a_m[9]), .B(a_m[10]), .C(n1096), .Y(n699) );
  oa22d1_hd U1459 ( .A(n88), .B(n958), .C(n197), .D(n697), .Y(n686) );
  ao21d1_hd U1460 ( .A(n71), .B(n411), .C(n686), .Y(n690) );
  nr2d1_hd U1461 ( .A(n688), .B(n687), .Y(n703) );
  nr3d1_hd U1462 ( .A(n690), .B(n693), .C(n466), .Y(n689) );
  ao211d1_hd U1463 ( .A(n690), .B(n466), .C(n703), .D(n689), .Y(intadd_20_A_0_) );
  ao21d1_hd U1464 ( .A(n693), .B(n692), .C(n691), .Y(intadd_20_B_0_) );
  scg4d1_hd U1465 ( .A(n515), .B(n216), .C(n505), .D(n402), .E(n405), .F(
        intadd_23_SUM_0_), .G(n145), .H(intadd_23_B_0_), .Y(n694) );
  ivd1_hd U1466 ( .A(intadd_20_SUM_0_), .Y(intadd_22_B_3_) );
  scg4d1_hd U1467 ( .A(n536), .B(n133), .C(n541), .D(n210), .E(n851), .F(n534), 
        .G(n389), .H(n40), .Y(n695) );
  ivd1_hd U1468 ( .A(intadd_21_SUM_6_), .Y(N186) );
  scg4d1_hd U1469 ( .A(n515), .B(n147), .C(n511), .D(n402), .E(n406), .F(n33), 
        .G(n519), .H(n217), .Y(n696) );
  scg4d1_hd U1470 ( .A(n504), .B(n218), .C(n180), .D(n149), .E(n409), .F(n124), 
        .G(n75), .H(n411), .Y(n701) );
  ivd1_hd U1471 ( .A(intadd_20_SUM_1_), .Y(intadd_22_A_4_) );
  scg4d1_hd U1472 ( .A(n528), .B(n140), .C(n523), .D(n391), .E(n534), .F(n363), 
        .G(n396), .H(n38), .Y(n704) );
  scg4d1_hd U1473 ( .A(n546), .B(n211), .C(n543), .D(n134), .E(n383), .F(n538), 
        .G(n389), .H(n44), .Y(n705) );
  ivd1_hd U1474 ( .A(intadd_21_SUM_7_), .Y(N187) );
  scg4d1_hd U1475 ( .A(n527), .B(n392), .C(n532), .D(n142), .E(n537), .F(n360), 
        .G(n909), .H(n42), .Y(n706) );
  scg4d1_hd U1476 ( .A(n509), .B(n219), .C(n178), .D(n408), .E(n73), .F(n414), 
        .G(n503), .H(n150), .Y(n707) );
  oa22d1_hd U1477 ( .A(n466), .B(a_m[12]), .C(n1386), .D(n84), .Y(n728) );
  ivd1_hd U1478 ( .A(n714), .Y(n718) );
  xo3d1_hd U1479 ( .A(n712), .B(n718), .C(n713), .Y(intadd_20_A_2_) );
  scg4d1_hd U1480 ( .A(n515), .B(n399), .C(n519), .D(n143), .E(n936), .F(n31), 
        .G(n523), .H(n214), .Y(n708) );
  ivd1_hd U1481 ( .A(intadd_20_SUM_2_), .Y(intadd_22_B_5_) );
  scg4d1_hd U1482 ( .A(intadd_23_B_9_), .B(n212), .C(n543), .D(n385), .E(n387), 
        .F(n46), .G(n545), .H(n135), .Y(n709) );
  ivd1_hd U1483 ( .A(intadd_21_SUM_8_), .Y(N188) );
  scg4d1_hd U1484 ( .A(n536), .B(n137), .C(n543), .D(n361), .E(n534), .F(n393), 
        .G(n909), .H(n40), .Y(n710) );
  scg4d1_hd U1485 ( .A(n527), .B(n215), .C(n519), .D(n402), .E(n936), .F(n35), 
        .G(n144), .H(intadd_23_B_3_), .Y(n711) );
  scg6d1_hd U1486 ( .A(n714), .B(n713), .C(n712), .Y(intadd_24_A_0_) );
  scg4d1_hd U1487 ( .A(n515), .B(n220), .C(n505), .D(n408), .E(n152), .F(n511), 
        .G(n413), .H(n29), .Y(n715) );
  nr2d1_hd U1488 ( .A(a_m[13]), .B(a_m[12]), .Y(n1101) );
  ao21d1_hd U1489 ( .A(a_m[12]), .B(a_m[13]), .C(n1101), .Y(n727) );
  oa22d1_hd U1490 ( .A(n462), .B(n1384), .C(a_m[13]), .D(n86), .Y(n726) );
  nr2d1_hd U1491 ( .A(n716), .B(n726), .Y(n995) );
  ao22d1_hd U1492 ( .A(n176), .B(n226), .C(n72), .D(n420), .Y(n717) );
  oa21d1_hd U1493 ( .A(n88), .B(n989), .C(n717), .Y(n721) );
  nr2d1_hd U1494 ( .A(n461), .B(n721), .Y(n719) );
  nr2d1_hd U1495 ( .A(n718), .B(n463), .Y(n720) );
  ivd1_hd U1496 ( .A(intadd_24_SUM_0_), .Y(intadd_20_B_3_) );
  ivd1_hd U1497 ( .A(intadd_20_SUM_3_), .Y(intadd_22_B_6_) );
  scg4d1_hd U1498 ( .A(n553), .B(n136), .C(n555), .D(n213), .E(n383), .F(n548), 
        .G(n389), .H(n48), .Y(n723) );
  ivd1_hd U1499 ( .A(intadd_21_SUM_9_), .Y(N189) );
  scg4d1_hd U1500 ( .A(n546), .B(n362), .C(n543), .D(n139), .E(n393), .F(n538), 
        .G(n397), .H(n44), .Y(n724) );
  scg4d1_hd U1501 ( .A(n515), .B(n153), .C(n511), .D(n407), .E(n518), .F(n221), 
        .G(n413), .H(n33), .Y(n725) );
  nr3d1_hd U1502 ( .A(n728), .B(n727), .C(n726), .Y(n994) );
  scg4d1_hd U1503 ( .A(n506), .B(n227), .C(n180), .D(n154), .E(n417), .F(n123), 
        .G(n76), .H(n420), .Y(n729) );
  nr2d1_hd U1504 ( .A(n731), .B(n730), .Y(n742) );
  scg6d1_hd U1505 ( .A(n731), .B(n730), .C(n742), .Y(intadd_24_B_1_) );
  ivd1_hd U1506 ( .A(intadd_24_SUM_1_), .Y(intadd_20_A_4_) );
  scg4d1_hd U1507 ( .A(n527), .B(n145), .C(n523), .D(n402), .E(n936), .F(n38), 
        .G(n532), .H(n216), .Y(n732) );
  ivd1_hd U1508 ( .A(intadd_20_SUM_4_), .Y(intadd_22_B_7_) );
  scg4d1_hd U1509 ( .A(n554), .B(n386), .C(n557), .D(n133), .E(n561), .F(n210), 
        .G(n389), .H(n50), .Y(n733) );
  ivd1_hd U1510 ( .A(intadd_21_SUM_10_), .Y(N190) );
  scg4d1_hd U1511 ( .A(n554), .B(n363), .C(n542), .D(n391), .E(n140), .F(n548), 
        .G(n397), .H(n46), .Y(n734) );
  scg4d1_hd U1512 ( .A(n527), .B(n399), .C(n532), .D(n147), .E(n936), .F(n42), 
        .G(n535), .H(n217), .Y(n735) );
  scg4d1_hd U1513 ( .A(n509), .B(n228), .C(n181), .D(n416), .E(n73), .F(n422), 
        .G(n503), .H(n159), .Y(n736) );
  ao22d1_hd U1514 ( .A(n86), .B(n1381), .C(a_m[15]), .D(n462), .Y(n757) );
  nr2d1_hd U1515 ( .A(n87), .B(n757), .Y(n745) );
  xn3d1_hd U1516 ( .A(n741), .B(n745), .C(n742), .Y(intadd_24_A_2_) );
  scg4d1_hd U1517 ( .A(n516), .B(n408), .C(n520), .D(n149), .E(n524), .F(n218), 
        .G(n413), .H(n31), .Y(n737) );
  ivd1_hd U1518 ( .A(intadd_24_SUM_2_), .Y(intadd_20_B_5_) );
  ivd1_hd U1519 ( .A(intadd_20_SUM_5_), .Y(intadd_22_B_8_) );
  scg4d1_hd U1520 ( .A(n564), .B(n211), .C(n557), .D(n385), .E(n390), .F(n54), 
        .G(n560), .H(n134), .Y(n738) );
  ivd1_hd U1521 ( .A(intadd_21_SUM_11_), .Y(N191) );
  scg4d1_hd U1522 ( .A(n554), .B(n142), .C(n557), .D(n360), .E(n546), .F(n393), 
        .G(n397), .H(n48), .Y(n739) );
  scg4d1_hd U1523 ( .A(n536), .B(n143), .C(n542), .D(n214), .E(n406), .F(
        intadd_23_SUM_6_), .G(n400), .H(n532), .Y(n740) );
  oa21d1_hd U1524 ( .A(n745), .B(n742), .C(n741), .Y(intadd_26_A_0_) );
  scg4d1_hd U1525 ( .A(n516), .B(n359), .C(n505), .D(n416), .E(n162), .F(n511), 
        .G(n421), .H(n29), .Y(n743) );
  nr2d1_hd U1526 ( .A(a_m[16]), .B(a_m[15]), .Y(n1100) );
  ao21d1_hd U1527 ( .A(a_m[15]), .B(a_m[16]), .C(n1100), .Y(n755) );
  ao22d1_hd U1528 ( .A(a_m[17]), .B(a_m[16]), .C(n1379), .D(n459), .Y(n756) );
  ao22d1_hd U1529 ( .A(n176), .B(n364), .C(n72), .D(n428), .Y(n744) );
  oa21d1_hd U1530 ( .A(n88), .B(n1014), .C(n744), .Y(n748) );
  nr2d1_hd U1531 ( .A(n458), .B(n748), .Y(n746) );
  nr2d1_hd U1532 ( .A(n745), .B(n460), .Y(n747) );
  scg4d1_hd U1533 ( .A(n527), .B(n219), .C(n520), .D(n407), .E(n150), .F(n525), 
        .G(n413), .H(n35), .Y(n750) );
  ivd1_hd U1534 ( .A(intadd_24_SUM_3_), .Y(intadd_20_B_6_) );
  ivd1_hd U1535 ( .A(intadd_20_SUM_6_), .Y(intadd_22_B_9_) );
  scg4d1_hd U1536 ( .A(n566), .B(n135), .C(n560), .D(n385), .E(n390), .F(n52), 
        .G(n212), .H(intadd_23_B_13_), .Y(n751) );
  ivd1_hd U1537 ( .A(intadd_21_SUM_12_), .Y(N192) );
  scg4d1_hd U1538 ( .A(n566), .B(n386), .C(n569), .D(n136), .E(n573), .F(n213), 
        .G(n389), .H(n56), .Y(n752) );
  scg4d1_hd U1539 ( .A(n545), .B(n215), .C(n542), .D(n144), .E(n406), .F(n44), 
        .G(n400), .H(n535), .Y(n753) );
  scg4d1_hd U1540 ( .A(b_m[4]), .B(n163), .C(b_m[3]), .D(n415), .E(n518), .F(
        n226), .G(n421), .H(n33), .Y(n754) );
  scg4d1_hd U1541 ( .A(n506), .B(n365), .C(n180), .D(n164), .E(n426), .F(n125), 
        .G(n76), .H(n428), .Y(n758) );
  nr2d1_hd U1542 ( .A(n760), .B(n759), .Y(n773) );
  scg6d1_hd U1543 ( .A(n760), .B(n759), .C(n773), .Y(intadd_26_B_1_) );
  scg4d1_hd U1544 ( .A(n527), .B(n152), .C(n522), .D(n407), .E(n534), .F(n220), 
        .G(n413), .H(n38), .Y(n761) );
  ivd1_hd U1545 ( .A(intadd_24_SUM_4_), .Y(intadd_20_B_7_) );
  ivd1_hd U1546 ( .A(intadd_20_SUM_7_), .Y(intadd_22_A_10_) );
  scg4d1_hd U1547 ( .A(n554), .B(n392), .C(n557), .D(n137), .E(n562), .F(n361), 
        .G(n397), .H(n50), .Y(n762) );
  ivd1_hd U1548 ( .A(intadd_21_SUM_13_), .Y(N193) );
  scg4d1_hd U1549 ( .A(intadd_23_B_15_), .B(n210), .C(n570), .D(n385), .E(n390), .F(n60), .G(n574), .H(n133), .Y(n763) );
  scg4d1_hd U1550 ( .A(n554), .B(n216), .C(n542), .D(n402), .E(n406), .F(n46), 
        .G(n145), .H(n545), .Y(n764) );
  scg4d1_hd U1551 ( .A(n509), .B(n366), .C(n176), .D(n425), .E(n74), .F(n430), 
        .G(n503), .H(n165), .Y(n765) );
  oa22d1_hd U1552 ( .A(n459), .B(n1376), .C(a_m[18]), .D(n92), .Y(n789) );
  xo3d1_hd U1553 ( .A(n773), .B(n772), .C(n777), .Y(intadd_26_A_2_) );
  scg4d1_hd U1554 ( .A(b_m[4]), .B(n416), .C(n520), .D(n154), .E(n524), .F(
        n227), .G(n421), .H(n31), .Y(n766) );
  scg4d1_hd U1555 ( .A(n528), .B(n408), .C(n532), .D(n153), .E(n537), .F(n221), 
        .G(n413), .H(n42), .Y(n767) );
  ivd1_hd U1556 ( .A(intadd_24_SUM_5_), .Y(intadd_20_B_8_) );
  ivd1_hd U1557 ( .A(intadd_20_SUM_8_), .Y(intadd_22_A_11_) );
  scg4d1_hd U1558 ( .A(n566), .B(n362), .C(n556), .D(n391), .E(n139), .F(n563), 
        .G(n396), .H(n54), .Y(n768) );
  ivd1_hd U1559 ( .A(intadd_21_SUM_14_), .Y(N194) );
  scg4d1_hd U1560 ( .A(n579), .B(n134), .C(n574), .D(n385), .E(n390), .F(n58), 
        .G(n211), .H(intadd_23_B_16_), .Y(n769) );
  scg4d1_hd U1561 ( .A(n553), .B(n147), .C(n556), .D(n217), .E(n406), .F(n48), 
        .G(n400), .H(n545), .Y(n770) );
  scg4d1_hd U1562 ( .A(n528), .B(n228), .C(n520), .D(n415), .E(n159), .F(n524), 
        .G(n421), .H(n35), .Y(n771) );
  scg16d1_hd U1563 ( .A(n777), .B(n773), .C(n772), .Y(intadd_25_A_0_) );
  scg4d1_hd U1564 ( .A(b_m[4]), .B(n367), .C(n505), .D(n425), .E(n166), .F(
        b_m[3]), .G(n429), .H(intadd_23_SUM_0_), .Y(n774) );
  oa22d1_hd U1565 ( .A(n113), .B(n1374), .C(a_m[19]), .D(n121), .Y(n787) );
  nr2d1_hd U1566 ( .A(n789), .B(n787), .Y(n1042) );
  oa22d1_hd U1567 ( .A(n1374), .B(n1376), .C(a_m[18]), .D(a_m[19]), .Y(n788)
         );
  oa22d1_hd U1568 ( .A(n87), .B(n1029), .C(n197), .D(n786), .Y(n776) );
  ao21d1_hd U1569 ( .A(n71), .B(n435), .C(n776), .Y(n780) );
  nr2d1_hd U1570 ( .A(n778), .B(n779), .Y(n792) );
  oa211d1_hd U1571 ( .A(n122), .B(n780), .C(n779), .D(n778), .Y(n781) );
  nd2bd1_hd U1572 ( .AN(n792), .B(n781), .Y(intadd_25_CI) );
  scg4d1_hd U1573 ( .A(n536), .B(n149), .C(n542), .D(n218), .E(n534), .F(n409), 
        .G(n412), .H(n40), .Y(n782) );
  ivd1_hd U1574 ( .A(intadd_24_SUM_6_), .Y(intadd_20_B_9_) );
  ivd1_hd U1575 ( .A(intadd_20_SUM_9_), .Y(intadd_22_A_12_) );
  scg4d1_hd U1576 ( .A(n566), .B(n140), .C(n560), .D(n394), .E(n571), .F(n363), 
        .G(n398), .H(n52), .Y(n783) );
  ivd1_hd U1577 ( .A(intadd_21_SUM_15_), .Y(N195) );
  scg4d1_hd U1578 ( .A(n553), .B(n399), .C(n556), .D(n143), .E(n405), .F(n50), 
        .G(n560), .H(n214), .Y(n784) );
  scg4d1_hd U1579 ( .A(n514), .B(n167), .C(n510), .D(n424), .E(b_m[5]), .F(
        n364), .G(n429), .H(intadd_23_SUM_1_), .Y(n785) );
  scg4d1_hd U1580 ( .A(n506), .B(n168), .C(n178), .D(n369), .E(n434), .F(n123), 
        .G(n75), .H(n435), .Y(n790) );
  oa21d1_hd U1581 ( .A(n792), .B(n791), .C(n810), .Y(intadd_25_B_1_) );
  scg4d1_hd U1582 ( .A(b_m[7]), .B(n162), .C(b_m[6]), .D(n415), .E(n533), .F(
        n359), .G(n421), .H(n38), .Y(n793) );
  scg4d1_hd U1583 ( .A(n545), .B(n219), .C(n542), .D(n150), .E(n409), .F(n538), 
        .G(n412), .H(intadd_23_SUM_7_), .Y(n794) );
  ivd1_hd U1584 ( .A(intadd_24_SUM_7_), .Y(intadd_20_B_10_) );
  ivd1_hd U1585 ( .A(intadd_20_SUM_10_), .Y(intadd_22_A_13_) );
  scg4d1_hd U1586 ( .A(n565), .B(n392), .C(n570), .D(n142), .E(n575), .F(n360), 
        .G(n398), .H(n56), .Y(n795) );
  scg4d1_hd U1587 ( .A(n580), .B(n851), .C(n581), .D(n135), .E(n588), .F(n212), 
        .G(n388), .H(n66), .Y(n796) );
  ivd1_hd U1588 ( .A(intadd_21_SUM_16_), .Y(N196) );
  scg4d1_hd U1589 ( .A(n590), .B(n213), .C(n582), .D(n384), .E(n852), .F(n64), 
        .G(n586), .H(n136), .Y(n797) );
  scg4d1_hd U1590 ( .A(n565), .B(n215), .C(n556), .D(n401), .E(n403), .F(n54), 
        .G(n144), .H(intadd_23_B_11_), .Y(n798) );
  scg4d1_hd U1591 ( .A(b_m[7]), .B(n416), .C(n531), .D(n163), .E(n536), .F(
        n226), .G(n421), .H(n42), .Y(n799) );
  scg4d1_hd U1592 ( .A(n510), .B(n169), .C(n181), .D(n433), .E(n73), .F(n436), 
        .G(n504), .H(n370), .Y(n800) );
  xo3d1_hd U1593 ( .A(n814), .B(n809), .C(n810), .Y(intadd_25_A_2_) );
  scg4d1_hd U1594 ( .A(n514), .B(n425), .C(n520), .D(n164), .E(n524), .F(n365), 
        .G(n429), .H(intadd_23_SUM_2_), .Y(n801) );
  scg4d1_hd U1595 ( .A(n553), .B(n220), .C(n543), .D(n407), .E(n152), .F(n547), 
        .G(n412), .H(intadd_23_SUM_8_), .Y(n802) );
  ivd1_hd U1596 ( .A(intadd_24_SUM_8_), .Y(intadd_20_B_11_) );
  ivd1_hd U1597 ( .A(intadd_20_SUM_11_), .Y(intadd_22_A_14_) );
  scg4d1_hd U1598 ( .A(n580), .B(n361), .C(n570), .D(n908), .E(n137), .F(n576), 
        .G(n398), .H(n60), .Y(n803) );
  ivd1_hd U1599 ( .A(intadd_21_SUM_17_), .Y(N197) );
  oa22d1_hd U1600 ( .A(n594), .B(n601), .C(n596), .D(intadd_23_A_17_), .Y(n804) );
  ivd1_hd U1601 ( .A(n804), .Y(n1068) );
  scg4d1_hd U1602 ( .A(n593), .B(n133), .C(n587), .D(n384), .E(n852), .F(n67), 
        .G(n210), .H(n597), .Y(n805) );
  scg4d1_hd U1603 ( .A(n565), .B(n145), .C(b_m[14]), .D(n401), .E(n403), .F(
        n52), .G(intadd_23_B_13_), .H(n216), .Y(n806) );
  scg4d1_hd U1604 ( .A(n536), .B(n154), .C(n543), .D(n227), .E(n533), .F(n417), 
        .G(n419), .H(n40), .Y(n807) );
  scg4d1_hd U1605 ( .A(b_m[7]), .B(n366), .C(n521), .D(n424), .E(n165), .F(
        n525), .G(n429), .H(intadd_23_SUM_3_), .Y(n808) );
  ao21d1_hd U1606 ( .A(n814), .B(n810), .C(n809), .Y(intadd_27_A_0_) );
  nr2d1_hd U1607 ( .A(n619), .B(a_m[22]), .Y(n1095) );
  ao21d1_hd U1608 ( .A(a_m[22]), .B(n616), .C(n1095), .Y(n829) );
  ao22d1_hd U1609 ( .A(n180), .B(n182), .C(n72), .D(n443), .Y(n813) );
  oa21d1_hd U1610 ( .A(n88), .B(n1050), .C(n813), .Y(n817) );
  nr2d1_hd U1611 ( .A(n615), .B(n817), .Y(n815) );
  nr2bd1_hd U1612 ( .AN(n814), .B(n610), .Y(n816) );
  ao211d1_hd U1613 ( .A(n610), .B(n817), .C(n816), .D(n815), .Y(n818) );
  nr2bd1_hd U1614 ( .AN(n833), .B(n818), .Y(intadd_27_B_0_) );
  scg4d1_hd U1615 ( .A(n514), .B(n170), .C(n506), .D(n433), .E(n371), .F(
        b_m[3]), .G(n436), .H(n29), .Y(n819) );
  ivd1_hd U1616 ( .A(intadd_27_SUM_0_), .Y(intadd_25_B_3_) );
  scg4d1_hd U1617 ( .A(n553), .B(n153), .C(n556), .D(n221), .E(n547), .F(n409), 
        .G(n412), .H(intadd_23_SUM_9_), .Y(n820) );
  ivd1_hd U1618 ( .A(intadd_24_SUM_9_), .Y(intadd_20_B_12_) );
  ivd1_hd U1619 ( .A(intadd_20_SUM_12_), .Y(intadd_22_A_15_) );
  scg4d1_hd U1620 ( .A(n580), .B(n139), .C(n574), .D(n391), .E(n583), .F(n362), 
        .G(n396), .H(n58), .Y(n821) );
  ivd1_hd U1621 ( .A(intadd_21_SUM_18_), .Y(N198) );
  scg4d1_hd U1622 ( .A(n593), .B(n851), .C(n598), .D(n134), .E(b_m[23]), .F(
        n211), .G(n388), .H(n27), .Y(n824) );
  scg4d1_hd U1623 ( .A(n565), .B(n399), .C(n571), .D(n147), .E(n403), .F(n56), 
        .G(n574), .H(n217), .Y(n825) );
  scg4d1_hd U1624 ( .A(n546), .B(n228), .C(b_m[10]), .D(n159), .E(n417), .F(
        b_m[9]), .G(n419), .H(n44), .Y(n826) );
  scg4d1_hd U1625 ( .A(n526), .B(n166), .C(n522), .D(n424), .E(n533), .F(n367), 
        .G(n429), .H(intadd_23_SUM_4_), .Y(n827) );
  scg4d1_hd U1626 ( .A(n504), .B(n183), .C(n176), .D(n373), .E(n442), .F(n125), 
        .G(n76), .H(n443), .Y(n832) );
  nr2d1_hd U1627 ( .A(n834), .B(n833), .Y(n856) );
  ao21d1_hd U1628 ( .A(n834), .B(n833), .C(n856), .Y(intadd_27_A_1_) );
  scg4d1_hd U1629 ( .A(b_m[4]), .B(n368), .C(n510), .D(n432), .E(b_m[5]), .F(
        n175), .G(n437), .H(n33), .Y(n835) );
  ivd1_hd U1630 ( .A(intadd_27_SUM_1_), .Y(intadd_25_B_4_) );
  scg4d1_hd U1631 ( .A(n553), .B(n408), .C(n556), .D(n149), .E(n562), .F(n218), 
        .G(n412), .H(intadd_23_SUM_10_), .Y(n836) );
  ivd1_hd U1632 ( .A(intadd_24_SUM_10_), .Y(intadd_20_B_13_) );
  ivd1_hd U1633 ( .A(intadd_20_SUM_13_), .Y(intadd_22_A_16_) );
  scg4d1_hd U1634 ( .A(n580), .B(n393), .C(n582), .D(n140), .E(n588), .F(n363), 
        .G(n398), .H(n66), .Y(n837) );
  ivd1_hd U1635 ( .A(intadd_21_SUM_19_), .Y(N199) );
  scg4d1_hd U1636 ( .A(n580), .B(n214), .C(n571), .D(n401), .E(n403), .F(n60), 
        .G(n143), .H(intadd_23_B_14_), .Y(n838) );
  scg4d1_hd U1637 ( .A(n551), .B(n359), .C(b_m[10]), .D(n415), .E(n162), .F(
        n548), .G(n419), .H(n46), .Y(n839) );
  scg4d1_hd U1638 ( .A(n526), .B(n425), .C(n531), .D(n167), .E(n537), .F(n364), 
        .G(n429), .H(intadd_23_SUM_5_), .Y(n840) );
  scg4d1_hd U1639 ( .A(n509), .B(n184), .C(n178), .D(n441), .E(n74), .F(n445), 
        .G(n503), .H(n374), .Y(n842) );
  xo3d1_hd U1640 ( .A(n857), .B(n856), .C(n858), .Y(intadd_27_A_2_) );
  scg4d1_hd U1641 ( .A(n514), .B(n433), .C(n521), .D(n369), .E(b_m[6]), .F(
        n168), .G(n436), .H(n31), .Y(n843) );
  ivd1_hd U1642 ( .A(intadd_27_SUM_2_), .Y(intadd_25_B_5_) );
  scg4d1_hd U1643 ( .A(n565), .B(n219), .C(n557), .D(n407), .E(n150), .F(n563), 
        .G(n414), .H(intadd_23_SUM_11_), .Y(n844) );
  ivd1_hd U1644 ( .A(intadd_24_SUM_11_), .Y(intadd_20_B_14_) );
  ivd1_hd U1645 ( .A(intadd_20_SUM_14_), .Y(intadd_22_A_17_) );
  scg4d1_hd U1646 ( .A(n593), .B(n360), .C(n582), .D(n908), .E(n142), .F(n589), 
        .G(n398), .H(n64), .Y(n845) );
  ao22d1_hd U1647 ( .A(n599), .B(n384), .C(n388), .D(n61), .Y(n848) );
  oa21d1_hd U1648 ( .A(n127), .B(n849), .C(n848), .Y(n850) );
  ivd1_hd U1649 ( .A(intadd_21_SUM_20_), .Y(N200) );
  ao21d1_hd U1650 ( .A(n1065), .B(n388), .C(n384), .Y(n853) );
  nr2d1_hd U1651 ( .A(n128), .B(n853), .Y(n854) );
  scg4d1_hd U1652 ( .A(n579), .B(n144), .C(n574), .D(n402), .E(n405), .F(n58), 
        .G(intadd_23_B_16_), .H(n215), .Y(n855) );
  ivd1_hd U1653 ( .A(n856), .Y(n859) );
  ao21d1_hd U1654 ( .A(n859), .B(n858), .C(n857), .Y(n874) );
  nr2d1_hd U1655 ( .A(n614), .B(n197), .Y(n873) );
  scg4d1_hd U1656 ( .A(n514), .B(n182), .C(b_m[2]), .D(n441), .E(n372), .F(
        n511), .G(n444), .H(intadd_23_SUM_0_), .Y(n860) );
  scg4d1_hd U1657 ( .A(n526), .B(n169), .C(n521), .D(n432), .E(n370), .F(n525), 
        .G(n436), .H(n35), .Y(n861) );
  ivd1_hd U1658 ( .A(intadd_27_SUM_3_), .Y(intadd_25_A_6_) );
  scg4d1_hd U1659 ( .A(n535), .B(n165), .C(b_m[10]), .D(n366), .E(n533), .F(
        n426), .G(n427), .H(intadd_23_SUM_6_), .Y(n862) );
  scg4d1_hd U1660 ( .A(n551), .B(n163), .C(n557), .D(n226), .E(n547), .F(n417), 
        .G(n995), .H(n48), .Y(n863) );
  scg4d1_hd U1661 ( .A(n565), .B(n152), .C(n561), .D(n410), .E(n571), .F(n220), 
        .G(n414), .H(intadd_23_SUM_12_), .Y(n864) );
  ivd1_hd U1662 ( .A(intadd_24_SUM_12_), .Y(intadd_20_B_15_) );
  ivd1_hd U1663 ( .A(intadd_20_SUM_15_), .Y(intadd_22_A_18_) );
  scg4d1_hd U1664 ( .A(n593), .B(n137), .C(n586), .D(n908), .E(n599), .F(n361), 
        .G(n395), .H(n68), .Y(n865) );
  ivd1_hd U1665 ( .A(intadd_21_SUM_21_), .Y(N201) );
  scg4d1_hd U1666 ( .A(n593), .B(n393), .C(n598), .D(n139), .E(n109), .F(n362), 
        .G(n909), .H(n27), .Y(n867) );
  scg4d1_hd U1667 ( .A(n579), .B(n935), .C(n583), .D(n145), .E(n405), .F(
        intadd_23_SUM_16_), .G(n586), .H(n216), .Y(n868) );
  scg4d1_hd U1668 ( .A(n566), .B(n408), .C(n570), .D(n153), .E(n575), .F(n221), 
        .G(n414), .H(intadd_23_SUM_13_), .Y(n869) );
  scg4d1_hd U1669 ( .A(b_m[12]), .B(n416), .C(b_m[13]), .D(n154), .E(n562), 
        .F(n227), .G(n995), .H(n50), .Y(n870) );
  scg4d1_hd U1670 ( .A(n545), .B(n365), .C(n541), .D(n164), .E(n426), .F(n538), 
        .G(n427), .H(intadd_23_SUM_7_), .Y(n871) );
  fad1_hd U1671 ( .A(n874), .B(n873), .CI(n872), .CO(n887), .S(intadd_27_A_3_)
         );
  scg4d1_hd U1672 ( .A(intadd_23_B_1_), .B(n375), .C(n510), .D(n440), .E(n518), 
        .F(n185), .G(n444), .H(intadd_23_SUM_1_), .Y(n875) );
  ivd1_hd U1673 ( .A(n876), .Y(n886) );
  scg4d1_hd U1674 ( .A(b_m[7]), .B(n371), .C(n523), .D(n432), .E(n533), .F(
        n170), .G(n1042), .H(n38), .Y(n877) );
  ivd1_hd U1675 ( .A(intadd_27_SUM_4_), .Y(intadd_25_B_7_) );
  ivd1_hd U1676 ( .A(intadd_24_SUM_13_), .Y(intadd_20_B_16_) );
  ivd1_hd U1677 ( .A(intadd_20_SUM_16_), .Y(intadd_21_B_22_) );
  ivd1_hd U1678 ( .A(intadd_21_SUM_22_), .Y(N202) );
  scg4d1_hd U1679 ( .A(n593), .B(n217), .C(b_m[19]), .D(n401), .E(n936), .F(
        intadd_23_SUM_17_), .G(n147), .H(intadd_23_B_17_), .Y(n878) );
  ao22d1_hd U1680 ( .A(b_m[22]), .B(n908), .C(n395), .D(n62), .Y(n879) );
  oa21d1_hd U1681 ( .A(n128), .B(n880), .C(n879), .Y(n881) );
  scg4d1_hd U1682 ( .A(n566), .B(n228), .C(b_m[13]), .D(n415), .E(n159), .F(
        n562), .G(n422), .H(n54), .Y(n882) );
  scg4d1_hd U1683 ( .A(n579), .B(n218), .C(b_m[16]), .D(n967), .E(n149), .F(
        n576), .G(n414), .H(intadd_23_SUM_14_), .Y(n883) );
  scg4d1_hd U1684 ( .A(b_m[12]), .B(n367), .C(n541), .D(n424), .E(n166), .F(
        n548), .G(n427), .H(intadd_23_SUM_8_), .Y(n884) );
  fad1_hd U1685 ( .A(n887), .B(n886), .CI(n885), .CO(intadd_27_A_5_), .S(
        intadd_27_B_4_) );
  fad1_hd U1686 ( .A(n473), .B(n889), .CI(n888), .CO(n900), .S(n876) );
  scg4d1_hd U1687 ( .A(n526), .B(n433), .C(n531), .D(n368), .E(n537), .F(n175), 
        .G(n1042), .H(n42), .Y(n890) );
  nr2d1_hd U1688 ( .A(n613), .B(n513), .Y(intadd_28_B_0_) );
  scg4d1_hd U1689 ( .A(intadd_23_B_1_), .B(n441), .C(n521), .D(n373), .E(n524), 
        .F(n183), .G(n444), .H(intadd_23_SUM_2_), .Y(n891) );
  ivd1_hd U1690 ( .A(intadd_28_SUM_0_), .Y(n898) );
  ivd1_hd U1691 ( .A(n892), .Y(intadd_27_B_5_) );
  ivd1_hd U1692 ( .A(intadd_27_SUM_5_), .Y(intadd_25_B_8_) );
  ivd1_hd U1693 ( .A(n893), .Y(intadd_20_B_17_) );
  scg4d1_hd U1694 ( .A(b_m[15]), .B(n162), .C(n561), .D(n418), .E(n570), .F(
        n359), .G(n422), .H(n52), .Y(n897) );
  fad1_hd U1695 ( .A(n900), .B(n899), .CI(n898), .CO(n901), .S(n892) );
  ivd1_hd U1696 ( .A(n901), .Y(intadd_28_A_1_) );
  nr2d1_hd U1697 ( .A(n613), .B(n517), .Y(intadd_32_B_0_) );
  scg4d1_hd U1698 ( .A(n526), .B(n184), .C(n521), .D(n440), .E(n374), .F(n525), 
        .G(n444), .H(intadd_23_SUM_3_), .Y(n902) );
  scg4d1_hd U1699 ( .A(n535), .B(n369), .C(n541), .D(n168), .E(b_m[8]), .F(
        n434), .G(n437), .H(n40), .Y(n903) );
  ivd1_hd U1700 ( .A(intadd_27_SUM_6_), .Y(intadd_25_A_9_) );
  scg4d1_hd U1701 ( .A(n551), .B(n167), .C(b_m[13]), .D(n364), .E(n547), .F(
        n426), .G(n1022), .H(intadd_23_SUM_9_), .Y(n904) );
  scg4d1_hd U1702 ( .A(n579), .B(n150), .C(n573), .D(n407), .E(n583), .F(n219), 
        .G(n412), .H(intadd_23_SUM_15_), .Y(n905) );
  fad1_hd U1703 ( .A(n907), .B(n906), .CI(intadd_25_SUM_8_), .CO(
        intadd_24_B_15_), .S(intadd_24_B_14_) );
  ivd1_hd U1704 ( .A(intadd_24_SUM_15_), .Y(n915) );
  ao21d1_hd U1705 ( .A(n395), .B(n1065), .C(n908), .Y(n910) );
  nr2d1_hd U1706 ( .A(n126), .B(n910), .Y(n911) );
  scg4d1_hd U1707 ( .A(n592), .B(n143), .C(n586), .D(n401), .E(n404), .F(n67), 
        .G(n597), .H(n214), .Y(n912) );
  scg4d1_hd U1708 ( .A(n579), .B(n409), .C(n582), .D(n153), .E(n587), .F(n221), 
        .G(n411), .H(n66), .Y(n916) );
  scg4d1_hd U1709 ( .A(b_m[15]), .B(n416), .C(b_m[16]), .D(n154), .E(n575), 
        .F(n227), .G(n422), .H(n56), .Y(n917) );
  scg4d1_hd U1710 ( .A(intadd_23_B_4_), .B(n372), .C(n522), .D(n440), .E(n533), 
        .F(n182), .G(n444), .H(intadd_23_SUM_4_), .Y(n918) );
  ivd1_hd U1711 ( .A(intadd_29_SUM_0_), .Y(intadd_32_B_1_) );
  scg4d1_hd U1712 ( .A(n546), .B(n169), .C(b_m[10]), .D(n370), .E(n434), .F(
        n538), .G(n437), .H(n44), .Y(n919) );
  scg4d1_hd U1713 ( .A(n552), .B(n425), .C(n555), .D(n164), .E(n562), .F(n365), 
        .G(n1022), .H(intadd_23_SUM_10_), .Y(n920) );
  ivd1_hd U1714 ( .A(intadd_27_SUM_7_), .Y(intadd_25_B_10_) );
  scg4d1_hd U1715 ( .A(n592), .B(n935), .C(n597), .D(n144), .E(n404), .F(n27), 
        .G(n1117), .H(n215), .Y(n921) );
  ivd1_hd U1716 ( .A(intadd_29_B_2_), .Y(intadd_29_A_1_) );
  scg4d1_hd U1717 ( .A(intadd_23_B_4_), .B(n441), .C(b_m[8]), .D(n375), .E(
        n537), .F(n185), .G(n444), .H(intadd_23_SUM_5_), .Y(n922) );
  ivd1_hd U1718 ( .A(intadd_29_SUM_1_), .Y(intadd_32_A_2_) );
  scg4d1_hd U1719 ( .A(n552), .B(n170), .C(n541), .D(n432), .E(n371), .F(n548), 
        .G(n437), .H(n46), .Y(n923) );
  scg4d1_hd U1720 ( .A(b_m[15]), .B(n366), .C(n555), .D(n424), .E(n165), .F(
        n563), .G(n430), .H(intadd_23_SUM_11_), .Y(n924) );
  scg4d1_hd U1721 ( .A(n578), .B(n226), .C(b_m[16]), .D(n994), .E(n163), .F(
        n575), .G(n422), .H(n60), .Y(n925) );
  ivd1_hd U1722 ( .A(intadd_27_SUM_8_), .Y(intadd_25_A_11_) );
  scg4d1_hd U1723 ( .A(n592), .B(n220), .C(n583), .D(n967), .E(n152), .F(n588), 
        .G(n414), .H(n64), .Y(n926) );
  ao22d1_hd U1724 ( .A(b_m[22]), .B(n400), .C(n404), .D(n61), .Y(n927) );
  oa21d1_hd U1725 ( .A(n127), .B(n928), .C(n927), .Y(n929) );
  ivd1_hd U1726 ( .A(intadd_39_SUM_2_), .Y(intadd_20_A_20_) );
  ivd1_hd U1727 ( .A(intadd_24_n1), .Y(intadd_20_B_20_) );
  scg4d1_hd U1728 ( .A(n592), .B(n149), .C(b_m[20]), .D(n967), .E(n598), .F(
        n218), .G(n968), .H(n68), .Y(n930) );
  ivd1_hd U1729 ( .A(intadd_25_n1), .Y(intadd_27_A_9_) );
  nr2d1_hd U1730 ( .A(n613), .B(n530), .Y(intadd_29_A_2_) );
  scg4d1_hd U1731 ( .A(n535), .B(n373), .C(n541), .D(n183), .E(b_m[8]), .F(
        n442), .G(n446), .H(intadd_23_SUM_6_), .Y(n931) );
  scg4d1_hd U1732 ( .A(n552), .B(n368), .C(n555), .D(n175), .E(n547), .F(n434), 
        .G(n437), .H(n48), .Y(n932) );
  ivd1_hd U1733 ( .A(intadd_38_SUM_0_), .Y(intadd_28_B_4_) );
  ivd1_hd U1734 ( .A(intadd_28_SUM_4_), .Y(intadd_37_A_0_) );
  scg4d1_hd U1735 ( .A(n564), .B(n166), .C(n561), .D(n1021), .E(n571), .F(n367), .G(n430), .H(intadd_23_SUM_12_), .Y(n933) );
  scg4d1_hd U1736 ( .A(n578), .B(n159), .C(b_m[17]), .D(n415), .E(n582), .F(
        n228), .G(n995), .H(n58), .Y(n934) );
  ivd1_hd U1737 ( .A(intadd_37_SUM_0_), .Y(intadd_27_B_9_) );
  ivd1_hd U1738 ( .A(intadd_27_SUM_9_), .Y(n948) );
  ao21d1_hd U1739 ( .A(n1065), .B(n404), .C(n400), .Y(n937) );
  nr2d1_hd U1740 ( .A(n127), .B(n937), .Y(n938) );
  ivd1_hd U1741 ( .A(n939), .Y(intadd_20_A_21_) );
  ivd1_hd U1742 ( .A(intadd_39_n1), .Y(intadd_20_B_21_) );
  scg4d1_hd U1743 ( .A(n546), .B(n184), .C(intadd_23_B_7_), .D(n374), .E(n442), 
        .F(n538), .G(n446), .H(intadd_23_SUM_7_), .Y(n940) );
  nr2bd1_hd U1744 ( .AN(n941), .B(intadd_29_A_2_), .Y(n952) );
  nr2d1_hd U1745 ( .A(n530), .B(n941), .Y(n951) );
  nr2d1_hd U1746 ( .A(n952), .B(n951), .Y(n942) );
  scg4d1_hd U1747 ( .A(n552), .B(n433), .C(b_m[13]), .D(n369), .E(n561), .F(
        n168), .G(n436), .H(n50), .Y(n943) );
  ivd1_hd U1748 ( .A(intadd_38_SUM_1_), .Y(intadd_28_A_5_) );
  scg4d1_hd U1749 ( .A(n564), .B(n425), .C(n569), .D(n167), .E(n575), .F(n364), 
        .G(n430), .H(intadd_23_SUM_13_), .Y(n944) );
  ivd1_hd U1750 ( .A(intadd_28_SUM_5_), .Y(intadd_37_A_1_) );
  scg4d1_hd U1751 ( .A(n578), .B(n417), .C(b_m[19]), .D(n162), .E(n587), .F(
        n359), .G(n422), .H(intadd_23_SUM_16_), .Y(n945) );
  ivd1_hd U1752 ( .A(intadd_37_SUM_1_), .Y(intadd_27_A_10_) );
  scg4d1_hd U1753 ( .A(n592), .B(n409), .C(n598), .D(n150), .E(b_m[23]), .F(
        n219), .G(n968), .H(n1048), .Y(n946) );
  ivd1_hd U1754 ( .A(intadd_31_A_0_), .Y(n963) );
  scg20d1_hd U1755 ( .A(n605), .B(n952), .C(n951), .Y(n962) );
  scg4d1_hd U1756 ( .A(n551), .B(n185), .C(intadd_23_B_7_), .D(n440), .E(n375), 
        .F(n548), .G(n1066), .H(intadd_23_SUM_8_), .Y(n953) );
  scg4d1_hd U1757 ( .A(n564), .B(n169), .C(n555), .D(n432), .E(n370), .F(n563), 
        .G(n438), .H(n54), .Y(n954) );
  scg4d1_hd U1758 ( .A(n578), .B(n365), .C(n569), .D(n423), .E(n164), .F(n576), 
        .G(n430), .H(intadd_23_SUM_14_), .Y(n955) );
  ivd1_hd U1759 ( .A(intadd_38_SUM_2_), .Y(intadd_28_A_6_) );
  scg4d1_hd U1760 ( .A(n592), .B(n226), .C(b_m[19]), .D(n994), .E(n163), .F(
        n589), .G(n419), .H(intadd_23_SUM_17_), .Y(n956) );
  ivd1_hd U1761 ( .A(intadd_28_SUM_6_), .Y(intadd_37_A_2_) );
  ao22d1_hd U1762 ( .A(b_m[22]), .B(n967), .C(n968), .D(n62), .Y(n957) );
  oa21d1_hd U1763 ( .A(n128), .B(n958), .C(n957), .Y(n959) );
  scg4d1_hd U1764 ( .A(n591), .B(n154), .C(n587), .D(n994), .E(n599), .F(n227), 
        .G(n420), .H(n67), .Y(n960) );
  ivd1_hd U1765 ( .A(intadd_38_n1), .Y(intadd_28_A_7_) );
  fad1_hd U1766 ( .A(n963), .B(n962), .CI(n961), .CO(intadd_29_A_5_), .S(
        intadd_29_A_4_) );
  nr2d1_hd U1767 ( .A(n613), .B(n544), .Y(intadd_31_B_0_) );
  scg4d1_hd U1768 ( .A(n552), .B(n372), .C(n555), .D(n182), .E(n547), .F(n442), 
        .G(n1066), .H(intadd_23_SUM_9_), .Y(n964) );
  ivd1_hd U1769 ( .A(intadd_31_SUM_0_), .Y(intadd_29_B_5_) );
  scg4d1_hd U1770 ( .A(b_m[15]), .B(n371), .C(b_m[14]), .D(n1041), .E(n570), 
        .F(n170), .G(n438), .H(n52), .Y(n965) );
  scg4d1_hd U1771 ( .A(n578), .B(n165), .C(b_m[17]), .D(n424), .E(n583), .F(
        n366), .G(n1022), .H(intadd_23_SUM_15_), .Y(n966) );
  ivd1_hd U1772 ( .A(intadd_36_SUM_0_), .Y(intadd_28_B_7_) );
  ivd1_hd U1773 ( .A(intadd_28_SUM_7_), .Y(n980) );
  ao21d1_hd U1774 ( .A(n968), .B(n196), .C(n967), .Y(n969) );
  nr2d1_hd U1775 ( .A(n126), .B(n969), .Y(n970) );
  scg4d1_hd U1776 ( .A(n552), .B(n441), .C(intadd_23_B_10_), .D(n373), .E(n562), .F(n183), .G(n1066), .H(intadd_23_SUM_10_), .Y(n972) );
  nr2d1_hd U1777 ( .A(intadd_23_B_8_), .B(intadd_23_B_6_), .Y(n973) );
  ao211d1_hd U1778 ( .A(intadd_23_B_8_), .B(intadd_23_B_6_), .C(n610), .D(n973), .Y(n974) );
  ivd1_hd U1779 ( .A(intadd_31_SUM_1_), .Y(intadd_29_A_6_) );
  scg4d1_hd U1780 ( .A(n564), .B(n433), .C(b_m[16]), .D(n369), .E(n573), .F(
        n168), .G(n438), .H(n56), .Y(n975) );
  scg4d1_hd U1781 ( .A(n577), .B(n426), .C(n581), .D(n166), .E(n588), .F(n364), 
        .G(n427), .H(n66), .Y(n976) );
  ivd1_hd U1782 ( .A(intadd_36_SUM_1_), .Y(intadd_28_A_8_) );
  scg4d1_hd U1783 ( .A(n591), .B(n417), .C(n597), .D(n159), .E(n109), .F(n228), 
        .G(n420), .H(n27), .Y(n978) );
  ivd1_hd U1784 ( .A(intadd_30_B_1_), .Y(intadd_30_A_0_) );
  nr2d1_hd U1785 ( .A(a_m[11]), .B(intadd_31_A_0_), .Y(n984) );
  ao211d1_hd U1786 ( .A(n84), .B(n540), .C(n610), .D(n550), .Y(n983) );
  nr2d1_hd U1787 ( .A(n984), .B(n983), .Y(intadd_30_B_0_) );
  scg4d1_hd U1788 ( .A(n564), .B(n184), .C(intadd_23_B_10_), .D(n440), .E(n374), .F(n563), .G(n445), .H(intadd_23_SUM_11_), .Y(n985) );
  ivd1_hd U1789 ( .A(intadd_30_SUM_0_), .Y(intadd_31_A_2_) );
  scg4d1_hd U1790 ( .A(n577), .B(n175), .C(n569), .D(n431), .E(n368), .F(n576), 
        .G(n438), .H(n60), .Y(n986) );
  ivd1_hd U1791 ( .A(intadd_31_SUM_2_), .Y(intadd_29_A_7_) );
  scg4d1_hd U1792 ( .A(n591), .B(n367), .C(n581), .D(n423), .E(n167), .F(n589), 
        .G(n430), .H(n64), .Y(n987) );
  ao22d1_hd U1793 ( .A(b_m[22]), .B(n994), .C(n420), .D(n61), .Y(n988) );
  oa21d1_hd U1794 ( .A(n127), .B(n989), .C(n988), .Y(n990) );
  scg4d1_hd U1795 ( .A(n591), .B(n164), .C(b_m[20]), .D(n423), .E(n599), .F(
        n365), .G(n428), .H(n68), .Y(n991) );
  ivd1_hd U1796 ( .A(intadd_29_n1), .Y(intadd_31_A_3_) );
  scg4d1_hd U1797 ( .A(intadd_23_B_12_), .B(n375), .C(n561), .D(n439), .E(n571), .F(n185), .G(n445), .H(intadd_23_SUM_12_), .Y(n992) );
  scg4d1_hd U1798 ( .A(n577), .B(n370), .C(n574), .D(n432), .E(n582), .F(n169), 
        .G(n436), .H(n58), .Y(n993) );
  nr2d1_hd U1799 ( .A(n613), .B(n559), .Y(intadd_30_A_1_) );
  ivd1_hd U1800 ( .A(intadd_35_SUM_0_), .Y(intadd_31_B_3_) );
  ivd1_hd U1801 ( .A(intadd_31_SUM_3_), .Y(n1006) );
  ao21d1_hd U1802 ( .A(n420), .B(n196), .C(n994), .Y(n996) );
  nr2d1_hd U1803 ( .A(n108), .B(n996), .Y(n997) );
  scg4d1_hd U1804 ( .A(intadd_23_B_12_), .B(n441), .C(n569), .D(n372), .E(n575), .F(n182), .G(n445), .H(intadd_23_SUM_13_), .Y(n999) );
  nr2bd1_hd U1805 ( .AN(n1000), .B(intadd_30_A_1_), .Y(n1010) );
  nr2d1_hd U1806 ( .A(n559), .B(n1000), .Y(n1009) );
  nr2d1_hd U1807 ( .A(n1010), .B(n1009), .Y(n1001) );
  scg4d1_hd U1808 ( .A(n577), .B(n434), .C(b_m[19]), .D(n371), .E(n588), .F(
        n170), .G(n438), .H(intadd_23_SUM_16_), .Y(n1002) );
  ivd1_hd U1809 ( .A(intadd_35_SUM_1_), .Y(intadd_31_A_4_) );
  scg4d1_hd U1810 ( .A(n591), .B(n426), .C(n597), .D(n165), .E(b_m[23]), .F(
        n366), .G(n428), .H(n1048), .Y(n1004) );
  nr2d1_hd U1811 ( .A(n614), .B(n568), .Y(n1019) );
  scg20d1_hd U1812 ( .A(n86), .B(n1010), .C(n1009), .Y(n1018) );
  scg4d1_hd U1813 ( .A(n578), .B(n183), .C(n569), .D(n439), .E(n373), .F(n576), 
        .G(n445), .H(intadd_23_SUM_14_), .Y(n1011) );
  scg4d1_hd U1814 ( .A(n590), .B(n175), .C(n581), .D(n431), .E(n368), .F(n589), 
        .G(n1042), .H(intadd_23_SUM_17_), .Y(n1012) );
  ao22d1_hd U1815 ( .A(n596), .B(n423), .C(n428), .D(n62), .Y(n1013) );
  oa21d1_hd U1816 ( .A(n128), .B(n1014), .C(n1013), .Y(n1015) );
  scg4d1_hd U1817 ( .A(n590), .B(n369), .C(n587), .D(n431), .E(n599), .F(n168), 
        .G(n435), .H(n67), .Y(n1016) );
  fad1_hd U1818 ( .A(n1019), .B(n1018), .CI(n1017), .CO(intadd_30_A_4_), .S(
        intadd_30_A_3_) );
  ivd1_hd U1819 ( .A(n1019), .Y(intadd_33_A_0_) );
  nr2d1_hd U1820 ( .A(n614), .B(n572), .Y(intadd_33_B_0_) );
  scg4d1_hd U1821 ( .A(b_m[18]), .B(n374), .C(n573), .D(n440), .E(n583), .F(
        n184), .G(n1066), .H(intadd_23_SUM_15_), .Y(n1020) );
  ivd1_hd U1822 ( .A(intadd_33_SUM_0_), .Y(intadd_30_B_4_) );
  ao21d1_hd U1823 ( .A(n428), .B(n196), .C(n1021), .Y(n1023) );
  nr2d1_hd U1824 ( .A(n126), .B(n1023), .Y(n1024) );
  ivd1_hd U1825 ( .A(n1025), .Y(intadd_20_A_30_) );
  ivd1_hd U1826 ( .A(intadd_35_n1), .Y(intadd_20_B_30_) );
  scg4d1_hd U1827 ( .A(b_m[18]), .B(n442), .C(n581), .D(n375), .E(n588), .F(
        n185), .G(n445), .H(n66), .Y(n1026) );
  nr2d1_hd U1828 ( .A(n568), .B(n1027), .Y(n1034) );
  nr2bd1_hd U1829 ( .AN(n1035), .B(n1034), .Y(n1028) );
  ivd1_hd U1830 ( .A(intadd_33_SUM_1_), .Y(intadd_30_A_5_) );
  scg4d1_hd U1831 ( .A(n591), .B(n434), .C(n598), .D(n370), .E(n109), .F(n169), 
        .G(n435), .H(n27), .Y(n1030) );
  fad1_hd U1832 ( .A(n1032), .B(intadd_30_SUM_4_), .CI(n1031), .CO(n1033), .S(
        n1025) );
  ivd1_hd U1833 ( .A(intadd_34_B_1_), .Y(intadd_34_A_0_) );
  ao21d1_hd U1834 ( .A(n459), .B(n1035), .C(n1034), .Y(intadd_34_B_0_) );
  ivd1_hd U1835 ( .A(intadd_34_SUM_0_), .Y(intadd_33_A_2_) );
  ao22d1_hd U1836 ( .A(b_m[22]), .B(n431), .C(n435), .D(n61), .Y(n1037) );
  oa21d1_hd U1837 ( .A(n108), .B(n1029), .C(n1037), .Y(n1038) );
  scg4d1_hd U1838 ( .A(n590), .B(n373), .C(n587), .D(n1064), .E(n599), .F(n183), .G(n443), .H(n68), .Y(n1040) );
  nr2d1_hd U1839 ( .A(n614), .B(n585), .Y(intadd_34_A_1_) );
  ao21d1_hd U1840 ( .A(n435), .B(n196), .C(n431), .Y(n1043) );
  nr2d1_hd U1841 ( .A(n126), .B(n1043), .Y(n1044) );
  nr2bd1_hd U1842 ( .AN(n1046), .B(intadd_34_A_1_), .Y(n1059) );
  nr2d1_hd U1843 ( .A(n585), .B(n1046), .Y(n1058) );
  nr2d1_hd U1844 ( .A(n1059), .B(n1058), .Y(n1047) );
  scg4d1_hd U1845 ( .A(n590), .B(n442), .C(n598), .D(n374), .E(n109), .F(n184), 
        .G(n443), .H(n1048), .Y(n1051) );
  ivd1_hd U1846 ( .A(intadd_34_SUM_2_), .Y(intadd_20_A_34_) );
  ivd1_hd U1847 ( .A(n1054), .Y(intadd_20_B_34_) );
  ao22d1_hd U1848 ( .A(n596), .B(n1064), .C(n443), .D(n62), .Y(n1056) );
  oa21d1_hd U1849 ( .A(n127), .B(n1050), .C(n1056), .Y(n1057) );
  nr2d1_hd U1850 ( .A(n614), .B(n595), .Y(n1075) );
  scg20d1_hd U1851 ( .A(a_m[20]), .B(n1059), .C(n1058), .Y(n1061) );
  fad1_hd U1852 ( .A(n1062), .B(n1075), .CI(n1061), .CO(n1063), .S(n1060) );
  ao21d1_hd U1853 ( .A(n443), .B(n196), .C(n1064), .Y(n1067) );
  nr2d1_hd U1854 ( .A(n108), .B(n1067), .Y(n1069) );
  oa21d1_hd U1855 ( .A(n617), .B(n1069), .C(n1072), .Y(n1074) );
  scg16d1_hd U1856 ( .A(n1072), .B(n1071), .C(n1070), .Y(intadd_20_B_36_) );
  oa211d1_hd U1857 ( .A(n595), .B(n1072), .C(n617), .D(n597), .Y(n1073) );
  oa21d1_hd U1858 ( .A(n1075), .B(n1074), .C(n1073), .Y(n1078) );
  oa211d1_hd U1859 ( .A(intadd_23_A_17_), .B(n126), .C(n617), .D(n1076), .Y(
        n1077) );
  ivd1_hd U1860 ( .A(b_e[9]), .Y(n1422) );
  ivd1_hd U1861 ( .A(a_e[9]), .Y(n1362) );
  ao22d1_hd U1862 ( .A(a_e[9]), .B(b_e[9]), .C(n1422), .D(n1362), .Y(n1081) );
  nr2d1_hd U1863 ( .A(DP_OP_125J2_130_6300_n12), .B(n1081), .Y(n1080) );
  ao211d1_hd U1864 ( .A(DP_OP_125J2_130_6300_n12), .B(n1081), .C(n498), .D(
        n1080), .Y(n1082) );
  ao21d1_hd U1865 ( .A(z_e[9]), .B(n90), .C(n1082), .Y(n1083) );
  ivd1_hd U1866 ( .A(n1188), .Y(n1427) );
  ao21d1_hd U1867 ( .A(n455), .B(product[25]), .C(n1085), .Y(n104) );
  nr2d1_hd U1868 ( .A(z_e[4]), .B(z_e[3]), .Y(n1087) );
  nr2d1_hd U1869 ( .A(z_e[6]), .B(z_e[5]), .Y(n1086) );
  nr3d1_hd U1870 ( .A(z_e[2]), .B(z_e[1]), .C(n1146), .Y(n1088) );
  oa21d1_hd U1871 ( .A(n1088), .B(n1145), .C(z_e[9]), .Y(n36) );
  ao22d1_hd U1872 ( .A(n482), .B(b[23]), .C(b_e[0]), .D(n102), .Y(n1371) );
  ivd1_hd U1873 ( .A(n1371), .Y(n1207) );
  nr4d1_hd U1874 ( .A(a_e[2]), .B(n10), .C(a_e[6]), .D(n1090), .Y(n1091) );
  ivd1_hd U1875 ( .A(n1091), .Y(n1092) );
  nr4d1_hd U1876 ( .A(a_e[9]), .B(a_e[0]), .C(a_e[8]), .D(n1092), .Y(n1137) );
  nr4d1_hd U1877 ( .A(n1093), .B(b_e[2]), .C(b_e[5]), .D(b_e[4]), .Y(n1106) );
  ivd1_hd U1878 ( .A(n1106), .Y(n1094) );
  nr4d1_hd U1879 ( .A(b_e[8]), .B(b_e[9]), .C(b_e[0]), .D(n1094), .Y(n1135) );
  nr2d1_hd U1880 ( .A(n1137), .B(n1135), .Y(n1144) );
  nd3d1_hd U1881 ( .A(n85), .B(n467), .C(n607), .Y(n1105) );
  nd4d1_hd U1882 ( .A(n1098), .B(n1097), .C(n1096), .D(n1095), .Y(n1104) );
  nr4d1_hd U1883 ( .A(a_m[3]), .B(a_m[0]), .C(a_m[2]), .D(a_m[1]), .Y(n1102)
         );
  nr4d1_hd U1884 ( .A(n120), .B(a_m[21]), .C(a_m[19]), .D(a_m[18]), .Y(n1099)
         );
  nd4d1_hd U1885 ( .A(n1102), .B(n1101), .C(n1100), .D(n1099), .Y(n1103) );
  nr4d1_hd U1886 ( .A(a_m[17]), .B(n1105), .C(n1104), .D(n1103), .Y(n1131) );
  nr2d1_hd U1887 ( .A(intadd_23_B_0_), .B(n502), .Y(n1107) );
  nd4d1_hd U1888 ( .A(n1108), .B(n1107), .C(n594), .D(n127), .Y(n1114) );
  nr4d1_hd U1889 ( .A(intadd_23_B_9_), .B(intadd_23_B_8_), .C(intadd_23_B_4_), 
        .D(intadd_23_B_6_), .Y(n1112) );
  nr4d1_hd U1890 ( .A(intadd_23_B_5_), .B(intadd_23_B_1_), .C(intadd_23_B_3_), 
        .D(intadd_23_B_2_), .Y(n1111) );
  nr4d1_hd U1891 ( .A(intadd_23_B_13_), .B(intadd_23_B_11_), .C(
        intadd_23_B_10_), .D(intadd_23_B_7_), .Y(n1110) );
  nr4d1_hd U1892 ( .A(intadd_23_B_17_), .B(intadd_23_B_16_), .C(
        intadd_23_B_12_), .D(intadd_23_B_14_), .Y(n1109) );
  nd4d1_hd U1893 ( .A(n1112), .B(n1111), .C(n1110), .D(n1109), .Y(n1113) );
  nr4d1_hd U1894 ( .A(n596), .B(intadd_23_B_15_), .C(n1114), .D(n1113), .Y(
        n1133) );
  ao21d1_hd U1895 ( .A(n1363), .B(n99), .C(n482), .Y(n1355) );
  nr2d1_hd U1896 ( .A(n1356), .B(n10), .Y(n1349) );
  ivd1_hd U1897 ( .A(n1349), .Y(n1347) );
  ivd1_hd U1898 ( .A(DP_OP_113J2_124_6892_n3), .Y(n1348) );
  ao22d1_hd U1899 ( .A(DP_OP_113J2_124_6892_n3), .B(n1347), .C(n1349), .D(
        n1348), .Y(n1115) );
  ao22d1_hd U1900 ( .A(n70), .B(a_e[7]), .C(n195), .D(n1115), .Y(n141) );
  ao22d1_hd U1901 ( .A(n481), .B(b[30]), .C(n101), .D(b_e[7]), .Y(n1364) );
  ao22d1_hd U1902 ( .A(n79), .B(b_e[7]), .C(n1418), .D(n1118), .Y(n151) );
  nr3d1_hd U1903 ( .A(n1119), .B(n99), .C(n496), .Y(n156) );
  oa211d1_hd U1904 ( .A(n1123), .B(n77), .C(n1122), .D(n1148), .Y(n1124) );
  nr2d1_hd U1905 ( .A(n1227), .B(n1124), .Y(n160) );
  nr2d1_hd U1906 ( .A(n1126), .B(n1125), .Y(n161) );
  nr2d1_hd U1907 ( .A(n453), .B(n89), .Y(n171) );
  ao22d1_hd U1908 ( .A(z_m[23]), .B(n378), .C(n476), .D(n177), .Y(n172) );
  ao22d1_hd U1909 ( .A(n100), .B(n618), .C(b_m[23]), .D(n102), .Y(n173) );
  nr2d1_hd U1910 ( .A(n476), .B(o_Z_STB), .Y(n179) );
  ao22d1_hd U1911 ( .A(n1137), .B(n1136), .C(n1135), .D(n1134), .Y(n1138) );
  nr2d1_hd U1912 ( .A(n1138), .B(n1143), .Y(n1180) );
  ao22d1_hd U1913 ( .A(n1139), .B(N35), .C(n1179), .D(z_s), .Y(n1140) );
  nr2d1_hd U1914 ( .A(z_e[1]), .B(z_e[0]), .Y(n1172) );
  ivd1_hd U1915 ( .A(z_e[2]), .Y(n1168) );
  nr2d1_hd U1916 ( .A(z_e[3]), .B(n1167), .Y(n1164) );
  ivd1_hd U1917 ( .A(z_e[4]), .Y(n1161) );
  nr2d1_hd U1918 ( .A(z_e[5]), .B(n1160), .Y(n1157) );
  ivd1_hd U1919 ( .A(z_e[6]), .Y(n1154) );
  nr2d1_hd U1920 ( .A(z_m[23]), .B(z_e[0]), .Y(n1150) );
  ivd1_hd U1921 ( .A(z_e[1]), .Y(n1147) );
  nr4d1_hd U1922 ( .A(z_e[2]), .B(n1147), .C(n1146), .D(n1145), .Y(n1149) );
  ao21d1_hd U1923 ( .A(n1150), .B(n1149), .C(n1148), .Y(n1170) );
  oa211d1_hd U1924 ( .A(z_e[7]), .B(n1153), .C(n1170), .D(n1151), .Y(n1152) );
  scg15d1_hd U1925 ( .A(n1183), .B(z[30]), .C(n1176), .D(n1152), .Y(n230) );
  oa21d1_hd U1926 ( .A(n1157), .B(n1154), .C(n1153), .Y(n1155) );
  ao22d1_hd U1927 ( .A(n451), .B(z[29]), .C(n1170), .D(n1155), .Y(n1156) );
  ao21d1_hd U1928 ( .A(z_e[5]), .B(n1160), .C(n1157), .Y(n1159) );
  oa211d1_hd U1929 ( .A(n1159), .B(n1177), .C(n1176), .D(n1158), .Y(n232) );
  oa21d1_hd U1930 ( .A(n1164), .B(n1161), .C(n1160), .Y(n1162) );
  ao22d1_hd U1931 ( .A(n451), .B(z[27]), .C(n1170), .D(n1162), .Y(n1163) );
  ao21d1_hd U1932 ( .A(z_e[3]), .B(n1167), .C(n1164), .Y(n1166) );
  oa211d1_hd U1933 ( .A(n1166), .B(n1177), .C(n1176), .D(n1165), .Y(n234) );
  oa21d1_hd U1934 ( .A(n1172), .B(n1168), .C(n1167), .Y(n1169) );
  ao22d1_hd U1935 ( .A(n450), .B(z[25]), .C(n1170), .D(n1169), .Y(n1171) );
  ao21d1_hd U1936 ( .A(z_e[0]), .B(z_e[1]), .C(n1172), .Y(n1174) );
  oa211d1_hd U1937 ( .A(n1174), .B(n1177), .C(n1176), .D(n1173), .Y(n236) );
  oa211d1_hd U1938 ( .A(z_e[0]), .B(n1177), .C(n1176), .D(n1175), .Y(n237) );
  ao21d1_hd U1939 ( .A(n450), .B(z[22]), .C(n1180), .Y(n1181) );
  oa21d1_hd U1940 ( .A(n1311), .B(n1182), .C(n1181), .Y(n238) );
  nr2d1_hd U1941 ( .A(sticky), .B(round_bit), .Y(n1184) );
  nd3d1_hd U1942 ( .A(n1274), .B(z_m[4]), .C(z_m[3]), .Y(n1262) );
  ivd1_hd U1943 ( .A(n1262), .Y(n1263) );
  ivd1_hd U1944 ( .A(z_m[5]), .Y(n1266) );
  nd3d1_hd U1945 ( .A(n1254), .B(z_m[8]), .C(z_m[7]), .Y(n1244) );
  ivd1_hd U1946 ( .A(n1244), .Y(n1245) );
  ivd1_hd U1947 ( .A(z_m[9]), .Y(n1248) );
  nd3d1_hd U1948 ( .A(n1237), .B(z_m[12]), .C(n19), .Y(n1226) );
  ivd1_hd U1949 ( .A(n1226), .Y(n1228) );
  nd3d1_hd U1950 ( .A(n1228), .B(z_m[14]), .C(z_m[13]), .Y(n1217) );
  ivd1_hd U1951 ( .A(n1217), .Y(n1218) );
  nd3d1_hd U1952 ( .A(n1218), .B(z_m[16]), .C(n21), .Y(n1200) );
  ivd1_hd U1953 ( .A(n1200), .Y(n1201) );
  nd3d1_hd U1954 ( .A(n1201), .B(z_m[18]), .C(z_m[17]), .Y(n1191) );
  ivd1_hd U1955 ( .A(n1191), .Y(n1192) );
  nd3d1_hd U1956 ( .A(n1192), .B(z_m[20]), .C(n23), .Y(n1309) );
  ao21d1_hd U1957 ( .A(n201), .B(n1309), .C(n93), .Y(n1187) );
  oa21d1_hd U1958 ( .A(z_m[21]), .B(n96), .C(n1187), .Y(n1306) );
  nd2bd1_hd U1959 ( .AN(n1309), .B(n201), .Y(n1186) );
  oa21d1_hd U1960 ( .A(z_m[22]), .B(n1186), .C(n198), .Y(n1185) );
  scg4d1_hd U1961 ( .A(n1306), .B(z_m[22]), .C(n1185), .D(z_m[21]), .E(z_m[23]), .F(n1295), .G(n457), .H(product[48]), .Y(n261) );
  ivd1_hd U1962 ( .A(z_m[21]), .Y(n1310) );
  ao22d1_hd U1963 ( .A(z_m[21]), .B(n1187), .C(n1186), .D(n1310), .Y(n1190) );
  ao22d1_hd U1964 ( .A(n455), .B(product[47]), .C(z_m[22]), .D(n188), .Y(n1189) );
  oa21d1_hd U1965 ( .A(n94), .B(n1191), .C(n1261), .Y(n1195) );
  oa21d1_hd U1966 ( .A(n23), .B(n95), .C(n1195), .Y(n1194) );
  oa21d1_hd U1967 ( .A(z_m[20]), .B(n1199), .C(n198), .Y(n1193) );
  scg4d1_hd U1968 ( .A(n1194), .B(z_m[20]), .C(n1193), .D(z_m[19]), .E(z_m[21]), .F(n188), .G(n1308), .H(product[46]), .Y(n263) );
  ao22d1_hd U1969 ( .A(n455), .B(product[45]), .C(z_m[20]), .D(n187), .Y(n1198) );
  ivd1_hd U1970 ( .A(n1195), .Y(n1196) );
  ao22d1_hd U1971 ( .A(z_m[18]), .B(n97), .C(n23), .D(n1196), .Y(n1197) );
  oa211d1_hd U1972 ( .A(n23), .B(n1199), .C(n1198), .D(n1197), .Y(n264) );
  ao21d1_hd U1973 ( .A(n1227), .B(n1200), .C(n93), .Y(n1214) );
  oa21d1_hd U1974 ( .A(z_m[17]), .B(n96), .C(n1214), .Y(n1203) );
  oa21d1_hd U1975 ( .A(z_m[18]), .B(n1205), .C(n199), .Y(n1202) );
  scg4d1_hd U1976 ( .A(n1203), .B(z_m[18]), .C(n1202), .D(n193), .E(n23), .F(
        n186), .G(n1308), .H(product[44]), .Y(n265) );
  ivd1_hd U1977 ( .A(z_m[17]), .Y(n1204) );
  ao22d1_hd U1978 ( .A(z_m[17]), .B(n1214), .C(n1205), .D(n1204), .Y(n1216) );
  ao22d1_hd U1979 ( .A(n456), .B(product[43]), .C(z_m[18]), .D(n187), .Y(n1215) );
  oa21d1_hd U1980 ( .A(n93), .B(n1217), .C(n1261), .Y(n1221) );
  oa21d1_hd U1981 ( .A(n21), .B(n96), .C(n1221), .Y(n1220) );
  oa21d1_hd U1982 ( .A(z_m[16]), .B(n1225), .C(n199), .Y(n1219) );
  scg4d1_hd U1983 ( .A(n1220), .B(z_m[16]), .C(n1219), .D(z_m[15]), .E(n193), 
        .F(n187), .G(n454), .H(product[42]), .Y(n267) );
  ao22d1_hd U1984 ( .A(n456), .B(product[41]), .C(z_m[16]), .D(n186), .Y(n1224) );
  ivd1_hd U1985 ( .A(n1221), .Y(n1222) );
  ao22d1_hd U1986 ( .A(z_m[14]), .B(n98), .C(n21), .D(n1222), .Y(n1223) );
  oa211d1_hd U1987 ( .A(n21), .B(n1225), .C(n1224), .D(n1223), .Y(n268) );
  ao21d1_hd U1988 ( .A(n1227), .B(n1226), .C(n94), .Y(n1233) );
  oa21d1_hd U1989 ( .A(z_m[13]), .B(n95), .C(n1233), .Y(n1230) );
  oa21d1_hd U1990 ( .A(z_m[14]), .B(n1232), .C(n198), .Y(n1229) );
  scg4d1_hd U1991 ( .A(n1230), .B(z_m[14]), .C(n1229), .D(n192), .E(n21), .F(
        n189), .G(n454), .H(product[40]), .Y(n269) );
  ivd1_hd U1992 ( .A(z_m[13]), .Y(n1231) );
  ao22d1_hd U1993 ( .A(z_m[13]), .B(n1233), .C(n1232), .D(n1231), .Y(n1235) );
  ao22d1_hd U1994 ( .A(n455), .B(product[39]), .C(z_m[14]), .D(n186), .Y(n1234) );
  oa21d1_hd U1995 ( .A(n1272), .B(n1237), .C(n1271), .Y(n1240) );
  ivd1_hd U1996 ( .A(n1240), .Y(n1236) );
  oa21d1_hd U1997 ( .A(n19), .B(n95), .C(n1236), .Y(n1239) );
  oa21d1_hd U1998 ( .A(z_m[12]), .B(n1243), .C(n199), .Y(n1238) );
  scg4d1_hd U1999 ( .A(n1239), .B(z_m[12]), .C(n1238), .D(z_m[11]), .E(n192), 
        .F(n186), .G(n454), .H(product[38]), .Y(n271) );
  ao22d1_hd U2000 ( .A(n456), .B(product[37]), .C(z_m[12]), .D(n188), .Y(n1242) );
  ao22d1_hd U2001 ( .A(z_m[10]), .B(n97), .C(n19), .D(n1240), .Y(n1241) );
  oa211d1_hd U2002 ( .A(n19), .B(n1243), .C(n1242), .D(n1241), .Y(n272) );
  oa21d1_hd U2003 ( .A(n94), .B(n1244), .C(n1261), .Y(n1250) );
  oa21d1_hd U2004 ( .A(z_m[9]), .B(n96), .C(n1250), .Y(n1247) );
  oa21d1_hd U2005 ( .A(z_m[10]), .B(n1249), .C(n199), .Y(n1246) );
  scg4d1_hd U2006 ( .A(n1247), .B(z_m[10]), .C(n1246), .D(z_m[9]), .E(n19), 
        .F(n186), .G(n1308), .H(product[36]), .Y(n273) );
  ao22d1_hd U2007 ( .A(z_m[9]), .B(n1250), .C(n1249), .D(n1248), .Y(n1252) );
  ao22d1_hd U2008 ( .A(n457), .B(product[35]), .C(z_m[10]), .D(n189), .Y(n1251) );
  oa21d1_hd U2009 ( .A(n1272), .B(n1254), .C(n1271), .Y(n1257) );
  ivd1_hd U2010 ( .A(n1257), .Y(n1253) );
  oa21d1_hd U2011 ( .A(z_m[7]), .B(n95), .C(n1253), .Y(n1256) );
  oa21d1_hd U2012 ( .A(z_m[8]), .B(n1260), .C(n198), .Y(n1255) );
  scg4d1_hd U2013 ( .A(n1256), .B(z_m[8]), .C(n1255), .D(z_m[7]), .E(z_m[9]), 
        .F(n189), .G(n454), .H(product[34]), .Y(n275) );
  ao22d1_hd U2014 ( .A(n456), .B(product[33]), .C(z_m[8]), .D(n189), .Y(n1259)
         );
  ao22d1_hd U2015 ( .A(z_m[6]), .B(n97), .C(z_m[7]), .D(n1257), .Y(n1258) );
  oa211d1_hd U2016 ( .A(n190), .B(n1260), .C(n1259), .D(n1258), .Y(n276) );
  oa21d1_hd U2017 ( .A(n93), .B(n1262), .C(n1261), .Y(n1268) );
  oa21d1_hd U2018 ( .A(z_m[5]), .B(n96), .C(n1268), .Y(n1265) );
  oa21d1_hd U2019 ( .A(z_m[6]), .B(n1267), .C(n198), .Y(n1264) );
  scg4d1_hd U2020 ( .A(n1265), .B(z_m[6]), .C(n1264), .D(z_m[5]), .E(n190), 
        .F(n188), .G(n1308), .H(product[32]), .Y(n277) );
  ao22d1_hd U2021 ( .A(z_m[5]), .B(n1268), .C(n1267), .D(n1266), .Y(n1270) );
  ao22d1_hd U2022 ( .A(n457), .B(product[31]), .C(z_m[6]), .D(n188), .Y(n1269)
         );
  oa21d1_hd U2023 ( .A(n1272), .B(n1274), .C(n1271), .Y(n1277) );
  ivd1_hd U2024 ( .A(n1277), .Y(n1273) );
  oa21d1_hd U2025 ( .A(z_m[3]), .B(n95), .C(n1273), .Y(n1276) );
  oa21d1_hd U2026 ( .A(z_m[4]), .B(n1280), .C(n199), .Y(n1275) );
  scg4d1_hd U2027 ( .A(n1276), .B(z_m[4]), .C(n1275), .D(z_m[3]), .E(z_m[5]), 
        .F(n187), .G(n457), .H(product[30]), .Y(n279) );
  ao22d1_hd U2028 ( .A(n456), .B(product[29]), .C(z_m[4]), .D(n187), .Y(n1279)
         );
  ao22d1_hd U2029 ( .A(z_m[2]), .B(n98), .C(z_m[3]), .D(n1277), .Y(n1278) );
  oa211d1_hd U2030 ( .A(n191), .B(n1280), .C(n1279), .D(n1278), .Y(n280) );
  nr2d1_hd U2031 ( .A(n25), .B(n95), .Y(n1302) );
  nr2d1_hd U2032 ( .A(n94), .B(n1302), .Y(n1286) );
  nd2bd1_hd U2033 ( .AN(z_m[1]), .B(n200), .Y(n1285) );
  nd3bd1_hd U2034 ( .AN(z_m[2]), .B(n201), .C(n25), .Y(n1282) );
  scg4d1_hd U2035 ( .A(n1284), .B(z_m[2]), .C(n1283), .D(z_m[1]), .E(n191), 
        .F(n187), .G(n457), .H(product[28]), .Y(n281) );
  ivd1_hd U2036 ( .A(n1286), .Y(n1287) );
  scg4d1_hd U2037 ( .A(n1288), .B(n25), .C(n1287), .D(z_m[1]), .E(z_m[2]), .F(
        n189), .G(n457), .H(product[27]), .Y(n282) );
  nr4d1_hd U2038 ( .A(product[14]), .B(product[12]), .C(product[19]), .D(
        product[17]), .Y(n1292) );
  nr4d1_hd U2039 ( .A(product[15]), .B(product[8]), .C(product[20]), .D(
        product[4]), .Y(n1291) );
  nr4d1_hd U2040 ( .A(product[21]), .B(product[2]), .C(product[13]), .D(
        product[16]), .Y(n1290) );
  nr4d1_hd U2041 ( .A(product[23]), .B(product[5]), .C(product[22]), .D(
        product[18]), .Y(n1289) );
  nd4d1_hd U2042 ( .A(n1292), .B(n1291), .C(n1290), .D(n1289), .Y(n1293) );
  nr4d1_hd U2043 ( .A(product[9]), .B(product[7]), .C(n1294), .D(n1293), .Y(
        n1298) );
  ao22d1_hd U2044 ( .A(round_bit), .B(n1295), .C(sticky), .D(n1297), .Y(n1296)
         );
  oa21d1_hd U2045 ( .A(n1298), .B(n1297), .C(n1296), .Y(n283) );
  ao22d1_hd U2046 ( .A(n455), .B(product[24]), .C(round_bit), .D(n1299), .Y(
        n1300) );
  scg16d1_hd U2047 ( .A(n188), .B(net908), .C(n1300), .Y(n284) );
  ao22d1_hd U2048 ( .A(n455), .B(product[26]), .C(z_m[1]), .D(n186), .Y(n1304)
         );
  ao21d1_hd U2049 ( .A(n93), .B(z_m[0]), .C(n1302), .Y(n1303) );
  oa211d1_hd U2050 ( .A(net908), .B(n198), .C(n1304), .D(n1303), .Y(n285) );
  ao21d1_hd U2051 ( .A(n1281), .B(n1311), .C(n1306), .Y(n1316) );
  ao22d1_hd U2052 ( .A(n456), .B(product[49]), .C(z_m[22]), .D(n98), .Y(n1314)
         );
  nr3d1_hd U2053 ( .A(n1311), .B(n1310), .C(n1309), .Y(n1423) );
  nd3d1_hd U2054 ( .A(n200), .B(n1423), .C(n1315), .Y(n1313) );
  oa211d1_hd U2055 ( .A(n1316), .B(n1315), .C(n1314), .D(n1313), .Y(n286) );
  ao22d1_hd U2056 ( .A(n482), .B(b[22]), .C(intadd_23_A_17_), .D(n129), .Y(
        n1317) );
  oa21d1_hd U2057 ( .A(n600), .B(n112), .C(n1317), .Y(n287) );
  ao22d1_hd U2058 ( .A(n481), .B(b[20]), .C(intadd_23_B_16_), .D(n131), .Y(
        n1318) );
  ao22d1_hd U2059 ( .A(n481), .B(b[19]), .C(intadd_23_B_15_), .D(n130), .Y(
        n1319) );
  oa21d1_hd U2060 ( .A(n584), .B(n111), .C(n1319), .Y(n289) );
  ao22d1_hd U2061 ( .A(n481), .B(b[18]), .C(intadd_23_B_14_), .D(n130), .Y(
        n1320) );
  ao22d1_hd U2062 ( .A(n481), .B(b[17]), .C(intadd_23_B_13_), .D(n129), .Y(
        n1321) );
  ao22d1_hd U2063 ( .A(n481), .B(b[16]), .C(intadd_23_B_12_), .D(n129), .Y(
        n1322) );
  oa21d1_hd U2064 ( .A(n572), .B(n110), .C(n1322), .Y(n292) );
  ao22d1_hd U2065 ( .A(n480), .B(b[15]), .C(intadd_23_B_11_), .D(n132), .Y(
        n1323) );
  oa21d1_hd U2066 ( .A(n567), .B(n112), .C(n1323), .Y(n293) );
  ao22d1_hd U2067 ( .A(n480), .B(b[14]), .C(intadd_23_B_10_), .D(n132), .Y(
        n1324) );
  ao22d1_hd U2068 ( .A(n480), .B(b[13]), .C(intadd_23_B_9_), .D(n131), .Y(
        n1325) );
  oa21d1_hd U2069 ( .A(n558), .B(n111), .C(n1325), .Y(n295) );
  ao22d1_hd U2070 ( .A(n480), .B(b[12]), .C(intadd_23_B_8_), .D(n132), .Y(
        n1326) );
  ao22d1_hd U2071 ( .A(n480), .B(b[11]), .C(intadd_23_B_7_), .D(n130), .Y(
        n1327) );
  oa21d1_hd U2072 ( .A(n549), .B(n110), .C(n1327), .Y(n297) );
  ao22d1_hd U2073 ( .A(n480), .B(b[10]), .C(intadd_23_B_6_), .D(n129), .Y(
        n1328) );
  oa21d1_hd U2074 ( .A(n544), .B(n112), .C(n1328), .Y(n298) );
  ao22d1_hd U2075 ( .A(n479), .B(b[9]), .C(intadd_23_B_5_), .D(n132), .Y(n1329) );
  oa21d1_hd U2076 ( .A(n539), .B(n111), .C(n1329), .Y(n299) );
  ao22d1_hd U2077 ( .A(n479), .B(b[8]), .C(intadd_23_B_4_), .D(n131), .Y(n1330) );
  ao22d1_hd U2078 ( .A(n479), .B(b[7]), .C(intadd_23_B_3_), .D(n131), .Y(n1331) );
  oa21d1_hd U2079 ( .A(n529), .B(n110), .C(n1331), .Y(n301) );
  ao22d1_hd U2080 ( .A(n479), .B(b[6]), .C(intadd_23_B_2_), .D(n130), .Y(n1333) );
  ao22d1_hd U2081 ( .A(n479), .B(b[5]), .C(intadd_23_B_1_), .D(n129), .Y(n1334) );
  ao22d1_hd U2082 ( .A(n478), .B(b[4]), .C(intadd_23_B_0_), .D(n130), .Y(n1335) );
  oa21d1_hd U2083 ( .A(n517), .B(n112), .C(n1335), .Y(n304) );
  ao22d1_hd U2084 ( .A(n478), .B(b[3]), .C(n502), .D(n129), .Y(n1336) );
  oa21d1_hd U2085 ( .A(n513), .B(n111), .C(n1336), .Y(n305) );
  ao22d1_hd U2086 ( .A(n478), .B(b[2]), .C(n180), .D(n132), .Y(n1337) );
  oa21d1_hd U2087 ( .A(n507), .B(n110), .C(n1337), .Y(n306) );
  ao22d1_hd U2088 ( .A(n478), .B(b[1]), .C(n123), .D(n131), .Y(n1338) );
  oa21d1_hd U2089 ( .A(n197), .B(n112), .C(n1338), .Y(n307) );
  ao22d1_hd U2090 ( .A(n478), .B(b[21]), .C(intadd_23_B_17_), .D(n130), .Y(
        n1342) );
  oa21d1_hd U2091 ( .A(n594), .B(n111), .C(n1342), .Y(n309) );
  ivd1_hd U2092 ( .A(n1344), .Y(n1414) );
  ao22d1_hd U2093 ( .A(n102), .B(n596), .C(n1117), .D(n116), .Y(n1345) );
  oa21d1_hd U2094 ( .A(n1346), .B(n1414), .C(n1345), .Y(n310) );
  oa211d1_hd U2095 ( .A(n1356), .B(n1348), .C(n1363), .D(n1347), .Y(n1350) );
  ao211d1_hd U2096 ( .A(a_e[8]), .B(n100), .C(DP_OP_113J2_124_6892_n3), .D(
        n1349), .Y(n1360) );
  ao22d1_hd U2097 ( .A(a_e[8]), .B(n1350), .C(n1360), .D(n195), .Y(n1351) );
  ao22d1_hd U2098 ( .A(a_e[1]), .B(n69), .C(C81_DATA2_1), .D(n1358), .Y(n1353)
         );
  oa22d1_hd U2099 ( .A(n1355), .B(n1206), .C(n1354), .D(n1363), .Y(n318) );
  nr2d1_hd U2100 ( .A(n1356), .B(n1362), .Y(n1359) );
  oa211d1_hd U2101 ( .A(n1360), .B(n1359), .C(n1358), .D(n1357), .Y(n1361) );
  oa211d1_hd U2102 ( .A(n1363), .B(n1362), .C(n138), .D(n1361), .Y(n319) );
  ivd1_hd U2103 ( .A(n1364), .Y(n1366) );
  nr2d1_hd U2104 ( .A(DP_OP_116J2_127_7148_n3), .B(n1366), .Y(n1365) );
  oa21d1_hd U2105 ( .A(n1365), .B(n1416), .C(n1370), .Y(n1367) );
  ao211d1_hd U2106 ( .A(n101), .B(b_e[8]), .C(DP_OP_116J2_127_7148_n3), .D(
        n1366), .Y(n1420) );
  ao22d1_hd U2107 ( .A(b_e[8]), .B(n1367), .C(n1420), .D(n1418), .Y(n1368) );
  ao22d1_hd U2108 ( .A(b_e[1]), .B(n79), .C(C82_DATA2_1), .D(n1418), .Y(n1369)
         );
  ao22d1_hd U2109 ( .A(n478), .B(a[21]), .C(n205), .D(a_m[21]), .Y(n1372) );
  oa21d1_hd U2110 ( .A(n224), .B(n113), .C(n1372), .Y(n328) );
  ao22d1_hd U2111 ( .A(n477), .B(a[20]), .C(n202), .D(n120), .Y(n1373) );
  oa21d1_hd U2112 ( .A(n222), .B(n1374), .C(n1373), .Y(n329) );
  ao22d1_hd U2113 ( .A(n477), .B(a[19]), .C(n202), .D(a_m[19]), .Y(n1375) );
  oa21d1_hd U2114 ( .A(n225), .B(n1376), .C(n1375), .Y(n330) );
  oa22d1_hd U2115 ( .A(n223), .B(n459), .C(n1392), .D(n1376), .Y(n331) );
  ao22d1_hd U2116 ( .A(n479), .B(a[17]), .C(n204), .D(n92), .Y(n1378) );
  oa21d1_hd U2117 ( .A(n223), .B(n1379), .C(n1378), .Y(n332) );
  ao22d1_hd U2118 ( .A(n477), .B(a[16]), .C(n203), .D(a_m[16]), .Y(n1380) );
  oa21d1_hd U2119 ( .A(n224), .B(n1381), .C(n1380), .Y(n333) );
  oa22d1_hd U2120 ( .A(n224), .B(n462), .C(n1392), .D(n1381), .Y(n334) );
  ao22d1_hd U2121 ( .A(n477), .B(a[14]), .C(n204), .D(a_m[14]), .Y(n1383) );
  oa21d1_hd U2122 ( .A(n225), .B(n1384), .C(n1383), .Y(n335) );
  ao22d1_hd U2123 ( .A(n477), .B(a[13]), .C(n205), .D(a_m[13]), .Y(n1385) );
  oa21d1_hd U2124 ( .A(n223), .B(n1386), .C(n1385), .Y(n336) );
  oa22d1_hd U2125 ( .A(n225), .B(n466), .C(n1392), .D(n1386), .Y(n337) );
  ao22d1_hd U2126 ( .A(n1332), .B(a[11]), .C(n202), .D(a_m[11]), .Y(n1388) );
  oa21d1_hd U2127 ( .A(n224), .B(n1389), .C(n1388), .Y(n338) );
  ao22d1_hd U2128 ( .A(n487), .B(a[10]), .C(n203), .D(a_m[10]), .Y(n1390) );
  oa21d1_hd U2129 ( .A(n225), .B(n1391), .C(n1390), .Y(n339) );
  oa22d1_hd U2130 ( .A(n223), .B(n606), .C(n1392), .D(n1391), .Y(n340) );
  ao22d1_hd U2131 ( .A(n487), .B(a[8]), .C(n204), .D(n602), .Y(n1393) );
  oa21d1_hd U2132 ( .A(n223), .B(n1394), .C(n1393), .Y(n341) );
  ao22d1_hd U2133 ( .A(n487), .B(a[7]), .C(n205), .D(a_m[7]), .Y(n1395) );
  oa21d1_hd U2134 ( .A(n224), .B(n1396), .C(n1395), .Y(n342) );
  ao22d1_hd U2135 ( .A(n487), .B(a[6]), .C(n202), .D(a_m[6]), .Y(n1397) );
  oa21d1_hd U2136 ( .A(n225), .B(n470), .C(n1397), .Y(n343) );
  ao22d1_hd U2137 ( .A(n1332), .B(a[5]), .C(n203), .D(n82), .Y(n1399) );
  oa21d1_hd U2138 ( .A(n222), .B(n1400), .C(n1399), .Y(n344) );
  ao22d1_hd U2139 ( .A(n485), .B(a[4]), .C(n203), .D(a_m[4]), .Y(n1401) );
  oa21d1_hd U2140 ( .A(n223), .B(n1402), .C(n1401), .Y(n345) );
  ao22d1_hd U2141 ( .A(n486), .B(a[3]), .C(n204), .D(a_m[3]), .Y(n1403) );
  oa21d1_hd U2142 ( .A(n224), .B(n473), .C(n1403), .Y(n346) );
  ao22d1_hd U2143 ( .A(n477), .B(a[2]), .C(n203), .D(n106), .Y(n1405) );
  oa21d1_hd U2144 ( .A(n222), .B(n1406), .C(n1405), .Y(n347) );
  ao22d1_hd U2145 ( .A(n486), .B(a[1]), .C(n205), .D(a_m[1]), .Y(n1407) );
  oa21d1_hd U2146 ( .A(n225), .B(n1408), .C(n1407), .Y(n348) );
  ao22d1_hd U2147 ( .A(n486), .B(a[22]), .C(n202), .D(a_m[22]), .Y(n1410) );
  oa21d1_hd U2148 ( .A(n222), .B(n1411), .C(n1410), .Y(n354) );
  ao22d1_hd U2149 ( .A(a_m[22]), .B(n100), .C(n618), .D(n117), .Y(n1413) );
  oa21d1_hd U2150 ( .A(n1415), .B(n1414), .C(n1413), .Y(n355) );
  nr2d1_hd U2151 ( .A(n1422), .B(n1416), .Y(n1419) );
  oa211d1_hd U2152 ( .A(n1420), .B(n1419), .C(n1418), .D(n1417), .Y(n1421) );
  oa211d1_hd U2153 ( .A(n1370), .B(n1422), .C(n148), .D(n1421), .Y(n356) );
  ivd1_hd U2154 ( .A(state[3]), .Y(n1435) );
  ivd1_hd U2155 ( .A(n1429), .Y(n1436) );
  ivd1_hd U2156 ( .A(o_AB_ACK), .Y(n1437) );
endmodule


module iir_lpf ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   r_add_AB_STB, w_add_AB_ACK, w_add_Z_STB, r_add_Z_ACK, w_mult_1_AB_ACK,
         w_mult_2_AB_ACK, w_mult_1_Z_STB, w_mult_2_Z_STB, r_mult_AB_STB,
         r_mult_Z_ACK, N18, r_pstate_0_, N807, N814, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n207, n252, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097;
  wire   [31:0] r_add_A;
  wire   [31:0] r_add_B;
  wire   [31:0] w_add_Z;
  wire   [29:0] r_mult_1_A;
  wire   [31:0] r_mult_1_B;
  wire   [31:0] w_mult_1_Z;
  wire   [31:0] r_mult_2_A;
  wire   [31:0] r_mult_2_B;
  wire   [31:0] w_mult_2_Z;
  wire   [95:0] r_x_data;
  wire   [63:0] r_y_data;

  float_adder add ( .i_A(r_add_A), .i_B(r_add_B), .i_AB_STB(r_add_AB_STB), 
        .o_AB_ACK(w_add_AB_ACK), .o_Z(w_add_Z), .o_Z_STB(w_add_Z_STB), 
        .i_Z_ACK(r_add_Z_ACK), .i_CLK(i_CLK), .i_RST(N18) );
  float_multiplier_1 mult_1 ( .i_A({1'b0, 1'b0, r_mult_1_A[29:22], 1'b0, 
        r_mult_1_A[20:19], 1'b0, r_mult_1_A[17:14], 1'b0, r_mult_1_A[12:0]}), 
        .i_B(r_mult_1_B), .i_AB_STB(r_mult_AB_STB), .o_AB_ACK(w_mult_1_AB_ACK), 
        .o_Z(w_mult_1_Z), .o_Z_STB(w_mult_1_Z_STB), .i_Z_ACK(r_mult_Z_ACK), 
        .i_CLK(i_CLK), .i_RST(N18) );
  float_multiplier_0 mult_2 ( .i_A({r_mult_2_A[31], 1'b0, r_mult_2_A[29:24], 
        1'b0, r_mult_2_A[22:19], 1'b0, r_mult_2_A[17:16], 1'b0, 
        r_mult_2_A[14:13], 1'b0, r_mult_2_A[11:10], 1'b0, r_mult_2_A[8:0]}), 
        .i_B(r_mult_2_B), .i_AB_STB(r_mult_AB_STB), .o_AB_ACK(w_mult_2_AB_ACK), 
        .o_Z(w_mult_2_Z), .o_Z_STB(w_mult_2_Z_STB), .i_Z_ACK(r_mult_Z_ACK), 
        .i_CLK(i_CLK), .i_RST(N18) );
  fd3qd1_hd r_counter_reg_0_ ( .D(n163), .CK(i_CLK), .SN(i_RSTN), .Q(n164) );
  fd3qd1_hd r_counter_reg_1_ ( .D(n162), .CK(i_CLK), .SN(i_RSTN), .Q(n207) );
  fd3qd1_hd r_pstate_reg_1_ ( .D(n160), .CK(i_CLK), .SN(i_RSTN), .Q(n161) );
  nr2d1_hd U555 ( .A(n252), .B(N18), .Y(N814) );
  ivd1_hd U574 ( .A(i_RSTN), .Y(N18) );
  fd2qd1_hd r_mult_2_A_reg_22_ ( .D(n389), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[22]) );
  fd2qd1_hd r_mult_2_A_reg_19_ ( .D(n392), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[19]) );
  fd2qd1_hd r_mult_2_A_reg_2_ ( .D(n405), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[2]) );
  fd2qd1_hd r_mult_2_A_reg_1_ ( .D(n406), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_19_ ( .D(n417), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[19]) );
  fd2qd1_hd r_mult_1_A_reg_16_ ( .D(n419), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[16]) );
  fd2qd1_hd r_mult_1_A_reg_2_ ( .D(n432), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[2]) );
  fd2qd1_hd r_mult_1_A_reg_1_ ( .D(n433), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_0_ ( .D(n434), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[0]) );
  fd2qd1_hd r_mult_2_A_reg_31_ ( .D(n382), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[31]) );
  fd2qd1_hd r_mult_2_A_reg_25_ ( .D(n387), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[25]) );
  fd2qd1_hd r_mult_2_A_reg_24_ ( .D(n388), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[24]) );
  fd2qd1_hd r_mult_2_A_reg_21_ ( .D(n390), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[21]) );
  fd2qd1_hd r_mult_2_A_reg_14_ ( .D(n395), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[14]) );
  fd2qd1_hd r_mult_2_A_reg_13_ ( .D(n396), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[13]) );
  fd2qd1_hd r_mult_2_A_reg_8_ ( .D(n399), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[8]) );
  fd2qd1_hd r_mult_2_A_reg_4_ ( .D(n403), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[4]) );
  fd2qd1_hd r_mult_1_A_reg_25_ ( .D(n412), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[25]) );
  fd2qd1_hd r_mult_1_A_reg_24_ ( .D(n413), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[24]) );
  fd2qd1_hd r_mult_1_A_reg_15_ ( .D(n420), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[15]) );
  fd2qd1_hd r_mult_1_A_reg_14_ ( .D(n421), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[14]) );
  fd2qd1_hd r_mult_1_A_reg_12_ ( .D(n422), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[12]) );
  fd2qd1_hd r_mult_1_A_reg_9_ ( .D(n425), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[9]) );
  fd2qd1_hd r_mult_1_A_reg_8_ ( .D(n426), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[8]) );
  fd2qd1_hd r_mult_1_A_reg_4_ ( .D(n430), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[4]) );
  fd2qd1_hd r_mult_2_A_reg_29_ ( .D(n383), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[29]) );
  fd2qd1_hd r_mult_2_A_reg_28_ ( .D(n384), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[28]) );
  fd2qd1_hd r_mult_2_A_reg_27_ ( .D(n385), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[27]) );
  fd2qd1_hd r_mult_2_A_reg_26_ ( .D(n386), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[26]) );
  fd2qd1_hd r_mult_2_A_reg_20_ ( .D(n391), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[20]) );
  fd2qd1_hd r_mult_2_A_reg_17_ ( .D(n393), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[17]) );
  fd2qd1_hd r_mult_2_A_reg_16_ ( .D(n394), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[16]) );
  fd2qd1_hd r_mult_2_A_reg_11_ ( .D(n397), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[11]) );
  fd2qd1_hd r_mult_2_A_reg_10_ ( .D(n398), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[10]) );
  fd2qd1_hd r_mult_2_A_reg_7_ ( .D(n400), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[7]) );
  fd2qd1_hd r_mult_2_A_reg_6_ ( .D(n401), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[6]) );
  fd2qd1_hd r_mult_2_A_reg_5_ ( .D(n402), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[5]) );
  fd2qd1_hd r_mult_2_A_reg_3_ ( .D(n404), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[3]) );
  fd2qd1_hd r_mult_2_A_reg_0_ ( .D(n407), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[0]) );
  fd2qd1_hd r_mult_1_A_reg_29_ ( .D(n408), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_28_ ( .D(n409), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[28]) );
  fd2qd1_hd r_mult_1_A_reg_27_ ( .D(n410), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[27]) );
  fd2qd1_hd r_mult_1_A_reg_26_ ( .D(n411), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[26]) );
  fd2qd1_hd r_mult_1_A_reg_23_ ( .D(n414), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[23]) );
  fd2qd1_hd r_mult_1_A_reg_22_ ( .D(n415), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[22]) );
  fd2qd1_hd r_mult_1_A_reg_20_ ( .D(n416), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[20]) );
  fd2qd1_hd r_mult_1_A_reg_17_ ( .D(n418), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[17]) );
  fd2qd1_hd r_mult_1_A_reg_11_ ( .D(n423), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[11]) );
  fd2qd1_hd r_mult_1_A_reg_10_ ( .D(n424), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[10]) );
  fd2qd1_hd r_mult_1_A_reg_7_ ( .D(n427), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[7]) );
  fd2qd1_hd r_mult_1_A_reg_6_ ( .D(n428), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[6]) );
  fd2qd1_hd r_mult_1_A_reg_5_ ( .D(n429), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[5]) );
  fd2qd1_hd r_mult_1_A_reg_3_ ( .D(n431), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[3]) );
  fd2qd1_hd r_add_B_reg_0_ ( .D(n380), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[0])
         );
  fd2qd1_hd r_add_B_reg_1_ ( .D(n379), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[1])
         );
  fd2qd1_hd r_add_B_reg_2_ ( .D(n378), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[2])
         );
  fd2qd1_hd r_add_B_reg_3_ ( .D(n377), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[3])
         );
  fd2qd1_hd r_add_B_reg_4_ ( .D(n376), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[4])
         );
  fd2qd1_hd r_add_B_reg_5_ ( .D(n375), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[5])
         );
  fd2qd1_hd r_add_B_reg_6_ ( .D(n374), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[6])
         );
  fd2qd1_hd r_add_B_reg_7_ ( .D(n373), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[7])
         );
  fd2qd1_hd r_add_B_reg_8_ ( .D(n372), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[8])
         );
  fd2qd1_hd r_add_B_reg_9_ ( .D(n371), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[9])
         );
  fd2qd1_hd r_add_B_reg_10_ ( .D(n370), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[10]) );
  fd2qd1_hd r_add_B_reg_11_ ( .D(n369), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[11]) );
  fd2qd1_hd r_add_B_reg_12_ ( .D(n368), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[12]) );
  fd2qd1_hd r_add_B_reg_13_ ( .D(n367), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[13]) );
  fd2qd1_hd r_add_B_reg_14_ ( .D(n366), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[14]) );
  fd2qd1_hd r_add_B_reg_15_ ( .D(n365), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[15]) );
  fd2qd1_hd r_add_B_reg_16_ ( .D(n364), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[16]) );
  fd2qd1_hd r_add_B_reg_17_ ( .D(n363), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[17]) );
  fd2qd1_hd r_add_B_reg_18_ ( .D(n362), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[18]) );
  fd2qd1_hd r_add_B_reg_19_ ( .D(n361), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[19]) );
  fd2qd1_hd r_add_B_reg_20_ ( .D(n360), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[20]) );
  fd2qd1_hd r_add_B_reg_21_ ( .D(n359), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[21]) );
  fd2qd1_hd r_add_B_reg_22_ ( .D(n358), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[22]) );
  fd2qd1_hd r_add_B_reg_23_ ( .D(n357), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[23]) );
  fd2qd1_hd r_add_B_reg_24_ ( .D(n356), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[24]) );
  fd2qd1_hd r_add_B_reg_25_ ( .D(n355), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[25]) );
  fd2qd1_hd r_add_B_reg_26_ ( .D(n354), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[26]) );
  fd2qd1_hd r_add_B_reg_27_ ( .D(n353), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[27]) );
  fd2qd1_hd r_add_B_reg_28_ ( .D(n352), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[28]) );
  fd2qd1_hd r_add_B_reg_29_ ( .D(n351), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[29]) );
  fd2qd1_hd r_add_B_reg_30_ ( .D(n350), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[30]) );
  fd2qd1_hd r_add_B_reg_31_ ( .D(n349), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[31]) );
  fd2qd1_hd r_x_data_reg_64_ ( .D(n95), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[64]) );
  fd2qd1_hd r_x_data_reg_65_ ( .D(n94), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[65]) );
  fd2qd1_hd r_x_data_reg_66_ ( .D(n93), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[66]) );
  fd2qd1_hd r_x_data_reg_67_ ( .D(n92), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[67]) );
  fd2qd1_hd r_x_data_reg_68_ ( .D(n91), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[68]) );
  fd2qd1_hd r_x_data_reg_69_ ( .D(n90), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[69]) );
  fd2qd1_hd r_x_data_reg_70_ ( .D(n89), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[70]) );
  fd2qd1_hd r_x_data_reg_71_ ( .D(n88), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[71]) );
  fd2qd1_hd r_x_data_reg_72_ ( .D(n87), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[72]) );
  fd2qd1_hd r_x_data_reg_73_ ( .D(n86), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[73]) );
  fd2qd1_hd r_x_data_reg_74_ ( .D(n85), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[74]) );
  fd2qd1_hd r_x_data_reg_75_ ( .D(n84), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[75]) );
  fd2qd1_hd r_x_data_reg_76_ ( .D(n83), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[76]) );
  fd2qd1_hd r_x_data_reg_77_ ( .D(n82), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[77]) );
  fd2qd1_hd r_x_data_reg_78_ ( .D(n81), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[78]) );
  fd2qd1_hd r_x_data_reg_79_ ( .D(n80), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[79]) );
  fd2qd1_hd r_x_data_reg_80_ ( .D(n79), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[80]) );
  fd2qd1_hd r_x_data_reg_81_ ( .D(n78), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[81]) );
  fd2qd1_hd r_x_data_reg_82_ ( .D(n77), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[82]) );
  fd2qd1_hd r_x_data_reg_83_ ( .D(n76), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[83]) );
  fd2qd1_hd r_x_data_reg_84_ ( .D(n75), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[84]) );
  fd2qd1_hd r_x_data_reg_85_ ( .D(n74), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[85]) );
  fd2qd1_hd r_x_data_reg_86_ ( .D(n73), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[86]) );
  fd2qd1_hd r_x_data_reg_87_ ( .D(n72), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[87]) );
  fd2qd1_hd r_x_data_reg_88_ ( .D(n71), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[88]) );
  fd2qd1_hd r_x_data_reg_89_ ( .D(n70), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[89]) );
  fd2qd1_hd r_x_data_reg_90_ ( .D(n69), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[90]) );
  fd2qd1_hd r_x_data_reg_91_ ( .D(n68), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[91]) );
  fd2qd1_hd r_x_data_reg_92_ ( .D(n67), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[92]) );
  fd2qd1_hd r_x_data_reg_93_ ( .D(n66), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[93]) );
  fd2qd1_hd r_x_data_reg_94_ ( .D(n65), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[94]) );
  fd2qd1_hd r_x_data_reg_95_ ( .D(n64), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[95]) );
  fd2qd1_hd r_x_data_reg_32_ ( .D(n127), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[32]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(n126), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(n125), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[34]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(n124), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(n123), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(n122), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[37]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(n121), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(n120), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(n119), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(n118), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(n117), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(n116), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(n115), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(n114), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(n113), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(n112), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(n111), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(n110), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(n109), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(n108), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[51]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(n107), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(n106), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(n105), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(n104), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(n103), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(n102), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(n101), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[58]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(n100), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(n99), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(n98), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(n97), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(n96), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[63]) );
  fd2qd1_hd r_add_A_reg_0_ ( .D(n568), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[0])
         );
  fd2qd1_hd r_mult_2_B_reg_31_ ( .D(n533), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[31]) );
  fd2qd1_hd r_mult_2_B_reg_30_ ( .D(n436), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_30_ ( .D(n467), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[30]) );
  fd2qd1_hd r_mult_2_B_reg_29_ ( .D(n437), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[29]) );
  fd2qd1_hd r_mult_1_B_reg_29_ ( .D(n468), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[29]) );
  fd2qd1_hd r_mult_2_B_reg_28_ ( .D(n438), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[28]) );
  fd2qd1_hd r_mult_1_B_reg_28_ ( .D(n469), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[28]) );
  fd2qd1_hd r_mult_2_B_reg_27_ ( .D(n439), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[27]) );
  fd2qd1_hd r_mult_1_B_reg_27_ ( .D(n470), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[27]) );
  fd2qd1_hd r_mult_2_B_reg_26_ ( .D(n440), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[26]) );
  fd2qd1_hd r_mult_1_B_reg_26_ ( .D(n471), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[26]) );
  fd2qd1_hd r_mult_2_B_reg_25_ ( .D(n441), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[25]) );
  fd2qd1_hd r_mult_1_B_reg_25_ ( .D(n472), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[25]) );
  fd2qd1_hd r_mult_2_B_reg_24_ ( .D(n442), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[24]) );
  fd2qd1_hd r_mult_1_B_reg_24_ ( .D(n473), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[24]) );
  fd2qd1_hd r_mult_2_B_reg_23_ ( .D(n443), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[23]) );
  fd2qd1_hd r_mult_1_B_reg_23_ ( .D(n474), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[23]) );
  fd2qd1_hd r_mult_2_B_reg_22_ ( .D(n444), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[22]) );
  fd2qd1_hd r_mult_1_B_reg_22_ ( .D(n475), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[22]) );
  fd2qd1_hd r_mult_2_B_reg_21_ ( .D(n445), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[21]) );
  fd2qd1_hd r_mult_1_B_reg_21_ ( .D(n476), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[21]) );
  fd2qd1_hd r_mult_2_B_reg_20_ ( .D(n446), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[20]) );
  fd2qd1_hd r_mult_1_B_reg_20_ ( .D(n477), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[20]) );
  fd2qd1_hd r_mult_2_B_reg_19_ ( .D(n447), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[19]) );
  fd2qd1_hd r_mult_1_B_reg_19_ ( .D(n478), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[19]) );
  fd2qd1_hd r_mult_2_B_reg_18_ ( .D(n448), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[18]) );
  fd2qd1_hd r_mult_1_B_reg_18_ ( .D(n479), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[18]) );
  fd2qd1_hd r_mult_2_B_reg_17_ ( .D(n449), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[17]) );
  fd2qd1_hd r_mult_1_B_reg_17_ ( .D(n480), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[17]) );
  fd2qd1_hd r_mult_2_B_reg_16_ ( .D(n450), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[16]) );
  fd2qd1_hd r_mult_1_B_reg_16_ ( .D(n481), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[16]) );
  fd2qd1_hd r_mult_2_B_reg_15_ ( .D(n451), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[15]) );
  fd2qd1_hd r_mult_1_B_reg_15_ ( .D(n482), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[15]) );
  fd2qd1_hd r_mult_2_B_reg_14_ ( .D(n452), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[14]) );
  fd2qd1_hd r_mult_1_B_reg_14_ ( .D(n483), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[14]) );
  fd2qd1_hd r_mult_2_B_reg_13_ ( .D(n453), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[13]) );
  fd2qd1_hd r_mult_1_B_reg_13_ ( .D(n484), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[13]) );
  fd2qd1_hd r_mult_2_B_reg_12_ ( .D(n454), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[12]) );
  fd2qd1_hd r_mult_1_B_reg_12_ ( .D(n485), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[12]) );
  fd2qd1_hd r_mult_2_B_reg_11_ ( .D(n455), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[11]) );
  fd2qd1_hd r_mult_1_B_reg_11_ ( .D(n486), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[11]) );
  fd2qd1_hd r_mult_2_B_reg_10_ ( .D(n456), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[10]) );
  fd2qd1_hd r_mult_1_B_reg_10_ ( .D(n487), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[10]) );
  fd2qd1_hd r_mult_2_B_reg_9_ ( .D(n457), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[9]) );
  fd2qd1_hd r_mult_1_B_reg_9_ ( .D(n488), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[9]) );
  fd2qd1_hd r_mult_2_B_reg_8_ ( .D(n458), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[8]) );
  fd2qd1_hd r_mult_1_B_reg_8_ ( .D(n489), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[8]) );
  fd2qd1_hd r_mult_2_B_reg_7_ ( .D(n459), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[7]) );
  fd2qd1_hd r_mult_1_B_reg_7_ ( .D(n490), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[7]) );
  fd2qd1_hd r_mult_2_B_reg_6_ ( .D(n460), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[6]) );
  fd2qd1_hd r_mult_1_B_reg_6_ ( .D(n491), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[6]) );
  fd2qd1_hd r_mult_2_B_reg_5_ ( .D(n461), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[5]) );
  fd2qd1_hd r_mult_1_B_reg_5_ ( .D(n492), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[5]) );
  fd2qd1_hd r_mult_2_B_reg_4_ ( .D(n462), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[4]) );
  fd2qd1_hd r_mult_1_B_reg_4_ ( .D(n493), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[4]) );
  fd2qd1_hd r_mult_2_B_reg_3_ ( .D(n463), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[3]) );
  fd2qd1_hd r_mult_1_B_reg_3_ ( .D(n494), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[3]) );
  fd2qd1_hd r_mult_2_B_reg_2_ ( .D(n464), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[2]) );
  fd2qd1_hd r_mult_1_B_reg_2_ ( .D(n495), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[2]) );
  fd2qd1_hd r_mult_2_B_reg_1_ ( .D(n465), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[1]) );
  fd2qd1_hd r_mult_1_B_reg_1_ ( .D(n496), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[1]) );
  fd2qd1_hd r_mult_2_B_reg_0_ ( .D(n466), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[0]) );
  fd2qd1_hd r_mult_1_B_reg_0_ ( .D(n497), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[0]) );
  fd2qd1_hd r_add_A_reg_1_ ( .D(n527), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[1])
         );
  fd2qd1_hd r_add_A_reg_2_ ( .D(n526), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[2])
         );
  fd2qd1_hd r_add_A_reg_3_ ( .D(n525), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[3])
         );
  fd2qd1_hd r_add_A_reg_4_ ( .D(n524), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[4])
         );
  fd2qd1_hd r_add_A_reg_5_ ( .D(n523), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[5])
         );
  fd2qd1_hd r_add_A_reg_6_ ( .D(n522), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[6])
         );
  fd2qd1_hd r_add_A_reg_7_ ( .D(n521), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[7])
         );
  fd2qd1_hd r_add_A_reg_8_ ( .D(n520), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[8])
         );
  fd2qd1_hd r_add_A_reg_9_ ( .D(n519), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[9])
         );
  fd2qd1_hd r_add_A_reg_10_ ( .D(n518), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[10]) );
  fd2qd1_hd r_add_A_reg_11_ ( .D(n517), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[11]) );
  fd2qd1_hd r_add_A_reg_12_ ( .D(n516), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[12]) );
  fd2qd1_hd r_add_A_reg_13_ ( .D(n515), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[13]) );
  fd2qd1_hd r_add_A_reg_14_ ( .D(n514), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[14]) );
  fd2qd1_hd r_add_A_reg_15_ ( .D(n513), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[15]) );
  fd2qd1_hd r_add_A_reg_16_ ( .D(n512), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[16]) );
  fd2qd1_hd r_add_A_reg_17_ ( .D(n511), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[17]) );
  fd2qd1_hd r_add_A_reg_18_ ( .D(n510), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[18]) );
  fd2qd1_hd r_add_A_reg_19_ ( .D(n509), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[19]) );
  fd2qd1_hd r_add_A_reg_20_ ( .D(n508), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[20]) );
  fd2qd1_hd r_add_A_reg_21_ ( .D(n507), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[21]) );
  fd2qd1_hd r_add_A_reg_22_ ( .D(n506), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[22]) );
  fd2qd1_hd r_add_A_reg_23_ ( .D(n505), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[23]) );
  fd2qd1_hd r_add_A_reg_24_ ( .D(n504), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[24]) );
  fd2qd1_hd r_add_A_reg_25_ ( .D(n503), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[25]) );
  fd2qd1_hd r_add_A_reg_26_ ( .D(n502), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[26]) );
  fd2qd1_hd r_add_A_reg_27_ ( .D(n501), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[27]) );
  fd2qd1_hd r_add_A_reg_28_ ( .D(n500), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[28]) );
  fd2qd1_hd r_add_A_reg_29_ ( .D(n499), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[29]) );
  fd2qd1_hd r_add_A_reg_30_ ( .D(n498), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[30]) );
  fd2qd1_hd r_mult_1_B_reg_31_ ( .D(n565), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[31]) );
  fd2qd1_hd r_add_A_reg_31_ ( .D(n567), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[31]) );
  fd2qd1_hd r_y_data_reg_63_ ( .D(n165), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[63]) );
  fd2qd1_hd r_y_data_reg_62_ ( .D(n62), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[62]) );
  fd2qd1_hd r_y_data_reg_61_ ( .D(n60), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[61]) );
  fd2qd1_hd r_y_data_reg_60_ ( .D(n58), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[60]) );
  fd2qd1_hd r_y_data_reg_59_ ( .D(n56), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[59]) );
  fd2qd1_hd r_y_data_reg_58_ ( .D(n54), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[58]) );
  fd2qd1_hd r_y_data_reg_57_ ( .D(n52), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[57]) );
  fd2qd1_hd r_y_data_reg_56_ ( .D(n50), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[56]) );
  fd2qd1_hd r_y_data_reg_55_ ( .D(n48), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[55]) );
  fd2qd1_hd r_y_data_reg_54_ ( .D(n46), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[54]) );
  fd2qd1_hd r_y_data_reg_53_ ( .D(n44), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[53]) );
  fd2qd1_hd r_y_data_reg_52_ ( .D(n42), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[52]) );
  fd2qd1_hd r_y_data_reg_51_ ( .D(n40), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[51]) );
  fd2qd1_hd r_y_data_reg_50_ ( .D(n38), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[50]) );
  fd2qd1_hd r_y_data_reg_49_ ( .D(n36), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[49]) );
  fd2qd1_hd r_y_data_reg_48_ ( .D(n34), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[48]) );
  fd2qd1_hd r_y_data_reg_47_ ( .D(n32), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[47]) );
  fd2qd1_hd r_y_data_reg_46_ ( .D(n30), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[46]) );
  fd2qd1_hd r_y_data_reg_45_ ( .D(n28), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[45]) );
  fd2qd1_hd r_y_data_reg_44_ ( .D(n26), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[44]) );
  fd2qd1_hd r_y_data_reg_43_ ( .D(n24), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[43]) );
  fd2qd1_hd r_y_data_reg_42_ ( .D(n22), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[42]) );
  fd2qd1_hd r_y_data_reg_41_ ( .D(n20), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[41]) );
  fd2qd1_hd r_y_data_reg_40_ ( .D(n18), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[40]) );
  fd2qd1_hd r_y_data_reg_39_ ( .D(n16), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[39]) );
  fd2qd1_hd r_y_data_reg_38_ ( .D(n14), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[38]) );
  fd2qd1_hd r_y_data_reg_37_ ( .D(n12), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[37]) );
  fd2qd1_hd r_y_data_reg_36_ ( .D(n10), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[36]) );
  fd2qd1_hd r_y_data_reg_35_ ( .D(n8), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[35]) );
  fd2qd1_hd r_y_data_reg_34_ ( .D(n6), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[34]) );
  fd2qd1_hd r_y_data_reg_33_ ( .D(n4), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[33]) );
  fd2qd1_hd r_y_data_reg_32_ ( .D(n2), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[32]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(n159), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(n158), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(n157), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(n156), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(n155), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(n154), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[5]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(n153), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(n152), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(n151), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(n150), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(n149), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(n148), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(n147), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(n146), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(n145), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(n144), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(n143), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(n142), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(n141), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(n140), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(n139), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(n138), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(n137), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(n136), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(n135), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(n134), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(n133), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(n132), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(n131), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(n130), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(n129), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(n128), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[31]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(n166), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(n63), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(n61), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(n59), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(n57), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(n55), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(n53), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(n51), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(n49), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(n47), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(n45), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(n43), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(n41), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(n39), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(n37), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(n35), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(n33), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(n31), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(n29), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(n27), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(n25), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(n23), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(n21), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(n19), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(n17), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(n15), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(n13), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(n11), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(n9), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[3])
         );
  fd2qd1_hd r_y_data_reg_2_ ( .D(n7), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[2])
         );
  fd2qd1_hd r_y_data_reg_1_ ( .D(n5), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[1])
         );
  fd2qd1_hd r_y_data_reg_0_ ( .D(n3), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[0])
         );
  fd2qd1_hd r_add_Z_ACK_reg ( .D(n528), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_Z_ACK) );
  fd2qd1_hd r_add_AB_STB_reg ( .D(n532), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_AB_STB) );
  fd2qd1_hd r_mult_Z_ACK_reg ( .D(n529), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_Z_ACK) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(n566), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[31]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(n534), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(n535), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(n536), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(n537), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(n538), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(n539), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(n540), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(n541), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(n542), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(n543), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(n544), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(n545), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(n546), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(n547), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(n548), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(n549), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(n550), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(n551), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(n552), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(n553), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(n554), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(n555), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[9]) );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(n556), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[8]) );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(n557), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[7]) );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(n558), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[6]) );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(n559), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[5]) );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(n560), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[4]) );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(n561), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[3]) );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(n562), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[2]) );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(n563), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[1]) );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(n564), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[0]) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n381), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_mult_AB_STB_reg ( .D(n435), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_AB_STB) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n738), .E(N814), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(N807), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_pstate_0_) );
  clknd2d1_hd U586 ( .A(n207), .B(n164), .Y(n825) );
  clknd2d1_hd U587 ( .A(n832), .B(n997), .Y(n834) );
  clknd2d1_hd U588 ( .A(n570), .B(w_add_Z_STB), .Y(n762) );
  nid1_hd U589 ( .A(n696), .Y(n759) );
  clknd2d1_hd U590 ( .A(n990), .B(n207), .Y(n835) );
  clknd2d1_hd U591 ( .A(n823), .B(n1001), .Y(n824) );
  nid1_hd U592 ( .A(n688), .Y(n627) );
  clknd2d1_hd U593 ( .A(n1001), .B(n764), .Y(n986) );
  nid1_hd U594 ( .A(n759), .Y(n731) );
  nid1_hd U595 ( .A(n696), .Y(n756) );
  nid1_hd U596 ( .A(n569), .Y(n696) );
  nid1_hd U597 ( .A(n731), .Y(n730) );
  nid1_hd U598 ( .A(n757), .Y(n754) );
  nid1_hd U599 ( .A(n759), .Y(n755) );
  clknd2d1_hd U600 ( .A(n823), .B(n822), .Y(n965) );
  nid1_hd U601 ( .A(n967), .Y(n693) );
  nid1_hd U602 ( .A(n686), .Y(n597) );
  clknd2d1_hd U603 ( .A(n822), .B(n764), .Y(n983) );
  clknd2d1_hd U604 ( .A(n161), .B(n760), .Y(n252) );
  nid1_hd U605 ( .A(n755), .Y(n729) );
  nid1_hd U606 ( .A(n870), .Y(n678) );
  nid1_hd U607 ( .A(n695), .Y(n673) );
  nid1_hd U608 ( .A(n694), .Y(n665) );
  nid1_hd U609 ( .A(n870), .Y(n677) );
  nid1_hd U610 ( .A(n695), .Y(n672) );
  nid1_hd U611 ( .A(n694), .Y(n666) );
  nid1_hd U612 ( .A(n870), .Y(n676) );
  nid1_hd U613 ( .A(n695), .Y(n671) );
  nid1_hd U614 ( .A(n694), .Y(n667) );
  nid1_hd U615 ( .A(n870), .Y(n675) );
  nid1_hd U616 ( .A(n695), .Y(n670) );
  nid1_hd U617 ( .A(n694), .Y(n668) );
  clknd2d1_hd U618 ( .A(n833), .B(n834), .Y(n873) );
  nid1_hd U619 ( .A(n873), .Y(n694) );
  nid1_hd U620 ( .A(n870), .Y(n674) );
  nid1_hd U621 ( .A(n695), .Y(n669) );
  nid1_hd U622 ( .A(n694), .Y(n664) );
  nid1_hd U623 ( .A(n871), .Y(n695) );
  clknd2d1_hd U624 ( .A(r_pstate_0_), .B(n161), .Y(n877) );
  nid1_hd U625 ( .A(n758), .Y(n753) );
  nid1_hd U626 ( .A(n753), .Y(n752) );
  nid1_hd U627 ( .A(n753), .Y(n751) );
  nid1_hd U628 ( .A(n753), .Y(n750) );
  nid1_hd U629 ( .A(n758), .Y(n749) );
  nid1_hd U630 ( .A(n729), .Y(n739) );
  nid1_hd U631 ( .A(n757), .Y(n740) );
  nid1_hd U632 ( .A(n757), .Y(n741) );
  nid1_hd U633 ( .A(n757), .Y(n742) );
  nid1_hd U634 ( .A(n569), .Y(n758) );
  nid1_hd U635 ( .A(n966), .Y(n690) );
  nid1_hd U636 ( .A(n971), .Y(n691) );
  nid1_hd U637 ( .A(n693), .Y(n653) );
  nid1_hd U638 ( .A(n965), .Y(n642) );
  nid1_hd U639 ( .A(n690), .Y(n636) );
  nid1_hd U640 ( .A(n691), .Y(n641) );
  nid1_hd U641 ( .A(n984), .Y(n687) );
  nid1_hd U642 ( .A(n967), .Y(n654) );
  nid1_hd U643 ( .A(n692), .Y(n643) );
  nid1_hd U644 ( .A(n690), .Y(n635) );
  nid1_hd U645 ( .A(n691), .Y(n640) );
  nid1_hd U646 ( .A(n693), .Y(n655) );
  nid1_hd U647 ( .A(n965), .Y(n644) );
  nid1_hd U648 ( .A(n690), .Y(n634) );
  nid1_hd U649 ( .A(n691), .Y(n639) );
  nid1_hd U650 ( .A(n598), .Y(n586) );
  nid1_hd U651 ( .A(n967), .Y(n656) );
  nid1_hd U652 ( .A(n965), .Y(n645) );
  nid1_hd U653 ( .A(n690), .Y(n633) );
  nid1_hd U654 ( .A(n691), .Y(n638) );
  nid1_hd U655 ( .A(n598), .Y(n587) );
  nid1_hd U656 ( .A(n611), .Y(n599) );
  nid1_hd U657 ( .A(n967), .Y(n657) );
  nid1_hd U658 ( .A(n965), .Y(n646) );
  nid1_hd U659 ( .A(n584), .Y(n578) );
  nid1_hd U660 ( .A(n584), .Y(n579) );
  nid1_hd U661 ( .A(n611), .Y(n600) );
  nid1_hd U662 ( .A(n688), .Y(n616) );
  nid1_hd U663 ( .A(n583), .Y(n580) );
  nid1_hd U664 ( .A(n984), .Y(n605) );
  nid1_hd U665 ( .A(n688), .Y(n617) );
  nid1_hd U666 ( .A(n578), .Y(n581) );
  nid1_hd U667 ( .A(n627), .Y(n612) );
  nid1_hd U668 ( .A(n598), .Y(n588) );
  nid1_hd U669 ( .A(n984), .Y(n603) );
  nid1_hd U670 ( .A(n597), .Y(n591) );
  nid1_hd U671 ( .A(n983), .Y(n618) );
  nid1_hd U672 ( .A(n583), .Y(n582) );
  nid1_hd U673 ( .A(n627), .Y(n613) );
  nid1_hd U674 ( .A(n611), .Y(n601) );
  nid1_hd U675 ( .A(n597), .Y(n589) );
  nid1_hd U676 ( .A(n627), .Y(n619) );
  nid1_hd U677 ( .A(n627), .Y(n614) );
  nid1_hd U678 ( .A(n597), .Y(n590) );
  nid1_hd U679 ( .A(n610), .Y(n604) );
  nid1_hd U680 ( .A(n627), .Y(n615) );
  nid1_hd U681 ( .A(n610), .Y(n602) );
  nid1_hd U682 ( .A(n688), .Y(n620) );
  nid1_hd U683 ( .A(n598), .Y(n592) );
  nid1_hd U684 ( .A(n627), .Y(n621) );
  nid1_hd U685 ( .A(n598), .Y(n593) );
  nid1_hd U686 ( .A(n687), .Y(n611) );
  nid1_hd U687 ( .A(n690), .Y(n632) );
  nid1_hd U688 ( .A(n691), .Y(n637) );
  nid1_hd U689 ( .A(n756), .Y(n732) );
  clknd2d1_hd U690 ( .A(o_X_DATA_READY), .B(i_X_DATA_VALID), .Y(n569) );
  nid1_hd U691 ( .A(n731), .Y(n757) );
  nid1_hd U692 ( .A(n756), .Y(n737) );
  nid1_hd U693 ( .A(n756), .Y(n736) );
  nid1_hd U694 ( .A(n756), .Y(n735) );
  nid1_hd U695 ( .A(n756), .Y(n734) );
  nid1_hd U696 ( .A(n756), .Y(n733) );
  nid1_hd U697 ( .A(n754), .Y(n743) );
  nid1_hd U698 ( .A(n754), .Y(n744) );
  nid1_hd U699 ( .A(n754), .Y(n745) );
  nid1_hd U700 ( .A(n754), .Y(n746) );
  nid1_hd U701 ( .A(n754), .Y(n747) );
  nid1_hd U702 ( .A(n754), .Y(n748) );
  nid1_hd U703 ( .A(n652), .Y(n647) );
  nid1_hd U704 ( .A(n967), .Y(n658) );
  nid1_hd U705 ( .A(n826), .Y(n684) );
  nid1_hd U706 ( .A(n652), .Y(n648) );
  nid1_hd U707 ( .A(n967), .Y(n659) );
  nid1_hd U708 ( .A(n826), .Y(n683) );
  nid1_hd U709 ( .A(n693), .Y(n660) );
  nid1_hd U710 ( .A(n692), .Y(n649) );
  nid1_hd U711 ( .A(n687), .Y(n610) );
  nid1_hd U712 ( .A(n826), .Y(n682) );
  nid1_hd U713 ( .A(n610), .Y(n609) );
  nid1_hd U714 ( .A(n693), .Y(n661) );
  nid1_hd U715 ( .A(n692), .Y(n650) );
  nid1_hd U716 ( .A(n597), .Y(n595) );
  nid1_hd U717 ( .A(n826), .Y(n681) );
  nid1_hd U718 ( .A(n693), .Y(n662) );
  nid1_hd U719 ( .A(n965), .Y(n651) );
  nid1_hd U720 ( .A(n692), .Y(n652) );
  nid1_hd U721 ( .A(n826), .Y(n680) );
  nid1_hd U722 ( .A(n610), .Y(n608) );
  nid1_hd U723 ( .A(n818), .Y(n689) );
  nid1_hd U724 ( .A(n689), .Y(n631) );
  nid1_hd U725 ( .A(n689), .Y(n630) );
  nid1_hd U726 ( .A(n689), .Y(n629) );
  nid1_hd U727 ( .A(n689), .Y(n628) );
  nid1_hd U728 ( .A(n983), .Y(n622) );
  nid1_hd U729 ( .A(n597), .Y(n594) );
  nid1_hd U730 ( .A(n597), .Y(n596) );
  nid1_hd U731 ( .A(n983), .Y(n623) );
  nid1_hd U732 ( .A(n984), .Y(n607) );
  nid1_hd U733 ( .A(n686), .Y(n598) );
  nid1_hd U734 ( .A(n626), .Y(n624) );
  nid1_hd U735 ( .A(n984), .Y(n606) );
  nid1_hd U736 ( .A(n984), .Y(n686) );
  nid1_hd U737 ( .A(n983), .Y(n688) );
  nid1_hd U738 ( .A(n626), .Y(n625) );
  nid1_hd U739 ( .A(n688), .Y(n626) );
  nr2d1_hd U740 ( .A(r_pstate_0_), .B(n161), .Y(n1001) );
  nid1_hd U741 ( .A(n729), .Y(n738) );
  clknd2d1_hd U742 ( .A(n816), .B(n819), .Y(n817) );
  clknd2d1_hd U743 ( .A(n991), .B(n875), .Y(n816) );
  clknd2d1_hd U744 ( .A(n709), .B(i_X_DATA[31]), .Y(n1034) );
  clknd2d1_hd U745 ( .A(n711), .B(i_X_DATA[30]), .Y(n1036) );
  clknd2d1_hd U746 ( .A(n712), .B(i_X_DATA[29]), .Y(n1038) );
  clknd2d1_hd U747 ( .A(n710), .B(i_X_DATA[28]), .Y(n1040) );
  clknd2d1_hd U748 ( .A(n712), .B(i_X_DATA[27]), .Y(n1042) );
  clknd2d1_hd U749 ( .A(n712), .B(i_X_DATA[26]), .Y(n1044) );
  clknd2d1_hd U750 ( .A(n712), .B(i_X_DATA[25]), .Y(n1046) );
  clknd2d1_hd U751 ( .A(n710), .B(i_X_DATA[24]), .Y(n1048) );
  clknd2d1_hd U752 ( .A(n708), .B(i_X_DATA[23]), .Y(n1050) );
  clknd2d1_hd U753 ( .A(n712), .B(i_X_DATA[22]), .Y(n1052) );
  clknd2d1_hd U754 ( .A(n712), .B(i_X_DATA[21]), .Y(n1054) );
  clknd2d1_hd U755 ( .A(n711), .B(i_X_DATA[20]), .Y(n1056) );
  clknd2d1_hd U756 ( .A(n711), .B(i_X_DATA[19]), .Y(n1058) );
  clknd2d1_hd U757 ( .A(n710), .B(i_X_DATA[18]), .Y(n1060) );
  clknd2d1_hd U758 ( .A(n711), .B(i_X_DATA[17]), .Y(n1062) );
  clknd2d1_hd U759 ( .A(n707), .B(i_X_DATA[16]), .Y(n1064) );
  clknd2d1_hd U760 ( .A(n711), .B(i_X_DATA[15]), .Y(n1066) );
  clknd2d1_hd U761 ( .A(n711), .B(i_X_DATA[14]), .Y(n1068) );
  clknd2d1_hd U762 ( .A(n708), .B(i_X_DATA[13]), .Y(n1070) );
  clknd2d1_hd U763 ( .A(n710), .B(i_X_DATA[12]), .Y(n1072) );
  clknd2d1_hd U764 ( .A(n708), .B(i_X_DATA[11]), .Y(n1074) );
  clknd2d1_hd U765 ( .A(n710), .B(i_X_DATA[10]), .Y(n1076) );
  clknd2d1_hd U766 ( .A(n710), .B(i_X_DATA[9]), .Y(n1078) );
  clknd2d1_hd U767 ( .A(n709), .B(i_X_DATA[8]), .Y(n1080) );
  clknd2d1_hd U768 ( .A(n709), .B(i_X_DATA[7]), .Y(n1082) );
  clknd2d1_hd U769 ( .A(n709), .B(i_X_DATA[6]), .Y(n1084) );
  clknd2d1_hd U770 ( .A(n709), .B(i_X_DATA[5]), .Y(n1086) );
  clknd2d1_hd U771 ( .A(n709), .B(i_X_DATA[4]), .Y(n1088) );
  clknd2d1_hd U772 ( .A(n707), .B(i_X_DATA[3]), .Y(n1090) );
  clknd2d1_hd U773 ( .A(n708), .B(i_X_DATA[2]), .Y(n1092) );
  clknd2d1_hd U774 ( .A(n708), .B(i_X_DATA[1]), .Y(n1094) );
  clknd2d1_hd U775 ( .A(n708), .B(i_X_DATA[0]), .Y(n1096) );
  nid1_hd U776 ( .A(n826), .Y(n685) );
  nid1_hd U777 ( .A(n693), .Y(n663) );
  nid1_hd U778 ( .A(n870), .Y(n679) );
  nid1_hd U779 ( .A(n965), .Y(n692) );
  nid1_hd U780 ( .A(n585), .Y(n583) );
  scg10d1_hd U781 ( .A(n744), .B(r_x_data[53]), .C(r_x_data[85]), .D(n727), 
        .Y(n74) );
  scg10d1_hd U782 ( .A(n745), .B(r_x_data[47]), .C(r_x_data[79]), .D(n726), 
        .Y(n80) );
  scg10d1_hd U783 ( .A(n745), .B(r_x_data[48]), .C(r_x_data[80]), .D(n726), 
        .Y(n79) );
  scg10d1_hd U784 ( .A(n744), .B(r_x_data[52]), .C(r_x_data[84]), .D(n727), 
        .Y(n75) );
  scg10d1_hd U785 ( .A(n745), .B(r_x_data[51]), .C(r_x_data[83]), .D(n727), 
        .Y(n76) );
  scg10d1_hd U786 ( .A(n745), .B(r_x_data[50]), .C(r_x_data[82]), .D(n727), 
        .Y(n77) );
  scg10d1_hd U787 ( .A(n745), .B(r_x_data[49]), .C(r_x_data[81]), .D(n727), 
        .Y(n78) );
  scg10d1_hd U788 ( .A(n745), .B(r_x_data[46]), .C(r_x_data[78]), .D(n726), 
        .Y(n81) );
  scg10d1_hd U789 ( .A(n743), .B(r_x_data[63]), .C(r_x_data[95]), .D(n723), 
        .Y(n64) );
  scg10d1_hd U790 ( .A(n748), .B(r_x_data[32]), .C(r_x_data[64]), .D(n724), 
        .Y(n95) );
  scg10d1_hd U791 ( .A(n746), .B(r_x_data[45]), .C(r_x_data[77]), .D(n726), 
        .Y(n82) );
  scg10d1_hd U792 ( .A(n748), .B(r_x_data[33]), .C(r_x_data[65]), .D(n724), 
        .Y(n94) );
  scg10d1_hd U793 ( .A(n744), .B(r_x_data[54]), .C(r_x_data[86]), .D(n727), 
        .Y(n73) );
  scg10d1_hd U794 ( .A(n747), .B(r_x_data[34]), .C(r_x_data[66]), .D(n724), 
        .Y(n93) );
  scg10d1_hd U795 ( .A(n746), .B(r_x_data[44]), .C(r_x_data[76]), .D(n726), 
        .Y(n83) );
  scg10d1_hd U796 ( .A(n747), .B(r_x_data[35]), .C(r_x_data[67]), .D(n724), 
        .Y(n92) );
  scg10d1_hd U797 ( .A(n743), .B(r_x_data[62]), .C(r_x_data[94]), .D(n724), 
        .Y(n65) );
  scg10d1_hd U798 ( .A(n744), .B(r_x_data[55]), .C(r_x_data[87]), .D(n728), 
        .Y(n72) );
  scg10d1_hd U799 ( .A(n747), .B(r_x_data[36]), .C(r_x_data[68]), .D(n724), 
        .Y(n91) );
  scg10d1_hd U800 ( .A(n746), .B(r_x_data[43]), .C(r_x_data[75]), .D(n726), 
        .Y(n84) );
  scg10d1_hd U801 ( .A(n743), .B(r_x_data[61]), .C(r_x_data[93]), .D(n713), 
        .Y(n66) );
  scg10d1_hd U802 ( .A(n747), .B(r_x_data[37]), .C(r_x_data[69]), .D(n725), 
        .Y(n90) );
  scg10d1_hd U803 ( .A(n747), .B(r_x_data[38]), .C(r_x_data[70]), .D(n725), 
        .Y(n89) );
  scg10d1_hd U804 ( .A(n744), .B(r_x_data[56]), .C(r_x_data[88]), .D(n728), 
        .Y(n71) );
  scg10d1_hd U805 ( .A(n743), .B(r_x_data[60]), .C(r_x_data[92]), .D(n728), 
        .Y(n67) );
  scg10d1_hd U806 ( .A(n747), .B(r_x_data[39]), .C(r_x_data[71]), .D(n725), 
        .Y(n88) );
  scg10d1_hd U807 ( .A(n743), .B(r_x_data[59]), .C(r_x_data[91]), .D(n728), 
        .Y(n68) );
  scg10d1_hd U808 ( .A(n744), .B(r_x_data[57]), .C(r_x_data[89]), .D(n728), 
        .Y(n70) );
  scg10d1_hd U809 ( .A(n746), .B(r_x_data[40]), .C(r_x_data[72]), .D(n725), 
        .Y(n87) );
  scg10d1_hd U810 ( .A(n748), .B(r_y_data[15]), .C(r_y_data[47]), .D(n718), 
        .Y(n32) );
  scg10d1_hd U811 ( .A(n743), .B(r_x_data[58]), .C(r_x_data[90]), .D(n728), 
        .Y(n69) );
  scg10d1_hd U812 ( .A(n746), .B(r_x_data[42]), .C(r_x_data[74]), .D(n725), 
        .Y(n85) );
  scg10d1_hd U813 ( .A(n748), .B(r_y_data[16]), .C(r_y_data[48]), .D(n718), 
        .Y(n34) );
  scg10d1_hd U814 ( .A(n746), .B(r_x_data[41]), .C(r_x_data[73]), .D(n725), 
        .Y(n86) );
  scg10d1_hd U815 ( .A(n748), .B(o_Y_DATA[15]), .C(r_y_data[15]), .D(n718), 
        .Y(n33) );
  scg10d1_hd U816 ( .A(n748), .B(o_Y_DATA[14]), .C(r_y_data[14]), .D(n717), 
        .Y(n31) );
  scg10d1_hd U817 ( .A(n741), .B(o_Y_DATA[26]), .C(r_y_data[26]), .D(n722), 
        .Y(n55) );
  scg10d1_hd U818 ( .A(n741), .B(o_Y_DATA[25]), .C(r_y_data[25]), .D(n721), 
        .Y(n53) );
  scg10d1_hd U819 ( .A(n741), .B(o_Y_DATA[27]), .C(r_y_data[27]), .D(n722), 
        .Y(n57) );
  scg10d1_hd U820 ( .A(n740), .B(o_Y_DATA[24]), .C(r_y_data[24]), .D(n721), 
        .Y(n51) );
  scg10d1_hd U821 ( .A(n758), .B(r_y_data[31]), .C(r_y_data[63]), .D(n713), 
        .Y(n165) );
  scg10d1_hd U822 ( .A(n740), .B(o_Y_DATA[23]), .C(r_y_data[23]), .D(n721), 
        .Y(n49) );
  scg10d1_hd U823 ( .A(n740), .B(o_Y_DATA[22]), .C(r_y_data[22]), .D(n720), 
        .Y(n47) );
  scg10d1_hd U824 ( .A(n749), .B(o_Y_DATA[12]), .C(r_y_data[12]), .D(n717), 
        .Y(n27) );
  scg10d1_hd U825 ( .A(n739), .B(o_Y_DATA[21]), .C(r_y_data[21]), .D(n720), 
        .Y(n45) );
  scg10d1_hd U826 ( .A(n758), .B(o_Y_DATA[0]), .C(r_y_data[0]), .D(n713), .Y(
        n3) );
  scg10d1_hd U827 ( .A(n739), .B(o_Y_DATA[20]), .C(r_y_data[20]), .D(n720), 
        .Y(n43) );
  scg10d1_hd U828 ( .A(n753), .B(o_Y_DATA[1]), .C(r_y_data[1]), .D(n718), .Y(
        n5) );
  scg10d1_hd U829 ( .A(n739), .B(o_Y_DATA[19]), .C(r_y_data[19]), .D(n719), 
        .Y(n41) );
  scg10d1_hd U830 ( .A(n752), .B(o_Y_DATA[2]), .C(r_y_data[2]), .D(n713), .Y(
        n7) );
  scg10d1_hd U831 ( .A(n738), .B(o_Y_DATA[18]), .C(r_y_data[18]), .D(n719), 
        .Y(n39) );
  scg10d1_hd U832 ( .A(n738), .B(o_Y_DATA[17]), .C(r_y_data[17]), .D(n719), 
        .Y(n37) );
  scg10d1_hd U833 ( .A(n738), .B(o_Y_DATA[16]), .C(r_y_data[16]), .D(n718), 
        .Y(n35) );
  scg10d1_hd U834 ( .A(n749), .B(o_Y_DATA[13]), .C(r_y_data[13]), .D(n717), 
        .Y(n29) );
  scg10d1_hd U835 ( .A(n738), .B(r_y_data[17]), .C(r_y_data[49]), .D(n719), 
        .Y(n36) );
  scg10d1_hd U836 ( .A(n738), .B(r_y_data[18]), .C(r_y_data[50]), .D(n719), 
        .Y(n38) );
  scg10d1_hd U837 ( .A(n749), .B(r_y_data[14]), .C(r_y_data[46]), .D(n717), 
        .Y(n30) );
  scg10d1_hd U838 ( .A(n749), .B(r_y_data[13]), .C(r_y_data[45]), .D(n717), 
        .Y(n28) );
  scg10d1_hd U839 ( .A(n739), .B(r_y_data[19]), .C(r_y_data[51]), .D(n719), 
        .Y(n40) );
  scg10d1_hd U840 ( .A(n750), .B(r_y_data[11]), .C(r_y_data[43]), .D(n717), 
        .Y(n24) );
  scg10d1_hd U841 ( .A(n739), .B(r_y_data[20]), .C(r_y_data[52]), .D(n720), 
        .Y(n42) );
  scg10d1_hd U842 ( .A(n739), .B(r_y_data[21]), .C(r_y_data[53]), .D(n720), 
        .Y(n44) );
  scg10d1_hd U843 ( .A(n740), .B(r_y_data[22]), .C(r_y_data[54]), .D(n720), 
        .Y(n46) );
  scg10d1_hd U844 ( .A(n740), .B(r_y_data[23]), .C(r_y_data[55]), .D(n721), 
        .Y(n48) );
  scg10d1_hd U845 ( .A(n752), .B(r_y_data[4]), .C(r_y_data[36]), .D(n713), .Y(
        n10) );
  scg10d1_hd U846 ( .A(n753), .B(r_y_data[2]), .C(r_y_data[34]), .D(n713), .Y(
        n6) );
  scg10d1_hd U847 ( .A(n740), .B(r_y_data[24]), .C(r_y_data[56]), .D(n721), 
        .Y(n50) );
  scg10d1_hd U848 ( .A(n753), .B(r_y_data[0]), .C(r_y_data[32]), .D(n718), .Y(
        n2) );
  scg10d1_hd U849 ( .A(n742), .B(o_Y_DATA[28]), .C(r_y_data[28]), .D(n722), 
        .Y(n59) );
  scg10d1_hd U850 ( .A(n742), .B(r_y_data[30]), .C(r_y_data[62]), .D(n723), 
        .Y(n62) );
  scg10d1_hd U851 ( .A(n742), .B(r_y_data[28]), .C(r_y_data[60]), .D(n722), 
        .Y(n58) );
  scg10d1_hd U852 ( .A(n742), .B(o_Y_DATA[29]), .C(r_y_data[29]), .D(n723), 
        .Y(n61) );
  scg10d1_hd U853 ( .A(n741), .B(r_y_data[25]), .C(r_y_data[57]), .D(n721), 
        .Y(n52) );
  scg10d1_hd U854 ( .A(n741), .B(r_y_data[26]), .C(r_y_data[58]), .D(n722), 
        .Y(n54) );
  scg10d1_hd U855 ( .A(n741), .B(r_y_data[27]), .C(r_y_data[59]), .D(n722), 
        .Y(n56) );
  scg10d1_hd U856 ( .A(n742), .B(r_y_data[29]), .C(r_y_data[61]), .D(n723), 
        .Y(n60) );
  scg10d1_hd U857 ( .A(n742), .B(o_Y_DATA[30]), .C(r_y_data[30]), .D(n723), 
        .Y(n63) );
  scg10d1_hd U858 ( .A(n758), .B(o_Y_DATA[31]), .C(r_y_data[31]), .D(n723), 
        .Y(n166) );
  scg10d1_hd U859 ( .A(n750), .B(o_Y_DATA[10]), .C(r_y_data[10]), .D(n716), 
        .Y(n23) );
  scg10d1_hd U860 ( .A(n750), .B(o_Y_DATA[9]), .C(r_y_data[9]), .D(n716), .Y(
        n21) );
  scg10d1_hd U861 ( .A(n750), .B(o_Y_DATA[8]), .C(r_y_data[8]), .D(n716), .Y(
        n19) );
  scg10d1_hd U862 ( .A(n751), .B(o_Y_DATA[7]), .C(r_y_data[7]), .D(n714), .Y(
        n17) );
  scg10d1_hd U863 ( .A(n752), .B(o_Y_DATA[3]), .C(r_y_data[3]), .D(n715), .Y(
        n9) );
  scg10d1_hd U864 ( .A(n751), .B(o_Y_DATA[6]), .C(r_y_data[6]), .D(n714), .Y(
        n15) );
  scg10d1_hd U865 ( .A(n751), .B(o_Y_DATA[5]), .C(r_y_data[5]), .D(n714), .Y(
        n13) );
  scg10d1_hd U866 ( .A(n752), .B(o_Y_DATA[4]), .C(r_y_data[4]), .D(n714), .Y(
        n11) );
  scg10d1_hd U867 ( .A(n752), .B(r_y_data[3]), .C(r_y_data[35]), .D(n715), .Y(
        n8) );
  scg10d1_hd U868 ( .A(n752), .B(r_y_data[5]), .C(r_y_data[37]), .D(n714), .Y(
        n12) );
  scg10d1_hd U869 ( .A(n751), .B(r_y_data[6]), .C(r_y_data[38]), .D(n716), .Y(
        n14) );
  scg10d1_hd U870 ( .A(n751), .B(r_y_data[7]), .C(r_y_data[39]), .D(n714), .Y(
        n16) );
  scg10d1_hd U871 ( .A(n751), .B(r_y_data[8]), .C(r_y_data[40]), .D(n715), .Y(
        n18) );
  scg10d1_hd U872 ( .A(n750), .B(r_y_data[9]), .C(r_y_data[41]), .D(n715), .Y(
        n20) );
  scg10d1_hd U873 ( .A(n750), .B(r_y_data[10]), .C(r_y_data[42]), .D(n715), 
        .Y(n22) );
  scg10d1_hd U874 ( .A(n749), .B(r_y_data[12]), .C(r_y_data[44]), .D(n716), 
        .Y(n26) );
  scg10d1_hd U875 ( .A(n749), .B(o_Y_DATA[11]), .C(r_y_data[11]), .D(n716), 
        .Y(n25) );
  scg10d1_hd U876 ( .A(n758), .B(r_y_data[1]), .C(r_y_data[33]), .D(n715), .Y(
        n4) );
  ivd1_hd U877 ( .A(n991), .Y(n570) );
  scg12d1_hd U878 ( .A(n664), .B(n1001), .C(n835), .Y(n870) );
  nd2bd1_hd U879 ( .AN(n632), .B(n637), .Y(n826) );
  scg6d1_hd U880 ( .A(n832), .B(n821), .C(n876), .Y(n823) );
  nr2d1_hd U881 ( .A(n825), .B(n875), .Y(n984) );
  ivd1_hd U882 ( .A(n998), .Y(n875) );
  ivd1_hd U883 ( .A(n986), .Y(n584) );
  ivd1_hd U884 ( .A(n762), .Y(n832) );
  nr2d1_hd U885 ( .A(n825), .B(n824), .Y(n967) );
  ivd1_hd U886 ( .A(n731), .Y(n704) );
  ivd1_hd U887 ( .A(n733), .Y(n698) );
  ivd1_hd U888 ( .A(n755), .Y(n705) );
  ivd1_hd U889 ( .A(n755), .Y(n706) );
  ivd1_hd U890 ( .A(n986), .Y(n585) );
  ivd1_hd U891 ( .A(n579), .Y(n571) );
  ivd1_hd U892 ( .A(n834), .Y(n871) );
  scg6d1_hd U893 ( .A(n875), .B(n831), .C(n835), .Y(n833) );
  ivd1_hd U894 ( .A(n733), .Y(n697) );
  ivd1_hd U895 ( .A(n729), .Y(n707) );
  ivd1_hd U896 ( .A(n732), .Y(n700) );
  ivd1_hd U897 ( .A(n730), .Y(n712) );
  ivd1_hd U898 ( .A(n732), .Y(n701) );
  ivd1_hd U899 ( .A(n730), .Y(n711) );
  ivd1_hd U900 ( .A(n732), .Y(n699) );
  ivd1_hd U901 ( .A(n729), .Y(n728) );
  ivd1_hd U902 ( .A(n729), .Y(n727) );
  ivd1_hd U903 ( .A(n729), .Y(n726) );
  ivd1_hd U904 ( .A(n730), .Y(n719) );
  ivd1_hd U905 ( .A(n730), .Y(n717) );
  ivd1_hd U906 ( .A(n730), .Y(n718) );
  ivd1_hd U907 ( .A(n730), .Y(n713) );
  nr2d1_hd U908 ( .A(n586), .B(n579), .Y(n818) );
  ivd1_hd U909 ( .A(n584), .Y(n577) );
  ivd1_hd U910 ( .A(n583), .Y(n576) );
  ivd1_hd U911 ( .A(n578), .Y(n575) );
  ivd1_hd U912 ( .A(n578), .Y(n574) );
  ivd1_hd U913 ( .A(n578), .Y(n573) );
  ivd1_hd U914 ( .A(n578), .Y(n572) );
  ivd1_hd U915 ( .A(n877), .Y(n819) );
  nr2d1_hd U916 ( .A(n877), .B(n763), .Y(n998) );
  oa21d1_hd U917 ( .A(n825), .B(n831), .C(n877), .Y(n764) );
  ivd1_hd U918 ( .A(n696), .Y(n715) );
  ivd1_hd U919 ( .A(n696), .Y(n716) );
  ivd1_hd U920 ( .A(n696), .Y(n703) );
  nr2bd1_hd U921 ( .AN(n252), .B(n987), .Y(n995) );
  ivd1_hd U922 ( .A(n759), .Y(n714) );
  ivd1_hd U923 ( .A(n731), .Y(n709) );
  ivd1_hd U924 ( .A(n731), .Y(n708) );
  ivd1_hd U925 ( .A(n731), .Y(n710) );
  ivd1_hd U926 ( .A(n759), .Y(n721) );
  ivd1_hd U927 ( .A(n759), .Y(n722) );
  ivd1_hd U928 ( .A(n696), .Y(n702) );
  ivd1_hd U929 ( .A(n759), .Y(n720) );
  ivd1_hd U930 ( .A(n755), .Y(n723) );
  ivd1_hd U931 ( .A(n755), .Y(n725) );
  ivd1_hd U932 ( .A(n755), .Y(n724) );
  nr2d1_hd U933 ( .A(n824), .B(n835), .Y(n966) );
  nd2bd1_hd U934 ( .AN(n824), .B(n821), .Y(n971) );
  oa21d1_hd U935 ( .A(n825), .B(n763), .C(n819), .Y(n822) );
  nd3d1_hd U936 ( .A(n832), .B(w_mult_2_Z_STB), .C(w_mult_1_Z_STB), .Y(n831)
         );
  scg6d1_hd U937 ( .A(r_mult_1_A[15]), .B(n623), .C(n686), .Y(n420) );
  scg6d1_hd U938 ( .A(r_mult_2_A[13]), .B(n623), .C(n606), .Y(n396) );
  scg6d1_hd U939 ( .A(r_mult_1_A[12]), .B(n623), .C(n686), .Y(n422) );
  scg6d1_hd U940 ( .A(r_mult_1_A[24]), .B(n623), .C(n607), .Y(n413) );
  scg6d1_hd U941 ( .A(r_mult_1_A[25]), .B(n623), .C(n594), .Y(n412) );
  scg6d1_hd U942 ( .A(r_mult_1_A[14]), .B(n623), .C(n606), .Y(n421) );
  scg6d1_hd U943 ( .A(r_mult_1_A[4]), .B(n622), .C(n606), .Y(n430) );
  scg6d1_hd U944 ( .A(r_mult_1_A[8]), .B(n622), .C(n594), .Y(n426) );
  ivd1_hd U945 ( .A(r_x_data[1]), .Y(n1095) );
  ivd1_hd U946 ( .A(r_x_data[0]), .Y(n1097) );
  ivd1_hd U947 ( .A(r_x_data[12]), .Y(n1073) );
  ivd1_hd U948 ( .A(r_x_data[2]), .Y(n1093) );
  ivd1_hd U949 ( .A(r_x_data[11]), .Y(n1075) );
  ivd1_hd U950 ( .A(r_x_data[4]), .Y(n1089) );
  ivd1_hd U951 ( .A(r_x_data[5]), .Y(n1087) );
  ivd1_hd U952 ( .A(r_x_data[6]), .Y(n1085) );
  ivd1_hd U953 ( .A(r_x_data[8]), .Y(n1081) );
  ivd1_hd U954 ( .A(r_x_data[7]), .Y(n1083) );
  ivd1_hd U955 ( .A(r_x_data[13]), .Y(n1071) );
  ivd1_hd U956 ( .A(r_x_data[10]), .Y(n1077) );
  ivd1_hd U957 ( .A(r_x_data[9]), .Y(n1079) );
  ivd1_hd U958 ( .A(r_x_data[23]), .Y(n1051) );
  ivd1_hd U959 ( .A(r_x_data[24]), .Y(n1049) );
  ivd1_hd U960 ( .A(r_x_data[18]), .Y(n1061) );
  scg14d1_hd U961 ( .A(w_add_Z[30]), .B(n583), .C(n814), .Y(n436) );
  scg14d1_hd U962 ( .A(w_add_Z[17]), .B(n582), .C(n801), .Y(n449) );
  scg14d1_hd U963 ( .A(w_add_Z[20]), .B(n582), .C(n804), .Y(n446) );
  scg14d1_hd U964 ( .A(w_add_Z[18]), .B(n582), .C(n802), .Y(n448) );
  scg14d1_hd U965 ( .A(w_add_Z[21]), .B(n582), .C(n805), .Y(n445) );
  scg14d1_hd U966 ( .A(w_add_Z[19]), .B(n582), .C(n803), .Y(n447) );
  scg14d1_hd U967 ( .A(w_add_Z[22]), .B(n582), .C(n806), .Y(n444) );
  scg6d1_hd U968 ( .A(r_mult_2_A[25]), .B(n625), .C(n606), .Y(n387) );
  scg6d1_hd U969 ( .A(r_mult_2_A[31]), .B(n625), .C(n686), .Y(n382) );
  scg6d1_hd U970 ( .A(r_mult_2_A[4]), .B(n624), .C(n606), .Y(n403) );
  scg6d1_hd U971 ( .A(r_mult_2_A[14]), .B(n624), .C(n686), .Y(n395) );
  scg6d1_hd U972 ( .A(r_mult_2_A[21]), .B(n624), .C(n607), .Y(n390) );
  scg6d1_hd U973 ( .A(r_mult_2_A[8]), .B(n624), .C(n596), .Y(n399) );
  scg6d1_hd U974 ( .A(r_mult_1_A[9]), .B(n624), .C(n607), .Y(n425) );
  scg6d1_hd U975 ( .A(r_mult_2_A[24]), .B(n624), .C(n598), .Y(n388) );
  scg14d1_hd U976 ( .A(w_add_Z[1]), .B(n579), .C(n785), .Y(n465) );
  scg14d1_hd U977 ( .A(w_add_Z[23]), .B(n583), .C(n807), .Y(n443) );
  scg14d1_hd U978 ( .A(w_add_Z[24]), .B(n583), .C(n808), .Y(n442) );
  scg14d1_hd U979 ( .A(w_add_Z[2]), .B(n579), .C(n786), .Y(n464) );
  scg14d1_hd U980 ( .A(w_add_Z[3]), .B(n579), .C(n787), .Y(n463) );
  scg14d1_hd U981 ( .A(w_add_Z[4]), .B(n579), .C(n788), .Y(n462) );
  ivd1_hd U982 ( .A(r_x_data[44]), .Y(n1021) );
  ivd1_hd U983 ( .A(r_x_data[49]), .Y(n1016) );
  ivd1_hd U984 ( .A(r_x_data[43]), .Y(n1022) );
  ivd1_hd U985 ( .A(r_x_data[45]), .Y(n1020) );
  ivd1_hd U986 ( .A(r_x_data[47]), .Y(n1018) );
  ivd1_hd U987 ( .A(r_x_data[48]), .Y(n1017) );
  ivd1_hd U988 ( .A(r_x_data[31]), .Y(n1035) );
  ivd1_hd U989 ( .A(r_x_data[28]), .Y(n1041) );
  ivd1_hd U990 ( .A(o_Y_DATA[10]), .Y(n907) );
  ivd1_hd U991 ( .A(o_Y_DATA[6]), .Y(n895) );
  ivd1_hd U992 ( .A(o_Y_DATA[9]), .Y(n904) );
  ivd1_hd U993 ( .A(o_Y_DATA[5]), .Y(n892) );
  ivd1_hd U994 ( .A(o_Y_DATA[7]), .Y(n898) );
  ivd1_hd U995 ( .A(o_Y_DATA[24]), .Y(n949) );
  ivd1_hd U996 ( .A(o_Y_DATA[21]), .Y(n940) );
  ivd1_hd U997 ( .A(o_Y_DATA[23]), .Y(n946) );
  ivd1_hd U998 ( .A(o_Y_DATA[22]), .Y(n943) );
  ivd1_hd U999 ( .A(o_Y_DATA[12]), .Y(n913) );
  ivd1_hd U1000 ( .A(o_Y_DATA[19]), .Y(n934) );
  ivd1_hd U1001 ( .A(o_Y_DATA[8]), .Y(n901) );
  ivd1_hd U1002 ( .A(o_Y_DATA[20]), .Y(n937) );
  ivd1_hd U1003 ( .A(o_Y_DATA[11]), .Y(n910) );
  ivd1_hd U1004 ( .A(o_Y_DATA[4]), .Y(n889) );
  ivd1_hd U1005 ( .A(o_Y_DATA[2]), .Y(n883) );
  ivd1_hd U1006 ( .A(o_Y_DATA[31]), .Y(n837) );
  ivd1_hd U1007 ( .A(o_Y_DATA[3]), .Y(n886) );
  ivd1_hd U1008 ( .A(o_Y_DATA[1]), .Y(n880) );
  ivd1_hd U1009 ( .A(o_Y_DATA[0]), .Y(n840) );
  ivd1_hd U1010 ( .A(r_x_data[3]), .Y(n1091) );
  ivd1_hd U1011 ( .A(r_x_data[16]), .Y(n1065) );
  ivd1_hd U1012 ( .A(r_x_data[21]), .Y(n1055) );
  ivd1_hd U1013 ( .A(r_x_data[25]), .Y(n1047) );
  ivd1_hd U1014 ( .A(r_x_data[27]), .Y(n1043) );
  ivd1_hd U1015 ( .A(r_x_data[20]), .Y(n1057) );
  ivd1_hd U1016 ( .A(r_x_data[29]), .Y(n1039) );
  ivd1_hd U1017 ( .A(r_x_data[19]), .Y(n1059) );
  ivd1_hd U1018 ( .A(r_x_data[14]), .Y(n1069) );
  ivd1_hd U1019 ( .A(r_x_data[15]), .Y(n1067) );
  ivd1_hd U1020 ( .A(r_x_data[22]), .Y(n1053) );
  ivd1_hd U1021 ( .A(r_x_data[30]), .Y(n1037) );
  ivd1_hd U1022 ( .A(r_x_data[26]), .Y(n1045) );
  ivd1_hd U1023 ( .A(r_x_data[17]), .Y(n1063) );
  scg14d1_hd U1024 ( .A(r_mult_2_A[22]), .B(n626), .C(n577), .Y(n389) );
  scg14d1_hd U1025 ( .A(r_mult_2_A[19]), .B(n626), .C(n577), .Y(n392) );
  scg14d1_hd U1026 ( .A(r_mult_1_A[1]), .B(n625), .C(n577), .Y(n433) );
  scg14d1_hd U1027 ( .A(r_mult_1_A[2]), .B(n625), .C(n577), .Y(n432) );
  scg14d1_hd U1028 ( .A(r_mult_1_A[19]), .B(n626), .C(n577), .Y(n417) );
  scg14d1_hd U1029 ( .A(r_mult_1_A[0]), .B(n625), .C(n576), .Y(n434) );
  scg14d1_hd U1030 ( .A(r_mult_2_A[1]), .B(n626), .C(n576), .Y(n406) );
  scg14d1_hd U1031 ( .A(r_mult_1_A[16]), .B(n688), .C(n576), .Y(n419) );
  scg14d1_hd U1032 ( .A(r_mult_2_A[2]), .B(n625), .C(n576), .Y(n405) );
  scg14d1_hd U1033 ( .A(w_add_Z[31]), .B(n584), .C(n874), .Y(n533) );
  scg14d1_hd U1034 ( .A(w_add_Z[0]), .B(n578), .C(n784), .Y(n466) );
  scg4d1_hd U1035 ( .A(n685), .B(w_add_Z[30]), .C(n647), .D(r_add_B[30]), .E(
        n596), .F(r_x_data[94]), .G(n658), .H(w_mult_2_Z[30]), .Y(n350) );
  scg4d1_hd U1036 ( .A(n685), .B(w_add_Z[31]), .C(n647), .D(r_add_B[31]), .E(
        n610), .F(r_x_data[95]), .G(n658), .H(w_mult_2_Z[31]), .Y(n349) );
  scg4d1_hd U1037 ( .A(n684), .B(w_add_Z[24]), .C(n648), .D(r_add_B[24]), .E(
        n595), .F(r_x_data[88]), .G(n659), .H(w_mult_2_Z[24]), .Y(n356) );
  scg4d1_hd U1038 ( .A(n684), .B(w_add_Z[29]), .C(n647), .D(r_add_B[29]), .E(
        n609), .F(r_x_data[93]), .G(n658), .H(w_mult_2_Z[29]), .Y(n351) );
  scg4d1_hd U1039 ( .A(n684), .B(w_add_Z[26]), .C(n648), .D(r_add_B[26]), .E(
        n596), .F(r_x_data[90]), .G(n659), .H(w_mult_2_Z[26]), .Y(n354) );
  scg4d1_hd U1040 ( .A(n683), .B(w_add_Z[23]), .C(n648), .D(r_add_B[23]), .E(
        n609), .F(r_x_data[87]), .G(n659), .H(w_mult_2_Z[23]), .Y(n357) );
  scg4d1_hd U1041 ( .A(n684), .B(w_add_Z[28]), .C(n647), .D(r_add_B[28]), .E(
        n595), .F(r_x_data[92]), .G(n658), .H(w_mult_2_Z[28]), .Y(n352) );
  scg4d1_hd U1042 ( .A(n684), .B(w_add_Z[25]), .C(n648), .D(r_add_B[25]), .E(
        n609), .F(r_x_data[89]), .G(n659), .H(w_mult_2_Z[25]), .Y(n355) );
  scg4d1_hd U1043 ( .A(n683), .B(w_add_Z[22]), .C(n648), .D(r_add_B[22]), .E(
        n596), .F(r_x_data[86]), .G(n659), .H(w_mult_2_Z[22]), .Y(n358) );
  scg4d1_hd U1044 ( .A(n684), .B(w_add_Z[27]), .C(n648), .D(r_add_B[27]), .E(
        n609), .F(r_x_data[91]), .G(n659), .H(w_mult_2_Z[27]), .Y(n353) );
  scg4d1_hd U1045 ( .A(n680), .B(w_add_Z[0]), .C(n652), .D(r_add_B[0]), .E(
        n608), .F(r_x_data[64]), .G(n663), .H(w_mult_2_Z[0]), .Y(n380) );
  scg4d1_hd U1046 ( .A(n680), .B(w_add_Z[3]), .C(n652), .D(r_add_B[3]), .E(
        n594), .F(r_x_data[67]), .G(n663), .H(w_mult_2_Z[3]), .Y(n377) );
  scg4d1_hd U1047 ( .A(n680), .B(w_add_Z[2]), .C(n652), .D(r_add_B[2]), .E(
        n607), .F(r_x_data[66]), .G(n663), .H(w_mult_2_Z[2]), .Y(n378) );
  scg4d1_hd U1048 ( .A(n680), .B(w_add_Z[1]), .C(n652), .D(r_add_B[1]), .E(
        n594), .F(r_x_data[65]), .G(n663), .H(w_mult_2_Z[1]), .Y(n379) );
  ivd1_hd U1049 ( .A(r_x_data[41]), .Y(n1024) );
  ivd1_hd U1050 ( .A(r_x_data[40]), .Y(n1025) );
  ivd1_hd U1051 ( .A(r_x_data[38]), .Y(n1027) );
  ivd1_hd U1052 ( .A(r_x_data[59]), .Y(n1006) );
  ivd1_hd U1053 ( .A(r_x_data[35]), .Y(n1030) );
  ivd1_hd U1054 ( .A(r_x_data[56]), .Y(n1009) );
  ivd1_hd U1055 ( .A(r_x_data[52]), .Y(n1013) );
  ivd1_hd U1056 ( .A(r_x_data[62]), .Y(n1003) );
  ivd1_hd U1057 ( .A(r_x_data[36]), .Y(n1029) );
  ivd1_hd U1058 ( .A(r_x_data[42]), .Y(n1023) );
  ivd1_hd U1059 ( .A(r_x_data[46]), .Y(n1019) );
  ivd1_hd U1060 ( .A(r_x_data[50]), .Y(n1015) );
  ivd1_hd U1061 ( .A(r_x_data[57]), .Y(n1008) );
  ivd1_hd U1062 ( .A(r_x_data[60]), .Y(n1005) );
  ivd1_hd U1063 ( .A(r_x_data[32]), .Y(n1033) );
  ivd1_hd U1064 ( .A(r_x_data[63]), .Y(n1002) );
  ivd1_hd U1065 ( .A(r_x_data[58]), .Y(n1007) );
  ivd1_hd U1066 ( .A(r_x_data[39]), .Y(n1026) );
  ivd1_hd U1067 ( .A(r_x_data[54]), .Y(n1011) );
  ivd1_hd U1068 ( .A(r_x_data[37]), .Y(n1028) );
  ivd1_hd U1069 ( .A(r_x_data[55]), .Y(n1010) );
  ivd1_hd U1070 ( .A(r_x_data[33]), .Y(n1032) );
  ivd1_hd U1071 ( .A(r_x_data[53]), .Y(n1012) );
  ivd1_hd U1072 ( .A(r_x_data[34]), .Y(n1031) );
  ivd1_hd U1073 ( .A(r_x_data[61]), .Y(n1004) );
  ivd1_hd U1074 ( .A(r_x_data[51]), .Y(n1014) );
  scg4d1_hd U1075 ( .A(n682), .B(w_add_Z[17]), .C(n649), .D(r_add_B[17]), .E(
        n608), .F(r_x_data[81]), .G(n660), .H(w_mult_2_Z[17]), .Y(n363) );
  scg4d1_hd U1076 ( .A(n683), .B(w_add_Z[21]), .C(n649), .D(r_add_B[21]), .E(
        n608), .F(r_x_data[85]), .G(n660), .H(w_mult_2_Z[21]), .Y(n359) );
  scg4d1_hd U1077 ( .A(n683), .B(w_add_Z[19]), .C(n649), .D(r_add_B[19]), .E(
        n609), .F(r_x_data[83]), .G(n660), .H(w_mult_2_Z[19]), .Y(n361) );
  scg4d1_hd U1078 ( .A(n683), .B(w_add_Z[20]), .C(n649), .D(r_add_B[20]), .E(
        n595), .F(r_x_data[84]), .G(n660), .H(w_mult_2_Z[20]), .Y(n360) );
  scg4d1_hd U1079 ( .A(n683), .B(w_add_Z[18]), .C(n649), .D(r_add_B[18]), .E(
        n595), .F(r_x_data[82]), .G(n660), .H(w_mult_2_Z[18]), .Y(n362) );
  scg4d1_hd U1080 ( .A(n682), .B(w_add_Z[16]), .C(n649), .D(r_add_B[16]), .E(
        n596), .F(r_x_data[80]), .G(n660), .H(w_mult_2_Z[16]), .Y(n364) );
  scg4d1_hd U1081 ( .A(n681), .B(w_add_Z[10]), .C(n650), .D(r_add_B[10]), .E(
        n607), .F(r_x_data[74]), .G(n661), .H(w_mult_2_Z[10]), .Y(n370) );
  scg4d1_hd U1082 ( .A(n680), .B(w_add_Z[5]), .C(n651), .D(r_add_B[5]), .E(
        n594), .F(r_x_data[69]), .G(n662), .H(w_mult_2_Z[5]), .Y(n375) );
  scg4d1_hd U1083 ( .A(n681), .B(w_add_Z[6]), .C(n651), .D(r_add_B[6]), .E(
        n607), .F(r_x_data[70]), .G(n662), .H(w_mult_2_Z[6]), .Y(n374) );
  scg4d1_hd U1084 ( .A(n681), .B(w_add_Z[7]), .C(n651), .D(r_add_B[7]), .E(
        n594), .F(r_x_data[71]), .G(n662), .H(w_mult_2_Z[7]), .Y(n373) );
  scg4d1_hd U1085 ( .A(n681), .B(w_add_Z[9]), .C(n651), .D(r_add_B[9]), .E(
        n595), .F(r_x_data[73]), .G(n662), .H(w_mult_2_Z[9]), .Y(n371) );
  scg4d1_hd U1086 ( .A(n682), .B(w_add_Z[14]), .C(n650), .D(r_add_B[14]), .E(
        n608), .F(r_x_data[78]), .G(n661), .H(w_mult_2_Z[14]), .Y(n366) );
  scg4d1_hd U1087 ( .A(n681), .B(w_add_Z[8]), .C(n651), .D(r_add_B[8]), .E(
        n608), .F(r_x_data[72]), .G(n662), .H(w_mult_2_Z[8]), .Y(n372) );
  scg4d1_hd U1088 ( .A(n680), .B(w_add_Z[4]), .C(n651), .D(r_add_B[4]), .E(
        n608), .F(r_x_data[68]), .G(n662), .H(w_mult_2_Z[4]), .Y(n376) );
  scg4d1_hd U1089 ( .A(n682), .B(w_add_Z[13]), .C(n650), .D(r_add_B[13]), .E(
        n595), .F(r_x_data[77]), .G(n661), .H(w_mult_2_Z[13]), .Y(n367) );
  scg4d1_hd U1090 ( .A(n681), .B(w_add_Z[11]), .C(n650), .D(r_add_B[11]), .E(
        n596), .F(r_x_data[75]), .G(n661), .H(w_mult_2_Z[11]), .Y(n369) );
  scg4d1_hd U1091 ( .A(n682), .B(w_add_Z[12]), .C(n650), .D(r_add_B[12]), .E(
        n609), .F(r_x_data[76]), .G(n661), .H(w_mult_2_Z[12]), .Y(n368) );
  scg4d1_hd U1092 ( .A(n682), .B(w_add_Z[15]), .C(n650), .D(r_add_B[15]), .E(
        n610), .F(r_x_data[79]), .G(n661), .H(w_mult_2_Z[15]), .Y(n365) );
  ivd1_hd U1093 ( .A(o_Y_DATA[27]), .Y(n958) );
  ivd1_hd U1094 ( .A(o_Y_DATA[13]), .Y(n916) );
  ivd1_hd U1095 ( .A(o_Y_DATA[14]), .Y(n919) );
  ivd1_hd U1096 ( .A(o_Y_DATA[17]), .Y(n928) );
  ivd1_hd U1097 ( .A(o_Y_DATA[26]), .Y(n955) );
  ivd1_hd U1098 ( .A(o_Y_DATA[18]), .Y(n931) );
  ivd1_hd U1099 ( .A(o_Y_DATA[15]), .Y(n922) );
  ivd1_hd U1100 ( .A(o_Y_DATA[25]), .Y(n952) );
  ivd1_hd U1101 ( .A(o_Y_DATA[16]), .Y(n925) );
  ivd1_hd U1102 ( .A(o_Y_DATA[29]), .Y(n964) );
  ivd1_hd U1103 ( .A(o_Y_DATA[28]), .Y(n961) );
  ivd1_hd U1104 ( .A(o_Y_DATA[30]), .Y(n970) );
  oa21d1_hd U1105 ( .A(n992), .B(n831), .C(n877), .Y(n876) );
  nr2d1_hd U1106 ( .A(n207), .B(n990), .Y(n821) );
  ivd1_hd U1107 ( .A(n164), .Y(n990) );
  scg14d1_hd U1108 ( .A(w_add_Z[11]), .B(n580), .C(n795), .Y(n455) );
  scg14d1_hd U1109 ( .A(w_add_Z[5]), .B(n580), .C(n789), .Y(n461) );
  scg14d1_hd U1110 ( .A(w_add_Z[6]), .B(n580), .C(n790), .Y(n460) );
  scg14d1_hd U1111 ( .A(w_add_Z[7]), .B(n580), .C(n791), .Y(n459) );
  scg14d1_hd U1112 ( .A(w_add_Z[8]), .B(n580), .C(n792), .Y(n458) );
  scg14d1_hd U1113 ( .A(w_add_Z[9]), .B(n581), .C(n793), .Y(n457) );
  scg14d1_hd U1114 ( .A(w_add_Z[10]), .B(n580), .C(n794), .Y(n456) );
  scg14d1_hd U1115 ( .A(w_add_Z[14]), .B(n581), .C(n798), .Y(n452) );
  scg14d1_hd U1116 ( .A(w_add_Z[12]), .B(n581), .C(n796), .Y(n454) );
  scg14d1_hd U1117 ( .A(w_add_Z[13]), .B(n581), .C(n797), .Y(n453) );
  scg14d1_hd U1118 ( .A(w_add_Z[15]), .B(n581), .C(n799), .Y(n451) );
  scg14d1_hd U1119 ( .A(w_add_Z[16]), .B(n581), .C(n800), .Y(n450) );
  nd3d1_hd U1120 ( .A(w_mult_2_AB_ACK), .B(w_add_AB_ACK), .C(w_mult_1_AB_ACK), 
        .Y(n763) );
  ivd1_hd U1121 ( .A(r_pstate_0_), .Y(n760) );
  nd2bd1_hd U1122 ( .AN(r_mult_1_A[6]), .B(n818), .Y(n428) );
  nd2bd1_hd U1123 ( .AN(r_mult_1_A[7]), .B(n818), .Y(n427) );
  nr2d1_hd U1124 ( .A(n207), .B(n164), .Y(n997) );
  ivd1_hd U1125 ( .A(n207), .Y(n992) );
  ivd1_hd U1126 ( .A(n1001), .Y(n991) );
  nd2bd1_hd U1127 ( .AN(r_mult_1_A[3]), .B(n689), .Y(n431) );
  nd2bd1_hd U1128 ( .AN(r_mult_1_A[5]), .B(n689), .Y(n429) );
  ao21d1_hd U1130 ( .A(w_mult_2_Z_STB), .B(w_mult_1_Z_STB), .C(n992), .Y(n996)
         );
  nr2d1_hd U1131 ( .A(n996), .B(n762), .Y(n987) );
  ao211d1_hd U1132 ( .A(i_Y_ACK), .B(o_Y_DATA_VALID), .C(n161), .D(n760), .Y(
        n999) );
  ao211d1_hd U1133 ( .A(n819), .B(n763), .C(n987), .D(n999), .Y(n761) );
  oa21d1_hd U1134 ( .A(n252), .B(n733), .C(n761), .Y(N807) );
  ao22d1_hd U1135 ( .A(n605), .B(r_y_data[12]), .C(r_mult_1_B[12]), .D(n619), 
        .Y(n765) );
  oa21d1_hd U1136 ( .A(n1021), .B(n571), .C(n765), .Y(n485) );
  ao22d1_hd U1137 ( .A(n589), .B(r_y_data[13]), .C(r_mult_1_B[13]), .D(n612), 
        .Y(n766) );
  oa21d1_hd U1138 ( .A(n571), .B(n1020), .C(n766), .Y(n484) );
  ao22d1_hd U1139 ( .A(n601), .B(r_y_data[14]), .C(r_mult_1_B[14]), .D(n612), 
        .Y(n767) );
  oa21d1_hd U1140 ( .A(n572), .B(n1019), .C(n767), .Y(n483) );
  ao22d1_hd U1141 ( .A(n588), .B(r_y_data[15]), .C(r_mult_1_B[15]), .D(n612), 
        .Y(n768) );
  oa21d1_hd U1142 ( .A(n571), .B(n1018), .C(n768), .Y(n482) );
  ao22d1_hd U1143 ( .A(n601), .B(r_y_data[16]), .C(r_mult_1_B[16]), .D(n612), 
        .Y(n769) );
  oa21d1_hd U1144 ( .A(n571), .B(n1017), .C(n769), .Y(n481) );
  ao22d1_hd U1145 ( .A(n588), .B(r_y_data[17]), .C(r_mult_1_B[17]), .D(n612), 
        .Y(n770) );
  oa21d1_hd U1146 ( .A(n571), .B(n1016), .C(n770), .Y(n480) );
  ao22d1_hd U1147 ( .A(n601), .B(r_y_data[18]), .C(r_mult_1_B[18]), .D(n613), 
        .Y(n771) );
  oa21d1_hd U1148 ( .A(n572), .B(n1015), .C(n771), .Y(n479) );
  ao22d1_hd U1149 ( .A(n589), .B(r_y_data[19]), .C(r_mult_1_B[19]), .D(n613), 
        .Y(n772) );
  oa21d1_hd U1150 ( .A(n572), .B(n1014), .C(n772), .Y(n478) );
  ao22d1_hd U1151 ( .A(n601), .B(r_y_data[20]), .C(r_mult_1_B[20]), .D(n613), 
        .Y(n773) );
  oa21d1_hd U1152 ( .A(n572), .B(n1013), .C(n773), .Y(n477) );
  ao22d1_hd U1153 ( .A(n589), .B(r_y_data[21]), .C(r_mult_1_B[21]), .D(n613), 
        .Y(n774) );
  oa21d1_hd U1154 ( .A(n572), .B(n1012), .C(n774), .Y(n476) );
  ao22d1_hd U1155 ( .A(n601), .B(r_y_data[22]), .C(r_mult_1_B[22]), .D(n613), 
        .Y(n775) );
  oa21d1_hd U1156 ( .A(n574), .B(n1011), .C(n775), .Y(n475) );
  ao22d1_hd U1157 ( .A(n589), .B(r_y_data[23]), .C(r_mult_1_B[23]), .D(n613), 
        .Y(n776) );
  oa21d1_hd U1158 ( .A(n572), .B(n1010), .C(n776), .Y(n474) );
  ao22d1_hd U1159 ( .A(n601), .B(r_y_data[24]), .C(r_mult_1_B[24]), .D(n614), 
        .Y(n777) );
  oa21d1_hd U1160 ( .A(n573), .B(n1009), .C(n777), .Y(n473) );
  ao22d1_hd U1161 ( .A(n590), .B(r_y_data[25]), .C(r_mult_1_B[25]), .D(n614), 
        .Y(n778) );
  oa21d1_hd U1162 ( .A(n573), .B(n1008), .C(n778), .Y(n472) );
  ao22d1_hd U1163 ( .A(n602), .B(r_y_data[26]), .C(r_mult_1_B[26]), .D(n614), 
        .Y(n779) );
  oa21d1_hd U1164 ( .A(n573), .B(n1007), .C(n779), .Y(n471) );
  ao22d1_hd U1165 ( .A(n589), .B(r_y_data[27]), .C(r_mult_1_B[27]), .D(n614), 
        .Y(n780) );
  oa21d1_hd U1166 ( .A(n573), .B(n1006), .C(n780), .Y(n470) );
  ao22d1_hd U1167 ( .A(n602), .B(r_y_data[28]), .C(r_mult_1_B[28]), .D(n614), 
        .Y(n781) );
  oa21d1_hd U1168 ( .A(n573), .B(n1005), .C(n781), .Y(n469) );
  ao22d1_hd U1169 ( .A(n590), .B(r_y_data[29]), .C(r_mult_1_B[29]), .D(n614), 
        .Y(n782) );
  oa21d1_hd U1170 ( .A(n573), .B(n1004), .C(n782), .Y(n468) );
  ao22d1_hd U1171 ( .A(n602), .B(r_y_data[30]), .C(r_mult_1_B[30]), .D(n615), 
        .Y(n783) );
  oa21d1_hd U1172 ( .A(n574), .B(n1003), .C(n783), .Y(n467) );
  ao22d1_hd U1173 ( .A(n590), .B(r_y_data[32]), .C(r_mult_2_B[0]), .D(n615), 
        .Y(n784) );
  ao22d1_hd U1174 ( .A(n602), .B(r_y_data[33]), .C(r_mult_2_B[1]), .D(n615), 
        .Y(n785) );
  ao22d1_hd U1175 ( .A(n590), .B(r_y_data[34]), .C(r_mult_2_B[2]), .D(n615), 
        .Y(n786) );
  ao22d1_hd U1176 ( .A(n602), .B(r_y_data[35]), .C(r_mult_2_B[3]), .D(n615), 
        .Y(n787) );
  ao22d1_hd U1177 ( .A(n590), .B(r_y_data[36]), .C(r_mult_2_B[4]), .D(n615), 
        .Y(n788) );
  ao22d1_hd U1178 ( .A(n602), .B(r_y_data[37]), .C(r_mult_2_B[5]), .D(n616), 
        .Y(n789) );
  ao22d1_hd U1179 ( .A(n591), .B(r_y_data[38]), .C(r_mult_2_B[6]), .D(n616), 
        .Y(n790) );
  ao22d1_hd U1180 ( .A(n603), .B(r_y_data[39]), .C(r_mult_2_B[7]), .D(n616), 
        .Y(n791) );
  ao22d1_hd U1181 ( .A(n590), .B(r_y_data[40]), .C(r_mult_2_B[8]), .D(n616), 
        .Y(n792) );
  ao22d1_hd U1182 ( .A(n603), .B(r_y_data[41]), .C(r_mult_2_B[9]), .D(n616), 
        .Y(n793) );
  ao22d1_hd U1183 ( .A(n591), .B(r_y_data[42]), .C(r_mult_2_B[10]), .D(n616), 
        .Y(n794) );
  ao22d1_hd U1184 ( .A(n603), .B(r_y_data[43]), .C(r_mult_2_B[11]), .D(n617), 
        .Y(n795) );
  ao22d1_hd U1185 ( .A(n592), .B(r_y_data[44]), .C(r_mult_2_B[12]), .D(n617), 
        .Y(n796) );
  ao22d1_hd U1186 ( .A(n603), .B(r_y_data[45]), .C(r_mult_2_B[13]), .D(n617), 
        .Y(n797) );
  ao22d1_hd U1187 ( .A(n591), .B(r_y_data[46]), .C(r_mult_2_B[14]), .D(n617), 
        .Y(n798) );
  ao22d1_hd U1188 ( .A(n603), .B(r_y_data[47]), .C(r_mult_2_B[15]), .D(n617), 
        .Y(n799) );
  ao22d1_hd U1189 ( .A(n591), .B(r_y_data[48]), .C(r_mult_2_B[16]), .D(n617), 
        .Y(n800) );
  ao22d1_hd U1190 ( .A(n603), .B(r_y_data[49]), .C(r_mult_2_B[17]), .D(n618), 
        .Y(n801) );
  ao22d1_hd U1191 ( .A(n591), .B(r_y_data[50]), .C(r_mult_2_B[18]), .D(n618), 
        .Y(n802) );
  ao22d1_hd U1192 ( .A(n604), .B(r_y_data[51]), .C(r_mult_2_B[19]), .D(n618), 
        .Y(n803) );
  ao22d1_hd U1193 ( .A(n591), .B(r_y_data[52]), .C(r_mult_2_B[20]), .D(n618), 
        .Y(n804) );
  ao22d1_hd U1194 ( .A(n604), .B(r_y_data[53]), .C(r_mult_2_B[21]), .D(n618), 
        .Y(n805) );
  ao22d1_hd U1195 ( .A(n592), .B(r_y_data[54]), .C(r_mult_2_B[22]), .D(n618), 
        .Y(n806) );
  ao22d1_hd U1196 ( .A(n604), .B(r_y_data[55]), .C(r_mult_2_B[23]), .D(n619), 
        .Y(n807) );
  ao22d1_hd U1197 ( .A(n592), .B(r_y_data[56]), .C(r_mult_2_B[24]), .D(n619), 
        .Y(n808) );
  ao22d1_hd U1198 ( .A(n604), .B(r_y_data[57]), .C(r_mult_2_B[25]), .D(n619), 
        .Y(n809) );
  scg14d1_hd U1199 ( .A(w_add_Z[25]), .B(n585), .C(n809), .Y(n441) );
  ao22d1_hd U1200 ( .A(n592), .B(r_y_data[58]), .C(r_mult_2_B[26]), .D(n619), 
        .Y(n810) );
  scg14d1_hd U1201 ( .A(w_add_Z[26]), .B(n585), .C(n810), .Y(n440) );
  ao22d1_hd U1202 ( .A(n604), .B(r_y_data[59]), .C(r_mult_2_B[27]), .D(n619), 
        .Y(n811) );
  scg14d1_hd U1203 ( .A(w_add_Z[27]), .B(n585), .C(n811), .Y(n439) );
  ao22d1_hd U1204 ( .A(n592), .B(r_y_data[60]), .C(r_mult_2_B[28]), .D(n620), 
        .Y(n812) );
  scg14d1_hd U1205 ( .A(w_add_Z[28]), .B(n585), .C(n812), .Y(n438) );
  ao22d1_hd U1206 ( .A(n604), .B(r_y_data[61]), .C(r_mult_2_B[29]), .D(n620), 
        .Y(n813) );
  scg14d1_hd U1207 ( .A(w_add_Z[29]), .B(n585), .C(n813), .Y(n437) );
  ao22d1_hd U1208 ( .A(n592), .B(r_y_data[62]), .C(r_mult_2_B[30]), .D(n620), 
        .Y(n814) );
  ivd1_hd U1209 ( .A(r_mult_AB_STB), .Y(n815) );
  oa22d1_hd U1210 ( .A(n992), .B(n817), .C(n816), .D(n815), .Y(n435) );
  nd2bd1_hd U1211 ( .AN(r_mult_1_A[10]), .B(n631), .Y(n424) );
  nd2bd1_hd U1212 ( .AN(r_mult_1_A[11]), .B(n631), .Y(n423) );
  nd2bd1_hd U1213 ( .AN(r_mult_1_A[17]), .B(n631), .Y(n418) );
  nd2bd1_hd U1214 ( .AN(r_mult_1_A[20]), .B(n631), .Y(n416) );
  nd2bd1_hd U1215 ( .AN(r_mult_1_A[22]), .B(n631), .Y(n415) );
  nd2bd1_hd U1216 ( .AN(r_mult_1_A[23]), .B(n631), .Y(n414) );
  nd2bd1_hd U1217 ( .AN(r_mult_1_A[26]), .B(n630), .Y(n411) );
  nd2bd1_hd U1218 ( .AN(r_mult_1_A[27]), .B(n630), .Y(n410) );
  nd2bd1_hd U1219 ( .AN(r_mult_1_A[28]), .B(n630), .Y(n409) );
  nd2bd1_hd U1220 ( .AN(r_mult_1_A[29]), .B(n630), .Y(n408) );
  nd2bd1_hd U1221 ( .AN(r_mult_2_A[0]), .B(n630), .Y(n407) );
  nd2bd1_hd U1222 ( .AN(r_mult_2_A[3]), .B(n630), .Y(n404) );
  nd2bd1_hd U1223 ( .AN(r_mult_2_A[5]), .B(n629), .Y(n402) );
  nd2bd1_hd U1224 ( .AN(r_mult_2_A[6]), .B(n629), .Y(n401) );
  nd2bd1_hd U1225 ( .AN(r_mult_2_A[7]), .B(n629), .Y(n400) );
  nd2bd1_hd U1226 ( .AN(r_mult_2_A[10]), .B(n629), .Y(n398) );
  nd2bd1_hd U1227 ( .AN(r_mult_2_A[11]), .B(n629), .Y(n397) );
  nd2bd1_hd U1228 ( .AN(r_mult_2_A[16]), .B(n629), .Y(n394) );
  nd2bd1_hd U1229 ( .AN(r_mult_2_A[17]), .B(n628), .Y(n393) );
  nd2bd1_hd U1230 ( .AN(r_mult_2_A[20]), .B(n628), .Y(n391) );
  nd2bd1_hd U1231 ( .AN(r_mult_2_A[26]), .B(n628), .Y(n386) );
  nd2bd1_hd U1232 ( .AN(r_mult_2_A[27]), .B(n628), .Y(n385) );
  nd2bd1_hd U1233 ( .AN(r_mult_2_A[28]), .B(n628), .Y(n384) );
  nd2bd1_hd U1234 ( .AN(r_mult_2_A[29]), .B(n628), .Y(n383) );
  oa21d1_hd U1235 ( .A(n819), .B(n1001), .C(o_Y_DATA_VALID), .Y(n820) );
  nd2bd1_hd U1236 ( .AN(n999), .B(n820), .Y(n381) );
  ao22d1_hd U1237 ( .A(r_x_data[0]), .B(n611), .C(r_add_A[0]), .D(n647), .Y(
        n828) );
  ao22d1_hd U1238 ( .A(n658), .B(w_mult_1_Z[0]), .C(w_mult_2_Z[0]), .D(n632), 
        .Y(n827) );
  oa211d1_hd U1239 ( .A(n637), .B(n840), .C(n828), .D(n827), .Y(n568) );
  ao22d1_hd U1240 ( .A(r_x_data[31]), .B(n600), .C(r_add_A[31]), .D(n647), .Y(
        n830) );
  ao22d1_hd U1241 ( .A(n658), .B(w_mult_1_Z[31]), .C(n632), .D(w_mult_2_Z[31]), 
        .Y(n829) );
  oa211d1_hd U1242 ( .A(n637), .B(n837), .C(n830), .D(n829), .Y(n567) );
  ao22d1_hd U1243 ( .A(w_add_Z[31]), .B(n695), .C(w_mult_1_Z[31]), .D(n679), 
        .Y(n836) );
  oa21d1_hd U1244 ( .A(n837), .B(n664), .C(n836), .Y(n566) );
  ao22d1_hd U1245 ( .A(n605), .B(r_y_data[31]), .C(r_mult_1_B[31]), .D(n620), 
        .Y(n838) );
  oa21d1_hd U1246 ( .A(n574), .B(n1002), .C(n838), .Y(n565) );
  ao22d1_hd U1247 ( .A(w_add_Z[0]), .B(n871), .C(w_mult_1_Z[0]), .D(n679), .Y(
        n839) );
  oa21d1_hd U1248 ( .A(n840), .B(n664), .C(n839), .Y(n564) );
  ao22d1_hd U1249 ( .A(w_add_Z[1]), .B(n673), .C(w_mult_1_Z[1]), .D(n678), .Y(
        n841) );
  oa21d1_hd U1250 ( .A(n880), .B(n664), .C(n841), .Y(n563) );
  ao22d1_hd U1251 ( .A(w_add_Z[2]), .B(n673), .C(w_mult_1_Z[2]), .D(n678), .Y(
        n842) );
  oa21d1_hd U1252 ( .A(n883), .B(n664), .C(n842), .Y(n562) );
  ao22d1_hd U1253 ( .A(w_add_Z[3]), .B(n673), .C(w_mult_1_Z[3]), .D(n678), .Y(
        n843) );
  oa21d1_hd U1254 ( .A(n886), .B(n664), .C(n843), .Y(n561) );
  ao22d1_hd U1255 ( .A(w_add_Z[4]), .B(n673), .C(w_mult_1_Z[4]), .D(n678), .Y(
        n844) );
  oa21d1_hd U1256 ( .A(n889), .B(n665), .C(n844), .Y(n560) );
  ao22d1_hd U1257 ( .A(w_add_Z[5]), .B(n673), .C(w_mult_1_Z[5]), .D(n678), .Y(
        n845) );
  oa21d1_hd U1258 ( .A(n892), .B(n665), .C(n845), .Y(n559) );
  ao22d1_hd U1259 ( .A(w_add_Z[6]), .B(n673), .C(w_mult_1_Z[6]), .D(n678), .Y(
        n846) );
  oa21d1_hd U1260 ( .A(n895), .B(n665), .C(n846), .Y(n558) );
  ao22d1_hd U1261 ( .A(w_add_Z[7]), .B(n672), .C(w_mult_1_Z[7]), .D(n677), .Y(
        n847) );
  oa21d1_hd U1262 ( .A(n898), .B(n665), .C(n847), .Y(n557) );
  ao22d1_hd U1263 ( .A(w_add_Z[8]), .B(n672), .C(w_mult_1_Z[8]), .D(n677), .Y(
        n848) );
  oa21d1_hd U1264 ( .A(n901), .B(n665), .C(n848), .Y(n556) );
  ao22d1_hd U1265 ( .A(w_add_Z[9]), .B(n672), .C(w_mult_1_Z[9]), .D(n677), .Y(
        n849) );
  oa21d1_hd U1266 ( .A(n904), .B(n665), .C(n849), .Y(n555) );
  ao22d1_hd U1267 ( .A(w_add_Z[10]), .B(n672), .C(w_mult_1_Z[10]), .D(n677), 
        .Y(n850) );
  oa21d1_hd U1268 ( .A(n907), .B(n666), .C(n850), .Y(n554) );
  ao22d1_hd U1269 ( .A(w_add_Z[11]), .B(n672), .C(w_mult_1_Z[11]), .D(n677), 
        .Y(n851) );
  oa21d1_hd U1270 ( .A(n910), .B(n666), .C(n851), .Y(n553) );
  ao22d1_hd U1271 ( .A(w_add_Z[12]), .B(n672), .C(w_mult_1_Z[12]), .D(n677), 
        .Y(n852) );
  oa21d1_hd U1272 ( .A(n913), .B(n666), .C(n852), .Y(n552) );
  ao22d1_hd U1273 ( .A(w_add_Z[13]), .B(n671), .C(w_mult_1_Z[13]), .D(n676), 
        .Y(n853) );
  oa21d1_hd U1274 ( .A(n916), .B(n666), .C(n853), .Y(n551) );
  ao22d1_hd U1275 ( .A(w_add_Z[14]), .B(n671), .C(w_mult_1_Z[14]), .D(n676), 
        .Y(n854) );
  oa21d1_hd U1276 ( .A(n919), .B(n666), .C(n854), .Y(n550) );
  ao22d1_hd U1277 ( .A(w_add_Z[15]), .B(n671), .C(w_mult_1_Z[15]), .D(n676), 
        .Y(n855) );
  oa21d1_hd U1278 ( .A(n922), .B(n666), .C(n855), .Y(n549) );
  ao22d1_hd U1279 ( .A(w_add_Z[16]), .B(n671), .C(w_mult_1_Z[16]), .D(n676), 
        .Y(n856) );
  oa21d1_hd U1280 ( .A(n925), .B(n667), .C(n856), .Y(n548) );
  ao22d1_hd U1281 ( .A(w_add_Z[17]), .B(n671), .C(w_mult_1_Z[17]), .D(n676), 
        .Y(n857) );
  oa21d1_hd U1282 ( .A(n928), .B(n667), .C(n857), .Y(n547) );
  ao22d1_hd U1283 ( .A(w_add_Z[18]), .B(n671), .C(w_mult_1_Z[18]), .D(n676), 
        .Y(n858) );
  oa21d1_hd U1284 ( .A(n931), .B(n667), .C(n858), .Y(n546) );
  ao22d1_hd U1285 ( .A(w_add_Z[19]), .B(n670), .C(w_mult_1_Z[19]), .D(n675), 
        .Y(n859) );
  oa21d1_hd U1286 ( .A(n934), .B(n667), .C(n859), .Y(n545) );
  ao22d1_hd U1287 ( .A(w_add_Z[20]), .B(n670), .C(w_mult_1_Z[20]), .D(n675), 
        .Y(n860) );
  oa21d1_hd U1288 ( .A(n937), .B(n667), .C(n860), .Y(n544) );
  ao22d1_hd U1289 ( .A(w_add_Z[21]), .B(n670), .C(w_mult_1_Z[21]), .D(n675), 
        .Y(n861) );
  oa21d1_hd U1290 ( .A(n940), .B(n667), .C(n861), .Y(n543) );
  ao22d1_hd U1291 ( .A(w_add_Z[22]), .B(n670), .C(w_mult_1_Z[22]), .D(n675), 
        .Y(n862) );
  oa21d1_hd U1292 ( .A(n943), .B(n668), .C(n862), .Y(n542) );
  ao22d1_hd U1293 ( .A(w_add_Z[23]), .B(n670), .C(w_mult_1_Z[23]), .D(n675), 
        .Y(n863) );
  oa21d1_hd U1294 ( .A(n946), .B(n668), .C(n863), .Y(n541) );
  ao22d1_hd U1295 ( .A(w_add_Z[24]), .B(n670), .C(w_mult_1_Z[24]), .D(n675), 
        .Y(n864) );
  oa21d1_hd U1296 ( .A(n949), .B(n668), .C(n864), .Y(n540) );
  ao22d1_hd U1297 ( .A(w_add_Z[25]), .B(n669), .C(w_mult_1_Z[25]), .D(n674), 
        .Y(n865) );
  oa21d1_hd U1298 ( .A(n952), .B(n668), .C(n865), .Y(n539) );
  ao22d1_hd U1299 ( .A(w_add_Z[26]), .B(n669), .C(w_mult_1_Z[26]), .D(n674), 
        .Y(n866) );
  oa21d1_hd U1300 ( .A(n955), .B(n668), .C(n866), .Y(n538) );
  ao22d1_hd U1301 ( .A(w_add_Z[27]), .B(n669), .C(w_mult_1_Z[27]), .D(n674), 
        .Y(n867) );
  oa21d1_hd U1302 ( .A(n958), .B(n668), .C(n867), .Y(n537) );
  ao22d1_hd U1303 ( .A(w_add_Z[28]), .B(n669), .C(w_mult_1_Z[28]), .D(n674), 
        .Y(n868) );
  oa21d1_hd U1304 ( .A(n961), .B(n873), .C(n868), .Y(n536) );
  ao22d1_hd U1305 ( .A(w_add_Z[29]), .B(n669), .C(w_mult_1_Z[29]), .D(n674), 
        .Y(n869) );
  oa21d1_hd U1306 ( .A(n964), .B(n873), .C(n869), .Y(n535) );
  ao22d1_hd U1307 ( .A(w_add_Z[30]), .B(n669), .C(w_mult_1_Z[30]), .D(n674), 
        .Y(n872) );
  oa21d1_hd U1308 ( .A(n970), .B(n694), .C(n872), .Y(n534) );
  ao22d1_hd U1309 ( .A(n593), .B(r_y_data[63]), .C(r_mult_2_B[31]), .D(n621), 
        .Y(n874) );
  scg14d1_hd U1310 ( .A(r_add_AB_STB), .B(n991), .C(n875), .Y(n532) );
  ao22ad1_hd U1311 ( .A(n991), .B(n876), .C(n876), .D(r_mult_Z_ACK), .Y(n529)
         );
  scg6d1_hd U1312 ( .A(r_add_Z_ACK), .B(n877), .C(n987), .Y(n528) );
  ao22d1_hd U1313 ( .A(r_x_data[1]), .B(n588), .C(r_add_A[1]), .D(n646), .Y(
        n879) );
  ao22d1_hd U1314 ( .A(n657), .B(w_mult_1_Z[1]), .C(n632), .D(w_mult_2_Z[1]), 
        .Y(n878) );
  oa211d1_hd U1315 ( .A(n637), .B(n880), .C(n879), .D(n878), .Y(n527) );
  ao22d1_hd U1316 ( .A(r_x_data[2]), .B(n599), .C(r_add_A[2]), .D(n646), .Y(
        n882) );
  ao22d1_hd U1317 ( .A(n657), .B(w_mult_1_Z[2]), .C(n632), .D(w_mult_2_Z[2]), 
        .Y(n881) );
  oa211d1_hd U1318 ( .A(n637), .B(n883), .C(n882), .D(n881), .Y(n526) );
  ao22d1_hd U1319 ( .A(r_x_data[3]), .B(n587), .C(r_add_A[3]), .D(n646), .Y(
        n885) );
  ao22d1_hd U1320 ( .A(n657), .B(w_mult_1_Z[3]), .C(n632), .D(w_mult_2_Z[3]), 
        .Y(n884) );
  oa211d1_hd U1321 ( .A(n637), .B(n886), .C(n885), .D(n884), .Y(n525) );
  ao22d1_hd U1322 ( .A(r_x_data[4]), .B(n600), .C(r_add_A[4]), .D(n646), .Y(
        n888) );
  ao22d1_hd U1323 ( .A(n657), .B(w_mult_1_Z[4]), .C(n633), .D(w_mult_2_Z[4]), 
        .Y(n887) );
  oa211d1_hd U1324 ( .A(n638), .B(n889), .C(n888), .D(n887), .Y(n524) );
  ao22d1_hd U1325 ( .A(r_x_data[5]), .B(n588), .C(r_add_A[5]), .D(n646), .Y(
        n891) );
  ao22d1_hd U1326 ( .A(n657), .B(w_mult_1_Z[5]), .C(n633), .D(w_mult_2_Z[5]), 
        .Y(n890) );
  oa211d1_hd U1327 ( .A(n638), .B(n892), .C(n891), .D(n890), .Y(n523) );
  ao22d1_hd U1328 ( .A(r_x_data[6]), .B(n600), .C(r_add_A[6]), .D(n646), .Y(
        n894) );
  ao22d1_hd U1329 ( .A(n657), .B(w_mult_1_Z[6]), .C(n633), .D(w_mult_2_Z[6]), 
        .Y(n893) );
  oa211d1_hd U1330 ( .A(n638), .B(n895), .C(n894), .D(n893), .Y(n522) );
  ao22d1_hd U1331 ( .A(r_x_data[7]), .B(n588), .C(r_add_A[7]), .D(n645), .Y(
        n897) );
  ao22d1_hd U1332 ( .A(n656), .B(w_mult_1_Z[7]), .C(n633), .D(w_mult_2_Z[7]), 
        .Y(n896) );
  oa211d1_hd U1333 ( .A(n638), .B(n898), .C(n897), .D(n896), .Y(n521) );
  ao22d1_hd U1334 ( .A(r_x_data[8]), .B(n599), .C(r_add_A[8]), .D(n645), .Y(
        n900) );
  ao22d1_hd U1335 ( .A(n656), .B(w_mult_1_Z[8]), .C(n633), .D(w_mult_2_Z[8]), 
        .Y(n899) );
  oa211d1_hd U1336 ( .A(n638), .B(n901), .C(n900), .D(n899), .Y(n520) );
  ao22d1_hd U1337 ( .A(r_x_data[9]), .B(n586), .C(r_add_A[9]), .D(n645), .Y(
        n903) );
  ao22d1_hd U1338 ( .A(n656), .B(w_mult_1_Z[9]), .C(n633), .D(w_mult_2_Z[9]), 
        .Y(n902) );
  oa211d1_hd U1339 ( .A(n638), .B(n904), .C(n903), .D(n902), .Y(n519) );
  ao22d1_hd U1340 ( .A(r_x_data[10]), .B(n600), .C(r_add_A[10]), .D(n645), .Y(
        n906) );
  ao22d1_hd U1341 ( .A(n656), .B(w_mult_1_Z[10]), .C(n634), .D(w_mult_2_Z[10]), 
        .Y(n905) );
  oa211d1_hd U1342 ( .A(n639), .B(n907), .C(n906), .D(n905), .Y(n518) );
  ao22d1_hd U1343 ( .A(r_x_data[11]), .B(n600), .C(r_add_A[11]), .D(n645), .Y(
        n909) );
  ao22d1_hd U1344 ( .A(n656), .B(w_mult_1_Z[11]), .C(n634), .D(w_mult_2_Z[11]), 
        .Y(n908) );
  oa211d1_hd U1345 ( .A(n639), .B(n910), .C(n909), .D(n908), .Y(n517) );
  ao22d1_hd U1346 ( .A(r_x_data[12]), .B(n588), .C(r_add_A[12]), .D(n645), .Y(
        n912) );
  ao22d1_hd U1347 ( .A(n656), .B(w_mult_1_Z[12]), .C(n634), .D(w_mult_2_Z[12]), 
        .Y(n911) );
  oa211d1_hd U1348 ( .A(n639), .B(n913), .C(n912), .D(n911), .Y(n516) );
  ao22d1_hd U1349 ( .A(r_x_data[13]), .B(n599), .C(r_add_A[13]), .D(n644), .Y(
        n915) );
  ao22d1_hd U1350 ( .A(n655), .B(w_mult_1_Z[13]), .C(n634), .D(w_mult_2_Z[13]), 
        .Y(n914) );
  oa211d1_hd U1351 ( .A(n639), .B(n916), .C(n915), .D(n914), .Y(n515) );
  ao22d1_hd U1352 ( .A(r_x_data[14]), .B(n587), .C(r_add_A[14]), .D(n644), .Y(
        n918) );
  ao22d1_hd U1353 ( .A(n655), .B(w_mult_1_Z[14]), .C(n634), .D(w_mult_2_Z[14]), 
        .Y(n917) );
  oa211d1_hd U1354 ( .A(n639), .B(n919), .C(n918), .D(n917), .Y(n514) );
  ao22d1_hd U1355 ( .A(r_x_data[15]), .B(n599), .C(r_add_A[15]), .D(n644), .Y(
        n921) );
  ao22d1_hd U1356 ( .A(n655), .B(w_mult_1_Z[15]), .C(n634), .D(w_mult_2_Z[15]), 
        .Y(n920) );
  oa211d1_hd U1357 ( .A(n639), .B(n922), .C(n921), .D(n920), .Y(n513) );
  ao22d1_hd U1358 ( .A(r_x_data[16]), .B(n587), .C(r_add_A[16]), .D(n644), .Y(
        n924) );
  ao22d1_hd U1359 ( .A(n655), .B(w_mult_1_Z[16]), .C(n635), .D(w_mult_2_Z[16]), 
        .Y(n923) );
  oa211d1_hd U1360 ( .A(n640), .B(n925), .C(n924), .D(n923), .Y(n512) );
  ao22d1_hd U1361 ( .A(r_x_data[17]), .B(n599), .C(r_add_A[17]), .D(n644), .Y(
        n927) );
  ao22d1_hd U1362 ( .A(n655), .B(w_mult_1_Z[17]), .C(n635), .D(w_mult_2_Z[17]), 
        .Y(n926) );
  oa211d1_hd U1363 ( .A(n640), .B(n928), .C(n927), .D(n926), .Y(n511) );
  ao22d1_hd U1364 ( .A(r_x_data[18]), .B(n587), .C(r_add_A[18]), .D(n644), .Y(
        n930) );
  ao22d1_hd U1365 ( .A(n655), .B(w_mult_1_Z[18]), .C(n635), .D(w_mult_2_Z[18]), 
        .Y(n929) );
  oa211d1_hd U1366 ( .A(n640), .B(n931), .C(n930), .D(n929), .Y(n510) );
  ao22d1_hd U1367 ( .A(r_x_data[19]), .B(n687), .C(r_add_A[19]), .D(n643), .Y(
        n933) );
  ao22d1_hd U1368 ( .A(n654), .B(w_mult_1_Z[19]), .C(n635), .D(w_mult_2_Z[19]), 
        .Y(n932) );
  oa211d1_hd U1369 ( .A(n640), .B(n934), .C(n933), .D(n932), .Y(n509) );
  ao22d1_hd U1370 ( .A(r_x_data[20]), .B(n587), .C(r_add_A[20]), .D(n643), .Y(
        n936) );
  ao22d1_hd U1371 ( .A(n654), .B(w_mult_1_Z[20]), .C(n635), .D(w_mult_2_Z[20]), 
        .Y(n935) );
  oa211d1_hd U1372 ( .A(n640), .B(n937), .C(n936), .D(n935), .Y(n508) );
  ao22d1_hd U1373 ( .A(r_x_data[21]), .B(n599), .C(r_add_A[21]), .D(n643), .Y(
        n939) );
  ao22d1_hd U1374 ( .A(n654), .B(w_mult_1_Z[21]), .C(n635), .D(w_mult_2_Z[21]), 
        .Y(n938) );
  oa211d1_hd U1375 ( .A(n640), .B(n940), .C(n939), .D(n938), .Y(n507) );
  ao22d1_hd U1376 ( .A(r_x_data[22]), .B(n586), .C(r_add_A[22]), .D(n643), .Y(
        n942) );
  ao22d1_hd U1377 ( .A(n654), .B(w_mult_1_Z[22]), .C(n636), .D(w_mult_2_Z[22]), 
        .Y(n941) );
  oa211d1_hd U1378 ( .A(n641), .B(n943), .C(n942), .D(n941), .Y(n506) );
  ao22d1_hd U1379 ( .A(r_x_data[23]), .B(n611), .C(r_add_A[23]), .D(n643), .Y(
        n945) );
  ao22d1_hd U1380 ( .A(n654), .B(w_mult_1_Z[23]), .C(n636), .D(w_mult_2_Z[23]), 
        .Y(n944) );
  oa211d1_hd U1381 ( .A(n641), .B(n946), .C(n945), .D(n944), .Y(n505) );
  ao22d1_hd U1382 ( .A(r_x_data[24]), .B(n587), .C(r_add_A[24]), .D(n643), .Y(
        n948) );
  ao22d1_hd U1383 ( .A(n654), .B(w_mult_1_Z[24]), .C(n636), .D(w_mult_2_Z[24]), 
        .Y(n947) );
  oa211d1_hd U1384 ( .A(n641), .B(n949), .C(n948), .D(n947), .Y(n504) );
  ao22d1_hd U1385 ( .A(r_x_data[25]), .B(n687), .C(r_add_A[25]), .D(n642), .Y(
        n951) );
  ao22d1_hd U1386 ( .A(n653), .B(w_mult_1_Z[25]), .C(n636), .D(w_mult_2_Z[25]), 
        .Y(n950) );
  oa211d1_hd U1387 ( .A(n641), .B(n952), .C(n951), .D(n950), .Y(n503) );
  ao22d1_hd U1388 ( .A(r_x_data[26]), .B(n586), .C(r_add_A[26]), .D(n642), .Y(
        n954) );
  ao22d1_hd U1389 ( .A(n653), .B(w_mult_1_Z[26]), .C(n636), .D(w_mult_2_Z[26]), 
        .Y(n953) );
  oa211d1_hd U1390 ( .A(n641), .B(n955), .C(n954), .D(n953), .Y(n502) );
  ao22d1_hd U1391 ( .A(r_x_data[27]), .B(n687), .C(r_add_A[27]), .D(n642), .Y(
        n957) );
  ao22d1_hd U1392 ( .A(n653), .B(w_mult_1_Z[27]), .C(n636), .D(w_mult_2_Z[27]), 
        .Y(n956) );
  oa211d1_hd U1393 ( .A(n641), .B(n958), .C(n957), .D(n956), .Y(n501) );
  ao22d1_hd U1394 ( .A(r_x_data[28]), .B(n586), .C(r_add_A[28]), .D(n642), .Y(
        n960) );
  ao22d1_hd U1395 ( .A(n653), .B(w_mult_1_Z[28]), .C(n966), .D(w_mult_2_Z[28]), 
        .Y(n959) );
  oa211d1_hd U1396 ( .A(n971), .B(n961), .C(n960), .D(n959), .Y(n500) );
  ao22d1_hd U1397 ( .A(r_x_data[29]), .B(n611), .C(r_add_A[29]), .D(n642), .Y(
        n963) );
  ao22d1_hd U1398 ( .A(n653), .B(w_mult_1_Z[29]), .C(n966), .D(w_mult_2_Z[29]), 
        .Y(n962) );
  oa211d1_hd U1399 ( .A(n971), .B(n964), .C(n963), .D(n962), .Y(n499) );
  ao22d1_hd U1400 ( .A(r_x_data[30]), .B(n586), .C(r_add_A[30]), .D(n642), .Y(
        n969) );
  ao22d1_hd U1401 ( .A(n653), .B(w_mult_1_Z[30]), .C(n690), .D(w_mult_2_Z[30]), 
        .Y(n968) );
  oa211d1_hd U1402 ( .A(n691), .B(n970), .C(n969), .D(n968), .Y(n498) );
  ao22d1_hd U1403 ( .A(n605), .B(r_y_data[0]), .C(r_mult_1_B[0]), .D(n621), 
        .Y(n972) );
  oa21d1_hd U1404 ( .A(n575), .B(n1033), .C(n972), .Y(n497) );
  ao22d1_hd U1405 ( .A(n593), .B(r_y_data[1]), .C(r_mult_1_B[1]), .D(n620), 
        .Y(n973) );
  oa21d1_hd U1406 ( .A(n574), .B(n1032), .C(n973), .Y(n496) );
  ao22d1_hd U1407 ( .A(n605), .B(r_y_data[2]), .C(r_mult_1_B[2]), .D(n621), 
        .Y(n974) );
  oa21d1_hd U1408 ( .A(n574), .B(n1031), .C(n974), .Y(n495) );
  ao22d1_hd U1409 ( .A(n593), .B(r_y_data[3]), .C(r_mult_1_B[3]), .D(n621), 
        .Y(n975) );
  oa21d1_hd U1410 ( .A(n575), .B(n1030), .C(n975), .Y(n494) );
  ao22d1_hd U1411 ( .A(n605), .B(r_y_data[4]), .C(r_mult_1_B[4]), .D(n621), 
        .Y(n976) );
  oa21d1_hd U1412 ( .A(n575), .B(n1029), .C(n976), .Y(n493) );
  ao22d1_hd U1413 ( .A(n593), .B(r_y_data[5]), .C(r_mult_1_B[5]), .D(n622), 
        .Y(n977) );
  oa21d1_hd U1414 ( .A(n575), .B(n1028), .C(n977), .Y(n492) );
  ao22d1_hd U1415 ( .A(n606), .B(r_y_data[6]), .C(r_mult_1_B[6]), .D(n621), 
        .Y(n978) );
  oa21d1_hd U1416 ( .A(n574), .B(n1027), .C(n978), .Y(n491) );
  ao22d1_hd U1417 ( .A(n593), .B(r_y_data[7]), .C(r_mult_1_B[7]), .D(n622), 
        .Y(n979) );
  oa21d1_hd U1418 ( .A(n575), .B(n1026), .C(n979), .Y(n490) );
  ao22d1_hd U1419 ( .A(n605), .B(r_y_data[8]), .C(r_mult_1_B[8]), .D(n622), 
        .Y(n980) );
  oa21d1_hd U1420 ( .A(n576), .B(n1025), .C(n980), .Y(n489) );
  ao22d1_hd U1421 ( .A(n593), .B(r_y_data[9]), .C(r_mult_1_B[9]), .D(n622), 
        .Y(n981) );
  oa21d1_hd U1422 ( .A(n576), .B(n1024), .C(n981), .Y(n488) );
  ao22d1_hd U1423 ( .A(n600), .B(r_y_data[10]), .C(r_mult_1_B[10]), .D(n620), 
        .Y(n982) );
  oa21d1_hd U1424 ( .A(n575), .B(n1023), .C(n982), .Y(n487) );
  ao22d1_hd U1425 ( .A(n589), .B(r_y_data[11]), .C(r_mult_1_B[11]), .D(n612), 
        .Y(n985) );
  oa21d1_hd U1426 ( .A(n571), .B(n1022), .C(n985), .Y(n486) );
  nr2d1_hd U1427 ( .A(n995), .B(n991), .Y(n989) );
  nr2d1_hd U1428 ( .A(n164), .B(n995), .Y(n993) );
  ivd1_hd U1429 ( .A(n993), .Y(n988) );
  oa21d1_hd U1430 ( .A(n990), .B(n989), .C(n988), .Y(n163) );
  nr2d1_hd U1431 ( .A(n997), .B(n991), .Y(n994) );
  oa22d1_hd U1432 ( .A(n995), .B(n994), .C(n993), .D(n992), .Y(n162) );
  scg13d1_hd U1433 ( .A(n997), .B(n996), .C(w_add_Z_STB), .Y(n1000) );
  ao211d1_hd U1434 ( .A(n1001), .B(n1000), .C(n999), .D(n998), .Y(n160) );
  ao22d1_hd U1435 ( .A(n707), .B(n1035), .C(n1002), .D(n733), .Y(n96) );
  ao22d1_hd U1436 ( .A(n707), .B(n1037), .C(n1003), .D(n732), .Y(n97) );
  ao22d1_hd U1437 ( .A(n707), .B(n1039), .C(n1004), .D(n732), .Y(n98) );
  ao22d1_hd U1438 ( .A(n707), .B(n1041), .C(n1005), .D(n732), .Y(n99) );
  ao22d1_hd U1439 ( .A(n706), .B(n1043), .C(n1006), .D(n569), .Y(n100) );
  ao22d1_hd U1440 ( .A(n706), .B(n1045), .C(n1007), .D(n757), .Y(n101) );
  ao22d1_hd U1441 ( .A(n706), .B(n1047), .C(n1008), .D(n737), .Y(n102) );
  ao22d1_hd U1442 ( .A(n706), .B(n1049), .C(n1009), .D(n737), .Y(n103) );
  ao22d1_hd U1443 ( .A(n706), .B(n1051), .C(n1010), .D(n737), .Y(n104) );
  ao22d1_hd U1444 ( .A(n706), .B(n1053), .C(n1011), .D(n737), .Y(n105) );
  ao22d1_hd U1445 ( .A(n705), .B(n1055), .C(n1012), .D(n737), .Y(n106) );
  ao22d1_hd U1446 ( .A(n705), .B(n1057), .C(n1013), .D(n737), .Y(n107) );
  ao22d1_hd U1447 ( .A(n705), .B(n1059), .C(n1014), .D(n736), .Y(n108) );
  ao22d1_hd U1448 ( .A(n705), .B(n1061), .C(n1015), .D(n736), .Y(n109) );
  ao22d1_hd U1449 ( .A(n705), .B(n1063), .C(n1016), .D(n736), .Y(n110) );
  ao22d1_hd U1450 ( .A(n705), .B(n1065), .C(n1017), .D(n736), .Y(n111) );
  ao22d1_hd U1451 ( .A(n704), .B(n1067), .C(n1018), .D(n736), .Y(n112) );
  ao22d1_hd U1452 ( .A(n704), .B(n1069), .C(n1019), .D(n736), .Y(n113) );
  ao22d1_hd U1453 ( .A(n704), .B(n1071), .C(n1020), .D(n735), .Y(n114) );
  ao22d1_hd U1454 ( .A(n704), .B(n1073), .C(n1021), .D(n735), .Y(n115) );
  ao22d1_hd U1455 ( .A(n704), .B(n1075), .C(n1022), .D(n735), .Y(n116) );
  ao22d1_hd U1456 ( .A(n704), .B(n1077), .C(n1023), .D(n735), .Y(n117) );
  ao22d1_hd U1457 ( .A(n703), .B(n1079), .C(n1024), .D(n735), .Y(n118) );
  ao22d1_hd U1458 ( .A(n703), .B(n1081), .C(n1025), .D(n735), .Y(n119) );
  ao22d1_hd U1459 ( .A(n703), .B(n1083), .C(n1026), .D(n734), .Y(n120) );
  ao22d1_hd U1460 ( .A(n703), .B(n1085), .C(n1027), .D(n734), .Y(n121) );
  ao22d1_hd U1461 ( .A(n703), .B(n1087), .C(n1028), .D(n734), .Y(n122) );
  ao22d1_hd U1462 ( .A(n703), .B(n1089), .C(n1029), .D(n734), .Y(n123) );
  ao22d1_hd U1463 ( .A(n702), .B(n1091), .C(n1030), .D(n734), .Y(n124) );
  ao22d1_hd U1464 ( .A(n702), .B(n1093), .C(n1031), .D(n734), .Y(n125) );
  ao22d1_hd U1465 ( .A(n702), .B(n1095), .C(n1032), .D(n733), .Y(n126) );
  ao22d1_hd U1466 ( .A(n702), .B(n1097), .C(n1033), .D(n733), .Y(n127) );
  oa21d1_hd U1467 ( .A(n1035), .B(n702), .C(n1034), .Y(n128) );
  oa21d1_hd U1468 ( .A(n1037), .B(n702), .C(n1036), .Y(n129) );
  oa21d1_hd U1469 ( .A(n1039), .B(n701), .C(n1038), .Y(n130) );
  oa21d1_hd U1470 ( .A(n1041), .B(n701), .C(n1040), .Y(n131) );
  oa21d1_hd U1471 ( .A(n1043), .B(n701), .C(n1042), .Y(n132) );
  oa21d1_hd U1472 ( .A(n1045), .B(n701), .C(n1044), .Y(n133) );
  oa21d1_hd U1473 ( .A(n1047), .B(n701), .C(n1046), .Y(n134) );
  oa21d1_hd U1474 ( .A(n1049), .B(n701), .C(n1048), .Y(n135) );
  oa21d1_hd U1475 ( .A(n1051), .B(n700), .C(n1050), .Y(n136) );
  oa21d1_hd U1476 ( .A(n1053), .B(n700), .C(n1052), .Y(n137) );
  oa21d1_hd U1477 ( .A(n1055), .B(n700), .C(n1054), .Y(n138) );
  oa21d1_hd U1478 ( .A(n1057), .B(n700), .C(n1056), .Y(n139) );
  oa21d1_hd U1479 ( .A(n1059), .B(n700), .C(n1058), .Y(n140) );
  oa21d1_hd U1480 ( .A(n1061), .B(n700), .C(n1060), .Y(n141) );
  oa21d1_hd U1481 ( .A(n1063), .B(n699), .C(n1062), .Y(n142) );
  oa21d1_hd U1482 ( .A(n1065), .B(n699), .C(n1064), .Y(n143) );
  oa21d1_hd U1483 ( .A(n1067), .B(n699), .C(n1066), .Y(n144) );
  oa21d1_hd U1484 ( .A(n1069), .B(n699), .C(n1068), .Y(n145) );
  oa21d1_hd U1485 ( .A(n1071), .B(n699), .C(n1070), .Y(n146) );
  oa21d1_hd U1486 ( .A(n1073), .B(n699), .C(n1072), .Y(n147) );
  oa21d1_hd U1487 ( .A(n1075), .B(n698), .C(n1074), .Y(n148) );
  oa21d1_hd U1488 ( .A(n1077), .B(n698), .C(n1076), .Y(n149) );
  oa21d1_hd U1489 ( .A(n1079), .B(n698), .C(n1078), .Y(n150) );
  oa21d1_hd U1490 ( .A(n1081), .B(n698), .C(n1080), .Y(n151) );
  oa21d1_hd U1491 ( .A(n1083), .B(n698), .C(n1082), .Y(n152) );
  oa21d1_hd U1492 ( .A(n1085), .B(n698), .C(n1084), .Y(n153) );
  oa21d1_hd U1493 ( .A(n1087), .B(n697), .C(n1086), .Y(n154) );
  oa21d1_hd U1494 ( .A(n1089), .B(n697), .C(n1088), .Y(n155) );
  oa21d1_hd U1495 ( .A(n1091), .B(n697), .C(n1090), .Y(n156) );
  oa21d1_hd U1496 ( .A(n1093), .B(n697), .C(n1092), .Y(n157) );
  oa21d1_hd U1497 ( .A(n1095), .B(n697), .C(n1094), .Y(n158) );
  oa21d1_hd U1498 ( .A(n1097), .B(n697), .C(n1096), .Y(n159) );
endmodule

