
module float_adder_1 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3, C91_DATA2_4,
         C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8, n1, n2, n27, n265,
         n266, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n509, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23,
         C2_Z_22, C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16,
         C2_Z_15, C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_43J2_124_6938_n58, DP_OP_43J2_124_6938_n57,
         DP_OP_43J2_124_6938_n56, DP_OP_43J2_124_6938_n55,
         DP_OP_43J2_124_6938_n54, DP_OP_43J2_124_6938_n53,
         DP_OP_43J2_124_6938_n52, DP_OP_43J2_124_6938_n51,
         DP_OP_43J2_124_6938_n50, DP_OP_43J2_124_6938_n49,
         DP_OP_43J2_124_6938_n48, DP_OP_43J2_124_6938_n47,
         DP_OP_43J2_124_6938_n46, DP_OP_43J2_124_6938_n45,
         DP_OP_43J2_124_6938_n44, DP_OP_43J2_124_6938_n43,
         DP_OP_43J2_124_6938_n42, DP_OP_43J2_124_6938_n41,
         DP_OP_43J2_124_6938_n40, DP_OP_43J2_124_6938_n39,
         DP_OP_43J2_124_6938_n38, DP_OP_43J2_124_6938_n37,
         DP_OP_43J2_124_6938_n36, DP_OP_43J2_124_6938_n35,
         DP_OP_43J2_124_6938_n34, DP_OP_43J2_124_6938_n33,
         DP_OP_43J2_124_6938_n32, DP_OP_43J2_124_6938_n27,
         DP_OP_43J2_124_6938_n26, DP_OP_43J2_124_6938_n25,
         DP_OP_43J2_124_6938_n24, DP_OP_43J2_124_6938_n23,
         DP_OP_43J2_124_6938_n22, DP_OP_43J2_124_6938_n21,
         DP_OP_43J2_124_6938_n20, DP_OP_43J2_124_6938_n19,
         DP_OP_43J2_124_6938_n18, DP_OP_43J2_124_6938_n17,
         DP_OP_43J2_124_6938_n16, DP_OP_43J2_124_6938_n15,
         DP_OP_43J2_124_6938_n14, DP_OP_43J2_124_6938_n13,
         DP_OP_43J2_124_6938_n12, DP_OP_43J2_124_6938_n11,
         DP_OP_43J2_124_6938_n10, DP_OP_43J2_124_6938_n9,
         DP_OP_43J2_124_6938_n8, DP_OP_43J2_124_6938_n7,
         DP_OP_43J2_124_6938_n6, DP_OP_43J2_124_6938_n5,
         DP_OP_43J2_124_6938_n4, DP_OP_43J2_124_6938_n3,
         DP_OP_43J2_124_6938_n2, DP_OP_43J2_124_6938_n1,
         DP_OP_154J2_137_6175_n9, DP_OP_154J2_137_6175_n8,
         DP_OP_154J2_137_6175_n7, DP_OP_154J2_137_6175_n6,
         DP_OP_154J2_137_6175_n5, DP_OP_154J2_137_6175_n4,
         DP_OP_154J2_137_6175_n3, DP_OP_154J2_137_6175_n2, n1283, n1313, n1895,
         n1896, n1897, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J2_137_6175_U10 ( .A(n1896), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J2_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J2_137_6175_U9 ( .A(n1896), .B(z_e[2]), .CI(
        DP_OP_154J2_137_6175_n9), .CO(DP_OP_154J2_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J2_137_6175_U8 ( .A(n1896), .B(z_e[3]), .CI(
        DP_OP_154J2_137_6175_n8), .CO(DP_OP_154J2_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J2_137_6175_U7 ( .A(n1896), .B(z_e[4]), .CI(
        DP_OP_154J2_137_6175_n7), .CO(DP_OP_154J2_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J2_137_6175_U6 ( .A(n1896), .B(z_e[5]), .CI(
        DP_OP_154J2_137_6175_n6), .CO(DP_OP_154J2_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J2_137_6175_U5 ( .A(n1896), .B(z_e[6]), .CI(
        DP_OP_154J2_137_6175_n5), .CO(DP_OP_154J2_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J2_137_6175_U4 ( .A(n1896), .B(z_e[7]), .CI(
        DP_OP_154J2_137_6175_n4), .CO(DP_OP_154J2_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J2_137_6175_U3 ( .A(n1896), .B(z_e[8]), .CI(
        DP_OP_154J2_137_6175_n3), .CO(DP_OP_154J2_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1580), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n509), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n509), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1580), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1580), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1580), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1580), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1580), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n1580), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n1580), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n1580), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n1580), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n1580), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n1580), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n1580), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n1580), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1580), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1580), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1580), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1580), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1580), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n509), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n509), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n509), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n509), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1580), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1580), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n1580), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1580), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1580), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1580), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n1570), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n1570), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n1570), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n1570), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n1569), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n1569), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n1570), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n1570), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n1570), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n1570), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n1570), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n1570), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n1570), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n1570), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n1570), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n1570), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n1570), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n1570), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n1570), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n1570), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n1570), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n1570), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n1570), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n1570), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n1570), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n1570), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n1570), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n1570), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n1570), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n1570), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n1570), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n1570), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n1570), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n1570), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n1570), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n1570), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n1570), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n1570), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n1570), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n1570), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n1570), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n1570), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n1570), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n1570), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n1570), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n1570), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n1570), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n1570), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n1570), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n1570), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n1570), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n1570), .CK(i_CLK), .Q(b[22]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n1569), .CK(i_CLK), .Q(sum[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n1569), .CK(i_CLK), .Q(sum[2]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n1569), .CK(i_CLK), .Q(sum[26]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n1569), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n1569), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n1569), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n1569), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n1569), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n1569), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n1569), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n1569), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n1569), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n1569), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n1569), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n1569), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n1569), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n1569), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n1569), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n1569), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n1569), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n1569), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n1569), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n1569), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n1569), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n1569), .CK(i_CLK), .Q(sum[25]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n1569), .CK(i_CLK), .Q(sum[1]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n1570), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n1570), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n1570), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n1570), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n1569), .CK(i_CLK), .Q(sum[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n1570), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n1570), .CK(i_CLK), .Q(b[28]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n1570), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n1570), .CK(i_CLK), .Q(b[25]) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n1570), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n1570), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n1570), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n1570), .CK(i_CLK), .Q(b[26]) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n1570), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n1570), .CK(i_CLK), .Q(b[23]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n265), .CK(i_CLK), .Q(guard) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1577), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1577), .CK(i_CLK), .Q(a_s) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n1895), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n1895), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J2_124_6938_U28 ( .A(C2_Z_0), .B(n1313), .CI(
        DP_OP_43J2_124_6938_n58), .CO(DP_OP_43J2_124_6938_n27), .S(N310) );
  fad1_hd DP_OP_43J2_124_6938_U27 ( .A(DP_OP_43J2_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J2_124_6938_n27), .CO(DP_OP_43J2_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J2_124_6938_U26 ( .A(DP_OP_43J2_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J2_124_6938_n26), .CO(DP_OP_43J2_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J2_124_6938_U25 ( .A(DP_OP_43J2_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J2_124_6938_n25), .CO(DP_OP_43J2_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J2_124_6938_U24 ( .A(DP_OP_43J2_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J2_124_6938_n24), .CO(DP_OP_43J2_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J2_124_6938_U23 ( .A(DP_OP_43J2_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J2_124_6938_n23), .CO(DP_OP_43J2_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J2_124_6938_U2 ( .A(DP_OP_43J2_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J2_124_6938_n2), .CO(DP_OP_43J2_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J2_124_6938_U3 ( .A(DP_OP_43J2_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J2_124_6938_n3), .CO(DP_OP_43J2_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J2_124_6938_U4 ( .A(DP_OP_43J2_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J2_124_6938_n4), .CO(DP_OP_43J2_124_6938_n3), .S(N334) );
  fad1_hd DP_OP_43J2_124_6938_U5 ( .A(DP_OP_43J2_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J2_124_6938_n5), .CO(DP_OP_43J2_124_6938_n4), .S(N333) );
  fad1_hd DP_OP_43J2_124_6938_U6 ( .A(DP_OP_43J2_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J2_124_6938_n6), .CO(DP_OP_43J2_124_6938_n5), .S(N332) );
  fad1_hd DP_OP_43J2_124_6938_U7 ( .A(DP_OP_43J2_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J2_124_6938_n7), .CO(DP_OP_43J2_124_6938_n6), .S(N331) );
  fad1_hd DP_OP_43J2_124_6938_U8 ( .A(DP_OP_43J2_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J2_124_6938_n8), .CO(DP_OP_43J2_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J2_124_6938_U9 ( .A(DP_OP_43J2_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J2_124_6938_n9), .CO(DP_OP_43J2_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J2_124_6938_U10 ( .A(DP_OP_43J2_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J2_124_6938_n10), .CO(DP_OP_43J2_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J2_124_6938_U11 ( .A(DP_OP_43J2_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J2_124_6938_n11), .CO(DP_OP_43J2_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J2_124_6938_U12 ( .A(DP_OP_43J2_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J2_124_6938_n12), .CO(DP_OP_43J2_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J2_124_6938_U13 ( .A(DP_OP_43J2_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J2_124_6938_n13), .CO(DP_OP_43J2_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J2_124_6938_U14 ( .A(DP_OP_43J2_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J2_124_6938_n14), .CO(DP_OP_43J2_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J2_124_6938_U15 ( .A(DP_OP_43J2_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J2_124_6938_n15), .CO(DP_OP_43J2_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J2_124_6938_U16 ( .A(DP_OP_43J2_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J2_124_6938_n16), .CO(DP_OP_43J2_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J2_124_6938_U17 ( .A(DP_OP_43J2_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J2_124_6938_n17), .CO(DP_OP_43J2_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J2_124_6938_U18 ( .A(DP_OP_43J2_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J2_124_6938_n18), .CO(DP_OP_43J2_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J2_124_6938_U19 ( .A(DP_OP_43J2_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J2_124_6938_n19), .CO(DP_OP_43J2_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J2_124_6938_U20 ( .A(DP_OP_43J2_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J2_124_6938_n20), .CO(DP_OP_43J2_124_6938_n19), .S(N318)
         );
  fad1_hd DP_OP_43J2_124_6938_U21 ( .A(DP_OP_43J2_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J2_124_6938_n21), .CO(DP_OP_43J2_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J2_124_6938_U22 ( .A(DP_OP_43J2_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J2_124_6938_n22), .CO(DP_OP_43J2_124_6938_n21), .S(N316)
         );
  fd1qd1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK) );
  nr2d1_hd U523 ( .A(n1991), .B(n1935), .Y(n1952) );
  clknd2d1_hd U524 ( .A(b_m[5]), .B(n2084), .Y(n1587) );
  clknd2d1_hd U525 ( .A(n1595), .B(n1594), .Y(n1596) );
  clknd2d1_hd U526 ( .A(b_m[18]), .B(n1611), .Y(n1612) );
  clknd2d1_hd U527 ( .A(b_m[8]), .B(n2078), .Y(n1592) );
  clknd2d1_hd U528 ( .A(n1590), .B(b_m[7]), .Y(n1591) );
  clknd2d1_hd U529 ( .A(b_m[12]), .B(n2070), .Y(n1600) );
  clknd2d1_hd U530 ( .A(b_m[11]), .B(n1598), .Y(n1599) );
  clknd2d1_hd U531 ( .A(b_m[17]), .B(n2060), .Y(n1610) );
  clknd2d1_hd U532 ( .A(b_e[8]), .B(n2102), .Y(n1697) );
  clknd2d1_hd U533 ( .A(n1680), .B(n1679), .Y(n1688) );
  clknd2d1_hd U534 ( .A(b_e[6]), .B(n2100), .Y(n1679) );
  clknd2d1_hd U535 ( .A(a_e[9]), .B(n1683), .Y(n1700) );
  clknd2d1_hd U536 ( .A(b_m[19]), .B(n2056), .Y(n1613) );
  clknd2d1_hd U537 ( .A(n1700), .B(n1699), .Y(n1701) );
  clknd2d1_hd U538 ( .A(a_e[8]), .B(n2169), .Y(n1694) );
  clknd2d1_hd U539 ( .A(n2189), .B(n1701), .Y(n2235) );
  clknd2d1_hd U540 ( .A(n1705), .B(n1727), .Y(n2231) );
  clknd2d1_hd U541 ( .A(n1712), .B(n2097), .Y(n1715) );
  clknd2d1_hd U542 ( .A(n1703), .B(z_e[1]), .Y(n1727) );
  clknd2d1_hd U543 ( .A(n1717), .B(n1715), .Y(n1719) );
  clknd2d1_hd U544 ( .A(n1750), .B(n1792), .Y(n1716) );
  clknd2d1_hd U545 ( .A(n2163), .B(n1711), .Y(n1717) );
  clknd2d1_hd U546 ( .A(a_e[4]), .B(n2121), .Y(n2099) );
  clknd2d1_hd U547 ( .A(state[0]), .B(n2243), .Y(n2228) );
  clknd2d1_hd U548 ( .A(n1974), .B(guard), .Y(n1966) );
  clknd2d1_hd U549 ( .A(n1575), .B(n2189), .Y(n2252) );
  clknd2d1_hd U550 ( .A(n1718), .B(n2263), .Y(n1707) );
  clknd2d1_hd U551 ( .A(n1573), .B(n2189), .Y(n2094) );
  clknd2d1_hd U552 ( .A(n2188), .B(n2166), .Y(n2173) );
  clknd2d1_hd U553 ( .A(n2249), .B(n2243), .Y(n2246) );
  clknd2d1_hd U554 ( .A(n2205), .B(n2215), .Y(n2213) );
  clknd2d1_hd U555 ( .A(b_e[2]), .B(n2204), .Y(n2198) );
  clknd2d1_hd U556 ( .A(a_e[2]), .B(n2136), .Y(n2130) );
  clknd2d1_hd U557 ( .A(n2139), .B(n2131), .Y(n2129) );
  clknd2d1_hd U558 ( .A(n2139), .B(n2148), .Y(n2146) );
  clknd2d1_hd U559 ( .A(n2120), .B(n2098), .Y(n2106) );
  clknd2d1_hd U560 ( .A(n2180), .B(n2176), .Y(n2256) );
  clknd2d1_hd U561 ( .A(b_e[5]), .B(n2183), .Y(n2182) );
  clknd2d1_hd U562 ( .A(n2194), .B(b_e[4]), .Y(n2165) );
  clknd2d1_hd U563 ( .A(n2190), .B(b[28]), .Y(n2184) );
  clknd2d1_hd U564 ( .A(state[2]), .B(n2263), .Y(n2247) );
  clknd2d1_hd U565 ( .A(N41), .B(n2262), .Y(n2264) );
  clknd2d1_hd U566 ( .A(n1958), .B(n1949), .Y(n1940) );
  clknd2d1_hd U567 ( .A(n1945), .B(n1940), .Y(n1936) );
  clknd2d1_hd U568 ( .A(n1958), .B(n1921), .Y(n1928) );
  clknd2d1_hd U569 ( .A(z_m[21]), .B(n1967), .Y(n1960) );
  clknd2d1_hd U570 ( .A(n1975), .B(sum[27]), .Y(n1972) );
  clknd2d1_hd U571 ( .A(n1958), .B(n1893), .Y(n1903) );
  clknd2d1_hd U572 ( .A(n1958), .B(n1869), .Y(n1876) );
  clknd2d1_hd U573 ( .A(n1958), .B(n1970), .Y(n1827) );
  clknd2d1_hd U574 ( .A(n1958), .B(n1845), .Y(n1852) );
  clknd2d1_hd U575 ( .A(z_m[20]), .B(n1823), .Y(n1961) );
  clknd2d1_hd U576 ( .A(z_m[19]), .B(z_m[20]), .Y(n1813) );
  clknd2d1_hd U577 ( .A(n2193), .B(n2124), .Y(n1758) );
  clknd2d1_hd U578 ( .A(n2167), .B(n2100), .Y(n1743) );
  clknd2d1_hd U579 ( .A(b_e[0]), .B(a_e[0]), .Y(n1786) );
  clknd2d1_hd U580 ( .A(n1751), .B(n1750), .Y(n1779) );
  clknd2d1_hd U581 ( .A(n1778), .B(n1773), .Y(n1772) );
  clknd2d1_hd U582 ( .A(n1764), .B(n1760), .Y(n1759) );
  clknd2d1_hd U583 ( .A(b_e[7]), .B(a_e[7]), .Y(n1738) );
  clknd2d1_hd U584 ( .A(n1749), .B(n1745), .Y(n1744) );
  clknd2d1_hd U585 ( .A(n1796), .B(n1735), .Y(n1790) );
  clknd2d1_hd U586 ( .A(n1726), .B(n1725), .Y(n1729) );
  clknd2d1_hd U587 ( .A(state[1]), .B(n2249), .Y(n2225) );
  clknd2d1_hd U588 ( .A(state[3]), .B(n1718), .Y(n2224) );
  clknd2d1_hd U589 ( .A(a[23]), .B(a[24]), .Y(n2150) );
  clknd2d1_hd U590 ( .A(n2137), .B(a[26]), .Y(n2133) );
  clknd2d1_hd U591 ( .A(b[23]), .B(b[24]), .Y(n2217) );
  clknd2d1_hd U592 ( .A(n2216), .B(n2213), .Y(n2209) );
  clknd2d1_hd U593 ( .A(a_e[5]), .B(n2115), .Y(n2114) );
  clknd2d1_hd U594 ( .A(n2122), .B(a[28]), .Y(n2116) );
  clknd2d1_hd U595 ( .A(b_e[4]), .B(n2205), .Y(n2197) );
  clknd2d1_hd U596 ( .A(n2206), .B(b[26]), .Y(n2201) );
  clknd2d1_hd U597 ( .A(n1579), .B(n2170), .Y(n2175) );
  clknd2d1_hd U598 ( .A(n2203), .B(n2202), .Y(n495) );
  clknd2d1_hd U599 ( .A(a[30]), .B(n2103), .Y(n2108) );
  clknd2d1_hd U600 ( .A(n2184), .B(n2177), .Y(n2179) );
  clknd2d1_hd U601 ( .A(n1959), .B(n1940), .Y(n1942) );
  clknd2d1_hd U602 ( .A(n1996), .B(n1995), .Y(n428) );
  clknd2d1_hd U603 ( .A(DP_OP_154J2_137_6175_n2), .B(n1994), .Y(n1992) );
  clknd2d1_hd U604 ( .A(n1973), .B(n1805), .Y(n265) );
  clknd2d1_hd U605 ( .A(n1808), .B(n1807), .Y(n393) );
  clknd2d1_hd U606 ( .A(n1789), .B(n1741), .Y(n362) );
  clknd2d1_hd U607 ( .A(n2139), .B(n2136), .Y(n2145) );
  clknd2d1_hd U608 ( .A(n2139), .B(n2121), .Y(n2128) );
  clknd2d1_hd U609 ( .A(n2205), .B(n2204), .Y(n2212) );
  clknd2d1_hd U610 ( .A(n2116), .B(n2109), .Y(n2110) );
  ivd4_hd U611 ( .A(n1656), .Y(n1568) );
  ivd3_hd U612 ( .A(n1283), .Y(n1569) );
  oa22d2_hd U613 ( .A(n1657), .B(n1709), .C(a_s), .D(b_s), .Y(n1791) );
  xo2d1_hd U614 ( .A(n1313), .B(DP_OP_43J2_124_6938_n1), .Y(N337) );
  ad2d4_hd U615 ( .A(n1313), .B(n1626), .Y(n1656) );
  oa21d1_hd U616 ( .A(n1623), .B(n1622), .C(n1621), .Y(n1624) );
  ao21d1_hd U617 ( .A(a_m[23]), .B(n2000), .C(n1620), .Y(n1623) );
  nid1_hd U618 ( .A(n1802), .Y(n1571) );
  nid6_hd U619 ( .A(n27), .Y(n1570) );
  ad3d1_hd U620 ( .A(n2223), .B(i_AB_STB), .C(o_AB_ACK), .Y(n27) );
  ivd2_hd U621 ( .A(n1791), .Y(n1313) );
  or2d2_hd U622 ( .A(n1707), .B(n2228), .Y(n1897) );
  ivd1_hd U623 ( .A(b_m[23]), .Y(n2000) );
  nr2d4_hd U624 ( .A(n1656), .B(n1791), .Y(n1654) );
  scg9d1_hd U625 ( .A(n2241), .B(n1701), .C(n1897), .Y(n2161) );
  scg2d1_hd U626 ( .A(b_e[9]), .B(n1698), .C(n1697), .D(n1696), .Y(n1699) );
  ad3d1_hd U627 ( .A(n2261), .B(n1576), .C(n2259), .Y(n2265) );
  ivd2_hd U628 ( .A(n1779), .Y(n1804) );
  ivd2_hd U629 ( .A(n1972), .Y(n1946) );
  or4d1_hd U630 ( .A(z_m[23]), .B(z_e[0]), .C(n1728), .D(n1727), .Y(n1735) );
  or4d1_hd U631 ( .A(n1678), .B(a_e[9]), .C(a_e[0]), .D(a_e[8]), .Y(n1792) );
  or2d1_hd U632 ( .A(n2246), .B(n2247), .Y(n1283) );
  ivd1_hd U633 ( .A(b_m[1]), .Y(n2043) );
  ivd1_hd U634 ( .A(b_m[2]), .Y(n2042) );
  or2d1_hd U635 ( .A(b_e[2]), .B(a_e[2]), .Y(n1771) );
  nr2d2_hd U636 ( .A(n1797), .B(n2227), .Y(n1803) );
  ivd2_hd U637 ( .A(n1952), .Y(n1959) );
  nr2ad1_hd U638 ( .A(n1976), .B(n1989), .Y(n1993) );
  nr2ad1_hd U639 ( .A(n2259), .B(n1935), .Y(n1941) );
  nr2ad1_hd U640 ( .A(n2225), .B(n2247), .Y(n1896) );
  ivd1_hd U641 ( .A(b_m[0]), .Y(n2044) );
  oa22ad1_hd U642 ( .A(n1589), .B(a_m[6]), .C(n1588), .D(b_m[6]), .Y(n1590) );
  ivd1_hd U643 ( .A(b_m[3]), .Y(n2041) );
  ivd1_hd U644 ( .A(b_m[4]), .Y(n2038) );
  ao22d1_hd U645 ( .A(a_m[26]), .B(n2253), .C(n1625), .D(n1624), .Y(n1626) );
  ivd1_hd U646 ( .A(a_m[3]), .Y(n2089) );
  ivd1_hd U647 ( .A(a_m[5]), .Y(n2084) );
  ivd1_hd U648 ( .A(b_m[5]), .Y(n2036) );
  nid2_hd U649 ( .A(n2260), .Y(n1576) );
  ivd1_hd U650 ( .A(n1958), .Y(n1934) );
  ivd1_hd U651 ( .A(n1987), .Y(n1989) );
  ivd1_hd U652 ( .A(n2096), .Y(n1574) );
  oa21d1_hd U653 ( .A(a_m[21]), .B(n2004), .C(n1617), .Y(n1618) );
  ivd1_hd U654 ( .A(a_m[4]), .Y(n2086) );
  ivd1_hd U655 ( .A(n1787), .Y(n1800) );
  ivd1_hd U656 ( .A(n1897), .Y(n1577) );
  nr2d1_hd U657 ( .A(n2261), .B(n1935), .Y(n1958) );
  ivd1_hd U658 ( .A(n1974), .Y(n2261) );
  nid2_hd U659 ( .A(n1947), .Y(n1572) );
  ivd1_hd U660 ( .A(n1941), .Y(n1948) );
  nr2d1_hd U661 ( .A(n2224), .B(n2246), .Y(n1974) );
  ivd1_hd U662 ( .A(n1896), .Y(n1991) );
  ivd2_hd U663 ( .A(n2161), .Y(n1575) );
  ivd2_hd U664 ( .A(n1574), .Y(n1573) );
  ivd1_hd U665 ( .A(n1895), .Y(n2226) );
  ivd1_hd U666 ( .A(n2241), .Y(n2189) );
  nd2bd1_hd U667 ( .AN(n1707), .B(n2237), .Y(n2241) );
  ivd1_hd U668 ( .A(b_m[24]), .Y(n1998) );
  ivd1_hd U669 ( .A(a_m[16]), .Y(n2062) );
  ivd1_hd U670 ( .A(b_m[10]), .Y(n2026) );
  ivd1_hd U671 ( .A(b_m[13]), .Y(n2020) );
  ivd1_hd U672 ( .A(a_m[15]), .Y(n2064) );
  ivd1_hd U673 ( .A(b_m[14]), .Y(n2018) );
  ivd1_hd U674 ( .A(a_m[17]), .Y(n2060) );
  ivd1_hd U675 ( .A(b_m[17]), .Y(n2012) );
  ivd1_hd U676 ( .A(b_m[21]), .Y(n2004) );
  nid2_hd U677 ( .A(n509), .Y(n1580) );
  nr3d1_hd U678 ( .A(n1751), .B(n1717), .C(n1716), .Y(n1802) );
  ivd1_hd U679 ( .A(n1715), .Y(n1751) );
  ivd2_hd U680 ( .A(n2252), .Y(n2039) );
  scg20d2_hd U681 ( .A(n1812), .B(n1966), .C(n265), .Y(n1935) );
  ivd1_hd U682 ( .A(n1975), .Y(n1805) );
  ivd2_hd U683 ( .A(n1897), .Y(n1578) );
  ivd2_hd U684 ( .A(n2094), .Y(n2087) );
  nr2d1_hd U685 ( .A(n2228), .B(n2247), .Y(n1975) );
  nd2bd1_hd U686 ( .AN(n2247), .B(n2237), .Y(n2259) );
  ivd1_hd U687 ( .A(n2205), .Y(n2255) );
  nr2d1_hd U688 ( .A(n2221), .B(n2241), .Y(n2205) );
  ao21d1_hd U689 ( .A(n2163), .B(n2162), .C(n1575), .Y(n2221) );
  ivd1_hd U690 ( .A(n1897), .Y(n1579) );
  ivd1_hd U691 ( .A(n2139), .Y(n2157) );
  nr2d1_hd U692 ( .A(n2154), .B(n2241), .Y(n2139) );
  ao21d1_hd U693 ( .A(n2097), .B(n2162), .C(n1573), .Y(n2154) );
  scg16d1_hd U694 ( .A(n2236), .B(n2235), .C(n1897), .Y(n2096) );
  ivd1_hd U695 ( .A(b_e[1]), .Y(n2215) );
  nr2d1_hd U696 ( .A(n1719), .B(n1716), .Y(n2162) );
  nr2d1_hd U697 ( .A(n1707), .B(n2225), .Y(n1895) );
  ivd1_hd U698 ( .A(b_e[6]), .Y(n2167) );
  ivd1_hd U699 ( .A(a_e[8]), .Y(n2102) );
  ivd1_hd U700 ( .A(a_e[5]), .Y(n2119) );
  ivd1_hd U701 ( .A(a_e[6]), .Y(n2100) );
  nr2d1_hd U702 ( .A(n2249), .B(n2243), .Y(n2237) );
  ivd1_hd U703 ( .A(state[0]), .Y(n2249) );
  ivd1_hd U704 ( .A(state[1]), .Y(n2243) );
  ivd1_hd U705 ( .A(state[3]), .Y(n2263) );
  ivd1_hd U706 ( .A(b_m[25]), .Y(n1628) );
  ivd1_hd U707 ( .A(b_m[19]), .Y(n2008) );
  ivd1_hd U708 ( .A(b_m[20]), .Y(n2006) );
  ivd1_hd U709 ( .A(a_m[20]), .Y(n2054) );
  ivd1_hd U710 ( .A(b_m[22]), .Y(n2002) );
  ivd1_hd U711 ( .A(a_m[22]), .Y(n2050) );
  ivd1_hd U712 ( .A(a_m[25]), .Y(n1668) );
  ivd1_hd U713 ( .A(b_m[26]), .Y(n2253) );
  ivd1_hd U714 ( .A(n2162), .Y(n2245) );
  nr2d1_hd U715 ( .A(n2225), .B(n2224), .Y(n509) );
  ivd1_hd U716 ( .A(n1796), .Y(n2227) );
  ivd1_hd U717 ( .A(z_m[1]), .Y(n1949) );
  ao21d1_hd U718 ( .A(n1796), .B(n1797), .C(n1734), .Y(n1789) );
  ivd1_hd U719 ( .A(n1710), .Y(n1793) );
  nr2d1_hd U720 ( .A(n2228), .B(n2224), .Y(n1796) );
  ivd1_hd U721 ( .A(z_m[20]), .Y(n1832) );
  ivd1_hd U722 ( .A(z_m[21]), .Y(n1826) );
  ivd1_hd U723 ( .A(n1935), .Y(n1955) );
  ivd1_hd U724 ( .A(z_m[22]), .Y(n1968) );
  ivd1_hd U725 ( .A(z_m[17]), .Y(n1850) );
  ivd1_hd U726 ( .A(z_m[18]), .Y(n1838) );
  ivd1_hd U727 ( .A(z_m[13]), .Y(n1874) );
  ivd1_hd U728 ( .A(z_m[14]), .Y(n1862) );
  ivd1_hd U729 ( .A(z_m[10]), .Y(n1886) );
  ivd1_hd U730 ( .A(z_m[9]), .Y(n1901) );
  ivd1_hd U731 ( .A(z_m[5]), .Y(n1926) );
  ivd1_hd U732 ( .A(z_m[6]), .Y(n1913) );
  ivd1_hd U733 ( .A(z_m[23]), .Y(n1967) );
  ivd1_hd U734 ( .A(z_e[0]), .Y(n1988) );
  ivd1_hd U735 ( .A(z_e[7]), .Y(n1733) );
  ivd1_hd U736 ( .A(z_e[8]), .Y(n1978) );
  ivd1_hd U737 ( .A(n2257), .Y(n2210) );
  nr2d1_hd U738 ( .A(n2226), .B(n2221), .Y(n2257) );
  ivd1_hd U739 ( .A(b[30]), .Y(n2176) );
  ivd1_hd U740 ( .A(n2159), .Y(n2143) );
  nr2d1_hd U741 ( .A(n2226), .B(n2154), .Y(n2159) );
  ivd1_hd U742 ( .A(a_e[7]), .Y(n2104) );
  ivd1_hd U743 ( .A(a_e[4]), .Y(n2124) );
  ivd1_hd U744 ( .A(a_e[2]), .Y(n2140) );
  ivd1_hd U745 ( .A(b_e[7]), .Y(n2171) );
  nr3d1_hd U746 ( .A(n1676), .B(n1675), .C(n1674), .Y(n1712) );
  ivd1_hd U747 ( .A(b_e[9]), .Y(n1683) );
  ivd1_hd U748 ( .A(b_e[0]), .Y(n2214) );
  ivd1_hd U749 ( .A(b_e[5]), .Y(n2187) );
  ivd1_hd U750 ( .A(b_e[8]), .Y(n2169) );
  ivd1_hd U751 ( .A(a_e[0]), .Y(n2147) );
  ivd1_hd U752 ( .A(a_e[1]), .Y(n2148) );
  ivd1_hd U753 ( .A(a_e[3]), .Y(n2131) );
  ivd1_hd U754 ( .A(state[2]), .Y(n1718) );
  ivd1_hd U755 ( .A(a_m[1]), .Y(n2091) );
  ivd1_hd U756 ( .A(a_m[2]), .Y(n2090) );
  ivd1_hd U757 ( .A(a_m[6]), .Y(n2082) );
  ivd1_hd U758 ( .A(b_m[6]), .Y(n2034) );
  ivd1_hd U759 ( .A(a_m[7]), .Y(n2080) );
  ivd1_hd U760 ( .A(b_m[7]), .Y(n2032) );
  ivd1_hd U761 ( .A(a_m[11]), .Y(n2072) );
  ivd1_hd U762 ( .A(b_m[11]), .Y(n2024) );
  ivd1_hd U763 ( .A(a_m[13]), .Y(n2068) );
  ivd1_hd U764 ( .A(a_m[14]), .Y(n2066) );
  ivd1_hd U765 ( .A(a_m[18]), .Y(n2058) );
  ivd1_hd U766 ( .A(b_m[18]), .Y(n2010) );
  ivd1_hd U767 ( .A(a_m[21]), .Y(n2052) );
  ivd1_hd U768 ( .A(a_m[23]), .Y(n2048) );
  ivd1_hd U769 ( .A(a_m[24]), .Y(n2046) );
  ivd1_hd U770 ( .A(a_m[19]), .Y(n2056) );
  ivd1_hd U771 ( .A(b_m[15]), .Y(n2016) );
  ivd1_hd U772 ( .A(b_m[16]), .Y(n2014) );
  ivd1_hd U773 ( .A(a_m[12]), .Y(n2070) );
  ivd1_hd U774 ( .A(a_m[8]), .Y(n2078) );
  ivd1_hd U775 ( .A(b_m[8]), .Y(n2030) );
  ivd1_hd U776 ( .A(b_m[9]), .Y(n2028) );
  ivd1_hd U777 ( .A(a_m[10]), .Y(n2074) );
  ivd1_hd U778 ( .A(a_m[9]), .Y(n2076) );
  ivd1_hd U779 ( .A(b_m[12]), .Y(n2022) );
  ivd1_hd U780 ( .A(a_m[26]), .Y(n2095) );
  ivd1_hd U781 ( .A(a_s), .Y(n1709) );
  ivd1_hd U782 ( .A(b_s), .Y(n1657) );
  ivd1_hd U783 ( .A(z_m[0]), .Y(n1956) );
  nr2d1_hd U784 ( .A(n1576), .B(n2226), .Y(n1787) );
  nd2bd1_hd U785 ( .AN(a[30]), .B(n2111), .Y(n2158) );
  ivd1_hd U786 ( .A(a_e[9]), .Y(n1698) );
  nr2d1_hd U787 ( .A(sum[27]), .B(n1805), .Y(n1947) );
  ao22d1_hd U788 ( .A(b_m[25]), .B(n1668), .C(b_m[26]), .D(n2095), .Y(n1625)
         );
  ao22d1_hd U789 ( .A(a_m[21]), .B(n2004), .C(a_m[22]), .D(n2002), .Y(n1619)
         );
  ao22d1_hd U790 ( .A(a_m[20]), .B(n2006), .C(a_m[19]), .D(n2008), .Y(n1616)
         );
  nr2d1_hd U791 ( .A(b_m[15]), .B(n2064), .Y(n1606) );
  ao22d1_hd U792 ( .A(a_m[13]), .B(n2020), .C(a_m[12]), .D(n2022), .Y(n1604)
         );
  ao22d1_hd U793 ( .A(b_m[9]), .B(n2076), .C(b_m[10]), .D(n2074), .Y(n1597) );
  ao22d1_hd U794 ( .A(a_m[9]), .B(n2028), .C(a_m[8]), .D(n2030), .Y(n1595) );
  ao211d1_hd U795 ( .A(a_m[1]), .B(n2043), .C(a_m[0]), .D(n2044), .Y(n1582) );
  oa22d1_hd U796 ( .A(a_m[1]), .B(n2043), .C(a_m[2]), .D(n2042), .Y(n1581) );
  oa22d1_hd U797 ( .A(b_m[3]), .B(n2089), .C(n1582), .D(n1581), .Y(n1583) );
  ao21d1_hd U798 ( .A(a_m[2]), .B(n2042), .C(n1583), .Y(n1585) );
  oa22d1_hd U799 ( .A(a_m[4]), .B(n2038), .C(a_m[3]), .D(n2041), .Y(n1584) );
  oa22d1_hd U800 ( .A(n1585), .B(n1584), .C(b_m[4]), .D(n2086), .Y(n1586) );
  ao22d1_hd U801 ( .A(a_m[5]), .B(n2036), .C(n1587), .D(n1586), .Y(n1588) );
  nr2d1_hd U802 ( .A(n1588), .B(b_m[6]), .Y(n1589) );
  nr2d1_hd U803 ( .A(n1590), .B(b_m[7]), .Y(n1593) );
  oa211d1_hd U804 ( .A(a_m[7]), .B(n1593), .C(n1592), .D(n1591), .Y(n1594) );
  ao22d1_hd U805 ( .A(a_m[10]), .B(n2026), .C(n1597), .D(n1596), .Y(n1598) );
  nr2d1_hd U806 ( .A(b_m[11]), .B(n1598), .Y(n1601) );
  oa211d1_hd U807 ( .A(a_m[11]), .B(n1601), .C(n1600), .D(n1599), .Y(n1603) );
  oa22d1_hd U808 ( .A(a_m[13]), .B(n2020), .C(a_m[14]), .D(n2018), .Y(n1602)
         );
  ao21d1_hd U809 ( .A(n1604), .B(n1603), .C(n1602), .Y(n1605) );
  ao211d1_hd U810 ( .A(a_m[14]), .B(n2018), .C(n1606), .D(n1605), .Y(n1608) );
  oa22d1_hd U811 ( .A(a_m[16]), .B(n2014), .C(a_m[15]), .D(n2016), .Y(n1607)
         );
  oa22d1_hd U812 ( .A(n1608), .B(n1607), .C(b_m[16]), .D(n2062), .Y(n1609) );
  ao22d1_hd U813 ( .A(a_m[17]), .B(n2012), .C(n1610), .D(n1609), .Y(n1611) );
  nr2d1_hd U814 ( .A(b_m[18]), .B(n1611), .Y(n1614) );
  oa211d1_hd U815 ( .A(a_m[18]), .B(n1614), .C(n1613), .D(n1612), .Y(n1615) );
  ao22d1_hd U816 ( .A(b_m[20]), .B(n2054), .C(n1616), .D(n1615), .Y(n1617) );
  ao22d1_hd U817 ( .A(b_m[22]), .B(n2050), .C(n1619), .D(n1618), .Y(n1620) );
  oa22d1_hd U818 ( .A(a_m[23]), .B(n2000), .C(a_m[24]), .D(n1998), .Y(n1622)
         );
  ao22d1_hd U819 ( .A(a_m[24]), .B(n1998), .C(a_m[25]), .D(n1628), .Y(n1621)
         );
  ivd1_hd U820 ( .A(a_m[0]), .Y(n2092) );
  ao22d1_hd U821 ( .A(n1656), .B(n2044), .C(n2092), .D(n1568), .Y(C2_Z_0) );
  ao22d1_hd U822 ( .A(n1656), .B(n2043), .C(n2091), .D(n1568), .Y(C2_Z_1) );
  ao22d1_hd U823 ( .A(n1656), .B(n2026), .C(n2074), .D(n1568), .Y(C2_Z_10) );
  ao22d1_hd U824 ( .A(n1656), .B(n2024), .C(n2072), .D(n1568), .Y(C2_Z_11) );
  ao22d1_hd U825 ( .A(n1656), .B(n2022), .C(n2070), .D(n1568), .Y(C2_Z_12) );
  ao22d1_hd U826 ( .A(n1656), .B(n2020), .C(n2068), .D(n1568), .Y(C2_Z_13) );
  ao22d1_hd U827 ( .A(n1656), .B(n2018), .C(n2066), .D(n1568), .Y(C2_Z_14) );
  ao22d1_hd U828 ( .A(n1656), .B(n2016), .C(n2064), .D(n1568), .Y(C2_Z_15) );
  ao22d1_hd U829 ( .A(n1656), .B(n2014), .C(n2062), .D(n1568), .Y(C2_Z_16) );
  ao22d1_hd U830 ( .A(n1656), .B(n2012), .C(n2060), .D(n1568), .Y(C2_Z_17) );
  ao22d1_hd U831 ( .A(n1656), .B(n2010), .C(n2058), .D(n1568), .Y(C2_Z_18) );
  ao22d1_hd U832 ( .A(n1656), .B(n2008), .C(n2056), .D(n1568), .Y(C2_Z_19) );
  ao22d1_hd U833 ( .A(n1656), .B(n2042), .C(n2090), .D(n1568), .Y(C2_Z_2) );
  ao22d1_hd U834 ( .A(n1656), .B(n2006), .C(n2054), .D(n1568), .Y(C2_Z_20) );
  ao22d1_hd U835 ( .A(n1656), .B(n2004), .C(n2052), .D(n1568), .Y(C2_Z_21) );
  ao22d1_hd U836 ( .A(n1656), .B(n2002), .C(n2050), .D(n1568), .Y(C2_Z_22) );
  ao22d1_hd U837 ( .A(n1656), .B(n2000), .C(n2048), .D(n1568), .Y(C2_Z_23) );
  ao22d1_hd U838 ( .A(n1656), .B(n1998), .C(n2046), .D(n1568), .Y(C2_Z_24) );
  ao22d1_hd U839 ( .A(n1656), .B(n1628), .C(n1668), .D(n1568), .Y(C2_Z_25) );
  oa21d1_hd U840 ( .A(n2253), .B(n1791), .C(n2095), .Y(C2_Z_26) );
  ao22d1_hd U841 ( .A(n1656), .B(n2041), .C(n2089), .D(n1568), .Y(C2_Z_3) );
  ao22d1_hd U842 ( .A(n1656), .B(n2038), .C(n2086), .D(n1568), .Y(C2_Z_4) );
  ao22d1_hd U843 ( .A(n1656), .B(n2036), .C(n2084), .D(n1568), .Y(C2_Z_5) );
  ao22d1_hd U844 ( .A(n1656), .B(n2034), .C(n2082), .D(n1568), .Y(C2_Z_6) );
  ao22d1_hd U845 ( .A(n1656), .B(n2032), .C(n2080), .D(n1568), .Y(C2_Z_7) );
  ao22d1_hd U846 ( .A(n1656), .B(n2030), .C(n2078), .D(n1568), .Y(C2_Z_8) );
  ao22d1_hd U847 ( .A(n1656), .B(n2028), .C(n2076), .D(n1568), .Y(C2_Z_9) );
  nr2d1_hd U848 ( .A(n2253), .B(n2095), .Y(n1627) );
  ao22d1_hd U849 ( .A(n1313), .B(n1627), .C(n2253), .D(n1791), .Y(
        DP_OP_43J2_124_6938_n32) );
  ao22d1_hd U850 ( .A(b_m[25]), .B(n1791), .C(n1654), .D(n1628), .Y(n1629) );
  oa21d1_hd U851 ( .A(a_m[25]), .B(n1568), .C(n1629), .Y(
        DP_OP_43J2_124_6938_n33) );
  ao22d1_hd U852 ( .A(b_m[24]), .B(n1791), .C(n1654), .D(n1998), .Y(n1630) );
  oa21d1_hd U853 ( .A(a_m[24]), .B(n1568), .C(n1630), .Y(
        DP_OP_43J2_124_6938_n34) );
  ao22d1_hd U854 ( .A(b_m[23]), .B(n1791), .C(n1654), .D(n2000), .Y(n1631) );
  oa21d1_hd U855 ( .A(a_m[23]), .B(n1568), .C(n1631), .Y(
        DP_OP_43J2_124_6938_n35) );
  ao22d1_hd U856 ( .A(n1656), .B(n2050), .C(n1654), .D(n2002), .Y(n1632) );
  oa21d1_hd U857 ( .A(n1313), .B(n2002), .C(n1632), .Y(DP_OP_43J2_124_6938_n36) );
  ao22d1_hd U858 ( .A(b_m[21]), .B(n1791), .C(n1654), .D(n2004), .Y(n1633) );
  oa21d1_hd U859 ( .A(a_m[21]), .B(n1568), .C(n1633), .Y(
        DP_OP_43J2_124_6938_n37) );
  ao22d1_hd U860 ( .A(n1656), .B(n2054), .C(n1654), .D(n2006), .Y(n1634) );
  oa21d1_hd U861 ( .A(n1313), .B(n2006), .C(n1634), .Y(DP_OP_43J2_124_6938_n38) );
  ao22d1_hd U862 ( .A(n1656), .B(n2056), .C(n1654), .D(n2008), .Y(n1635) );
  oa21d1_hd U863 ( .A(n1313), .B(n2008), .C(n1635), .Y(DP_OP_43J2_124_6938_n39) );
  ao22d1_hd U864 ( .A(b_m[18]), .B(n1791), .C(n1654), .D(n2010), .Y(n1636) );
  oa21d1_hd U865 ( .A(a_m[18]), .B(n1568), .C(n1636), .Y(
        DP_OP_43J2_124_6938_n40) );
  ao22d1_hd U866 ( .A(n1656), .B(n2060), .C(n1654), .D(n2012), .Y(n1637) );
  oa21d1_hd U867 ( .A(n1313), .B(n2012), .C(n1637), .Y(DP_OP_43J2_124_6938_n41) );
  ao22d1_hd U868 ( .A(n1656), .B(n2062), .C(n1654), .D(n2014), .Y(n1638) );
  oa21d1_hd U869 ( .A(n1313), .B(n2014), .C(n1638), .Y(DP_OP_43J2_124_6938_n42) );
  ao22d1_hd U870 ( .A(n1656), .B(n2064), .C(n1654), .D(n2016), .Y(n1639) );
  oa21d1_hd U871 ( .A(n1313), .B(n2016), .C(n1639), .Y(DP_OP_43J2_124_6938_n43) );
  ao22d1_hd U872 ( .A(b_m[14]), .B(n1791), .C(n1654), .D(n2018), .Y(n1640) );
  oa21d1_hd U873 ( .A(a_m[14]), .B(n1568), .C(n1640), .Y(
        DP_OP_43J2_124_6938_n44) );
  ao22d1_hd U874 ( .A(b_m[13]), .B(n1791), .C(n1654), .D(n2020), .Y(n1641) );
  oa21d1_hd U875 ( .A(a_m[13]), .B(n1568), .C(n1641), .Y(
        DP_OP_43J2_124_6938_n45) );
  ao22d1_hd U876 ( .A(n1656), .B(n2070), .C(n1654), .D(n2022), .Y(n1642) );
  oa21d1_hd U877 ( .A(n1313), .B(n2022), .C(n1642), .Y(DP_OP_43J2_124_6938_n46) );
  ao22d1_hd U878 ( .A(b_m[11]), .B(n1791), .C(n1654), .D(n2024), .Y(n1643) );
  oa21d1_hd U879 ( .A(a_m[11]), .B(n1568), .C(n1643), .Y(
        DP_OP_43J2_124_6938_n47) );
  ao22d1_hd U880 ( .A(n1656), .B(n2074), .C(n1654), .D(n2026), .Y(n1644) );
  oa21d1_hd U881 ( .A(n1313), .B(n2026), .C(n1644), .Y(DP_OP_43J2_124_6938_n48) );
  ao22d1_hd U882 ( .A(n1656), .B(n2076), .C(n1654), .D(n2028), .Y(n1645) );
  oa21d1_hd U883 ( .A(n1313), .B(n2028), .C(n1645), .Y(DP_OP_43J2_124_6938_n49) );
  ao22d1_hd U884 ( .A(n1656), .B(n2078), .C(n1654), .D(n2030), .Y(n1646) );
  oa21d1_hd U885 ( .A(n1313), .B(n2030), .C(n1646), .Y(DP_OP_43J2_124_6938_n50) );
  ao22d1_hd U886 ( .A(b_m[7]), .B(n1791), .C(n1654), .D(n2032), .Y(n1647) );
  oa21d1_hd U887 ( .A(a_m[7]), .B(n1568), .C(n1647), .Y(
        DP_OP_43J2_124_6938_n51) );
  ao22d1_hd U888 ( .A(b_m[6]), .B(n1791), .C(n1654), .D(n2034), .Y(n1648) );
  oa21d1_hd U889 ( .A(a_m[6]), .B(n1568), .C(n1648), .Y(
        DP_OP_43J2_124_6938_n52) );
  ao22d1_hd U890 ( .A(n1656), .B(n2084), .C(n1654), .D(n2036), .Y(n1649) );
  oa21d1_hd U891 ( .A(n1313), .B(n2036), .C(n1649), .Y(DP_OP_43J2_124_6938_n53) );
  ao22d1_hd U892 ( .A(n1656), .B(n2086), .C(n1654), .D(n2038), .Y(n1650) );
  oa21d1_hd U893 ( .A(n1313), .B(n2038), .C(n1650), .Y(DP_OP_43J2_124_6938_n54) );
  ao22d1_hd U894 ( .A(n1656), .B(n2089), .C(n1654), .D(n2041), .Y(n1651) );
  oa21d1_hd U895 ( .A(n1313), .B(n2041), .C(n1651), .Y(DP_OP_43J2_124_6938_n55) );
  ao22d1_hd U896 ( .A(b_m[2]), .B(n1791), .C(n1654), .D(n2042), .Y(n1652) );
  oa21d1_hd U897 ( .A(a_m[2]), .B(n1568), .C(n1652), .Y(
        DP_OP_43J2_124_6938_n56) );
  ao22d1_hd U898 ( .A(b_m[1]), .B(n1791), .C(n1654), .D(n2043), .Y(n1653) );
  oa21d1_hd U899 ( .A(a_m[1]), .B(n1568), .C(n1653), .Y(
        DP_OP_43J2_124_6938_n57) );
  ao22d1_hd U900 ( .A(b_m[0]), .B(n1791), .C(n1654), .D(n2044), .Y(n1655) );
  oa21d1_hd U901 ( .A(a_m[0]), .B(n1568), .C(n1655), .Y(
        DP_OP_43J2_124_6938_n58) );
  ao22d1_hd U902 ( .A(n1656), .B(n1657), .C(n1709), .D(n1568), .Y(N338) );
  nr4d1_hd U903 ( .A(a_e[1]), .B(a_e[2]), .C(a_e[3]), .D(a_e[4]), .Y(n1658) );
  nd4d1_hd U904 ( .A(a_e[7]), .B(n1658), .C(n2100), .D(n2119), .Y(n1678) );
  nr4d1_hd U905 ( .A(n1678), .B(n2147), .C(n1698), .D(n2102), .Y(n2097) );
  nr4d1_hd U906 ( .A(b_e[2]), .B(b_e[1]), .C(b_e[3]), .D(b_e[4]), .Y(n1659) );
  nd4d1_hd U907 ( .A(b_e[7]), .B(n1659), .C(n2187), .D(n2167), .Y(n1677) );
  nr4d1_hd U908 ( .A(n2169), .B(n1677), .C(n2214), .D(n1683), .Y(n2163) );
  nd4d1_hd U909 ( .A(n2036), .B(n2038), .C(n2028), .D(n2016), .Y(n1667) );
  nr4d1_hd U910 ( .A(b_m[0]), .B(b_m[1]), .C(b_m[2]), .D(b_m[3]), .Y(n1660) );
  nd4d1_hd U911 ( .A(n1660), .B(n2014), .C(n2034), .D(n2020), .Y(n1666) );
  nr4d1_hd U912 ( .A(b_m[25]), .B(b_m[23]), .C(b_m[22]), .D(b_m[26]), .Y(n1664) );
  nr4d1_hd U913 ( .A(b_m[18]), .B(b_m[11]), .C(b_m[14]), .D(b_m[24]), .Y(n1663) );
  nr4d1_hd U914 ( .A(b_m[8]), .B(b_m[7]), .C(b_m[10]), .D(b_m[12]), .Y(n1662)
         );
  nr4d1_hd U915 ( .A(b_m[17]), .B(b_m[19]), .C(b_m[20]), .D(b_m[21]), .Y(n1661) );
  nd4d1_hd U916 ( .A(n1664), .B(n1663), .C(n1662), .D(n1661), .Y(n1665) );
  nr3d1_hd U917 ( .A(n1667), .B(n1666), .C(n1665), .Y(n1711) );
  nd4d1_hd U918 ( .A(n2060), .B(n2078), .C(n2052), .D(n2046), .Y(n1676) );
  nr4d1_hd U919 ( .A(a_m[18]), .B(a_m[12]), .C(a_m[20]), .D(a_m[26]), .Y(n1669) );
  nd4d1_hd U920 ( .A(n1669), .B(n2048), .C(n2050), .D(n1668), .Y(n1675) );
  nr4d1_hd U921 ( .A(a_m[11]), .B(a_m[6]), .C(a_m[9]), .D(a_m[10]), .Y(n1673)
         );
  nr4d1_hd U922 ( .A(a_m[13]), .B(a_m[14]), .C(a_m[15]), .D(a_m[19]), .Y(n1672) );
  nr4d1_hd U923 ( .A(a_m[16]), .B(a_m[5]), .C(a_m[4]), .D(a_m[7]), .Y(n1671)
         );
  nr4d1_hd U924 ( .A(a_m[0]), .B(a_m[1]), .C(a_m[2]), .D(a_m[3]), .Y(n1670) );
  nd4d1_hd U925 ( .A(n1673), .B(n1672), .C(n1671), .D(n1670), .Y(n1674) );
  nr4d1_hd U926 ( .A(b_e[8]), .B(b_e[0]), .C(b_e[9]), .D(n1677), .Y(n1710) );
  nr2d1_hd U927 ( .A(n1710), .B(n2226), .Y(n1750) );
  ao22d1_hd U928 ( .A(b_e[2]), .B(n2140), .C(b_e[3]), .D(n2131), .Y(n1685) );
  nr2d1_hd U929 ( .A(a_e[1]), .B(n2215), .Y(n1681) );
  ao22d1_hd U930 ( .A(b_e[4]), .B(n2124), .C(b_e[5]), .D(n2119), .Y(n1680) );
  ao211d1_hd U931 ( .A(b_e[0]), .B(n2147), .C(n1681), .D(n1688), .Y(n1682) );
  oa211d1_hd U932 ( .A(a_e[7]), .B(n2171), .C(n1685), .D(n1682), .Y(n1684) );
  nd3bd1_hd U933 ( .AN(n1684), .B(n1697), .C(n1700), .Y(n2236) );
  ao211d1_hd U934 ( .A(b_e[6]), .B(n2100), .C(b_e[5]), .D(n2119), .Y(n1692) );
  ivd1_hd U935 ( .A(b_e[4]), .Y(n2193) );
  ivd1_hd U936 ( .A(b_e[3]), .Y(n2164) );
  ao22d1_hd U937 ( .A(a_e[4]), .B(n2193), .C(a_e[3]), .D(n2164), .Y(n1690) );
  ao211d1_hd U938 ( .A(b_e[1]), .B(n2148), .C(b_e[0]), .D(n2147), .Y(n1687) );
  oa22d1_hd U939 ( .A(b_e[1]), .B(n2148), .C(b_e[2]), .D(n2140), .Y(n1686) );
  oa21d1_hd U940 ( .A(n1687), .B(n1686), .C(n1685), .Y(n1689) );
  ao21d1_hd U941 ( .A(n1690), .B(n1689), .C(n1688), .Y(n1691) );
  ao211d1_hd U942 ( .A(a_e[6]), .B(n2167), .C(n1692), .D(n1691), .Y(n1695) );
  scg6d1_hd U943 ( .A(b_e[7]), .B(n1695), .C(n2104), .Y(n1693) );
  oa211d1_hd U944 ( .A(b_e[7]), .B(n1695), .C(n1694), .D(n1693), .Y(n1696) );
  oa21d1_hd U945 ( .A(n2097), .B(n2245), .C(n1574), .Y(n1) );
  oa21d1_hd U946 ( .A(n2163), .B(n2245), .C(n2161), .Y(n2) );
  nr2d1_hd U947 ( .A(n1733), .B(n1978), .Y(n1703) );
  nr4d1_hd U948 ( .A(z_e[2]), .B(z_e[3]), .C(z_e[4]), .D(z_e[5]), .Y(n1702) );
  ivd1_hd U949 ( .A(z_e[6]), .Y(n1745) );
  nd3d1_hd U950 ( .A(z_e[9]), .B(n1702), .C(n1745), .Y(n1728) );
  ivd1_hd U951 ( .A(z_e[9]), .Y(n1990) );
  ao21d1_hd U952 ( .A(n1703), .B(n1728), .C(n1990), .Y(n1705) );
  nr2d1_hd U953 ( .A(n2259), .B(n2231), .Y(n1806) );
  nr2d1_hd U954 ( .A(n1727), .B(n1988), .Y(n1704) );
  scg16d1_hd U955 ( .A(n1705), .B(n1704), .C(n1967), .Y(n2230) );
  nr2d1_hd U956 ( .A(n2230), .B(n1991), .Y(n1706) );
  nr2d1_hd U957 ( .A(n1806), .B(n1706), .Y(n1973) );
  ivd1_hd U958 ( .A(n2259), .Y(n2232) );
  scg4d1_hd U959 ( .A(n2232), .B(z_m[0]), .C(n1896), .D(round_bit), .E(n1572), 
        .F(sum[2]), .G(sum[3]), .H(n1946), .Y(n266) );
  nr2d1_hd U960 ( .A(n1707), .B(n2246), .Y(n2223) );
  nr2d1_hd U961 ( .A(a_s), .B(n1717), .Y(n1708) );
  oa21d1_hd U962 ( .A(n1715), .B(n1708), .C(n1793), .Y(n1714) );
  nr3d1_hd U963 ( .A(n1710), .B(n1792), .C(n1709), .Y(n1713) );
  oa22d1_hd U964 ( .A(n1712), .B(n1792), .C(n1711), .D(n1793), .Y(n1794) );
  ao211d1_hd U965 ( .A(b_s), .B(n1714), .C(n1713), .D(n1794), .Y(n1732) );
  ao21d1_hd U966 ( .A(n1792), .B(n1793), .C(n2226), .Y(n1734) );
  ao211d1_hd U967 ( .A(n1895), .B(n1719), .C(n1734), .D(n1796), .Y(n2260) );
  ao22d1_hd U968 ( .A(a_s), .B(n1571), .C(n1576), .D(z[31]), .Y(n1731) );
  ivd1_hd U969 ( .A(z_m[4]), .Y(n1919) );
  ivd1_hd U970 ( .A(z_m[3]), .Y(n1927) );
  nd4d1_hd U971 ( .A(n1949), .B(n1919), .C(n1927), .D(n1913), .Y(n1720) );
  nr4d1_hd U972 ( .A(z_m[0]), .B(z_m[19]), .C(z_m[2]), .D(n1720), .Y(n1726) );
  ivd1_hd U973 ( .A(z_m[12]), .Y(n1868) );
  ivd1_hd U974 ( .A(z_m[11]), .Y(n1875) );
  nd4d1_hd U975 ( .A(n1886), .B(n1868), .C(n1875), .D(n1862), .Y(n1724) );
  ivd1_hd U976 ( .A(z_m[8]), .Y(n1892) );
  ivd1_hd U977 ( .A(z_m[7]), .Y(n1902) );
  nd4d1_hd U978 ( .A(n1926), .B(n1892), .C(n1902), .D(n1901), .Y(n1723) );
  nd4d1_hd U979 ( .A(n1968), .B(n1826), .C(n1832), .D(n1850), .Y(n1722) );
  ivd1_hd U980 ( .A(z_m[16]), .Y(n1844) );
  ivd1_hd U981 ( .A(z_m[15]), .Y(n1851) );
  nd4d1_hd U982 ( .A(n1874), .B(n1844), .C(n1851), .D(n1838), .Y(n1721) );
  nr4d1_hd U983 ( .A(n1724), .B(n1723), .C(n1722), .D(n1721), .Y(n1725) );
  oa211d1_hd U984 ( .A(n1729), .B(n1735), .C(n1796), .D(z_s), .Y(n1730) );
  oa211d1_hd U985 ( .A(n1732), .B(n2226), .C(n1731), .D(n1730), .Y(n361) );
  ao21d1_hd U986 ( .A(n1733), .B(n1978), .C(z_e[9]), .Y(n1797) );
  nr2d1_hd U987 ( .A(z_e[1]), .B(z_e[0]), .Y(n1778) );
  ivd1_hd U988 ( .A(z_e[2]), .Y(n1773) );
  nr2d1_hd U989 ( .A(z_e[3]), .B(n1772), .Y(n1764) );
  ivd1_hd U990 ( .A(z_e[4]), .Y(n1760) );
  nr2d1_hd U991 ( .A(z_e[5]), .B(n1759), .Y(n1749) );
  nr2d1_hd U992 ( .A(z_e[7]), .B(n1744), .Y(n1736) );
  ao211d1_hd U993 ( .A(z_e[7]), .B(n1744), .C(n1790), .D(n1736), .Y(n1740) );
  nd3d1_hd U994 ( .A(n2215), .B(n2148), .C(n1786), .Y(n1780) );
  nr2d1_hd U995 ( .A(n1780), .B(n1771), .Y(n1770) );
  nd3d1_hd U996 ( .A(n1770), .B(n2164), .C(n2131), .Y(n1765) );
  nr2d1_hd U997 ( .A(n1765), .B(n1758), .Y(n1757) );
  nd3d1_hd U998 ( .A(n1757), .B(n2187), .C(n2119), .Y(n1752) );
  nr2d1_hd U999 ( .A(n1752), .B(n1743), .Y(n1742) );
  nr2d1_hd U1000 ( .A(n1742), .B(n1738), .Y(n1737) );
  ao211d1_hd U1001 ( .A(n1742), .B(n1738), .C(n1800), .D(n1737), .Y(n1739) );
  ao211d1_hd U1002 ( .A(n1576), .B(z[30]), .C(n1740), .D(n1739), .Y(n1741) );
  ao21d1_hd U1003 ( .A(n1752), .B(n1743), .C(n1742), .Y(n1748) );
  ivd1_hd U1004 ( .A(n1790), .Y(n1775) );
  oa21d1_hd U1005 ( .A(n1749), .B(n1745), .C(n1744), .Y(n1746) );
  ao22d1_hd U1006 ( .A(n1576), .B(z[29]), .C(n1775), .D(n1746), .Y(n1747) );
  oa211d1_hd U1007 ( .A(n1748), .B(n1800), .C(n1789), .D(n1747), .Y(n363) );
  ao21d1_hd U1008 ( .A(z_e[5]), .B(n1759), .C(n1749), .Y(n1756) );
  ao22d1_hd U1009 ( .A(b_e[5]), .B(n1804), .C(a_e[5]), .D(n1787), .Y(n1753) );
  oa22d1_hd U1010 ( .A(n1757), .B(n1753), .C(n1800), .D(n1752), .Y(n1754) );
  ao21d1_hd U1011 ( .A(n1576), .B(z[28]), .C(n1754), .Y(n1755) );
  oa211d1_hd U1012 ( .A(n1756), .B(n1790), .C(n1789), .D(n1755), .Y(n364) );
  ao21d1_hd U1013 ( .A(n1765), .B(n1758), .C(n1757), .Y(n1763) );
  oa21d1_hd U1014 ( .A(n1764), .B(n1760), .C(n1759), .Y(n1761) );
  ao22d1_hd U1015 ( .A(n1576), .B(z[27]), .C(n1775), .D(n1761), .Y(n1762) );
  oa211d1_hd U1016 ( .A(n1763), .B(n1800), .C(n1789), .D(n1762), .Y(n365) );
  ao21d1_hd U1017 ( .A(z_e[3]), .B(n1772), .C(n1764), .Y(n1769) );
  ao22d1_hd U1018 ( .A(b_e[3]), .B(n1804), .C(a_e[3]), .D(n1787), .Y(n1766) );
  oa22d1_hd U1019 ( .A(n1770), .B(n1766), .C(n1800), .D(n1765), .Y(n1767) );
  ao21d1_hd U1020 ( .A(n1576), .B(z[26]), .C(n1767), .Y(n1768) );
  oa211d1_hd U1021 ( .A(n1769), .B(n1790), .C(n1789), .D(n1768), .Y(n366) );
  ao21d1_hd U1022 ( .A(n1780), .B(n1771), .C(n1770), .Y(n1777) );
  oa21d1_hd U1023 ( .A(n1778), .B(n1773), .C(n1772), .Y(n1774) );
  ao22d1_hd U1024 ( .A(n1576), .B(z[25]), .C(n1775), .D(n1774), .Y(n1776) );
  oa211d1_hd U1025 ( .A(n1777), .B(n1800), .C(n1789), .D(n1776), .Y(n367) );
  ao21d1_hd U1026 ( .A(z_e[0]), .B(z_e[1]), .C(n1778), .Y(n1785) );
  nr3d1_hd U1027 ( .A(n2215), .B(n1786), .C(n1779), .Y(n1783) );
  nd2bd1_hd U1028 ( .AN(n1786), .B(a_e[1]), .Y(n1781) );
  ao21d1_hd U1029 ( .A(n1781), .B(n1780), .C(n1800), .Y(n1782) );
  ao211d1_hd U1030 ( .A(n1576), .B(z[24]), .C(n1783), .D(n1782), .Y(n1784) );
  oa211d1_hd U1031 ( .A(n1785), .B(n1790), .C(n1789), .D(n1784), .Y(n368) );
  ao22d1_hd U1032 ( .A(n1576), .B(z[23]), .C(n1787), .D(n1786), .Y(n1788) );
  oa211d1_hd U1033 ( .A(z_e[0]), .B(n1790), .C(n1789), .D(n1788), .Y(n369) );
  nr3d1_hd U1034 ( .A(n1793), .B(n1792), .C(n1791), .Y(n1795) );
  nr2d1_hd U1035 ( .A(n1795), .B(n1794), .Y(n1801) );
  ao22d1_hd U1036 ( .A(b_m[25]), .B(n1804), .C(z_m[22]), .D(n1803), .Y(n1799)
         );
  ao22d1_hd U1037 ( .A(a_m[25]), .B(n1571), .C(n1576), .D(z[22]), .Y(n1798) );
  oa211d1_hd U1038 ( .A(n1801), .B(n1800), .C(n1799), .D(n1798), .Y(n370) );
  scg4d1_hd U1039 ( .A(b_m[24]), .B(n1804), .C(z_m[21]), .D(n1803), .E(a_m[24]), .F(n1571), .G(n1576), .H(z[21]), .Y(n371) );
  scg4d1_hd U1040 ( .A(b_m[23]), .B(n1804), .C(z_m[20]), .D(n1803), .E(a_m[23]), .F(n1571), .G(n1576), .H(z[20]), .Y(n372) );
  scg4d1_hd U1041 ( .A(b_m[22]), .B(n1804), .C(z_m[19]), .D(n1803), .E(a_m[22]), .F(n1571), .G(n1576), .H(z[19]), .Y(n373) );
  scg4d1_hd U1042 ( .A(b_m[21]), .B(n1804), .C(z_m[18]), .D(n1803), .E(a_m[21]), .F(n1571), .G(n1576), .H(z[18]), .Y(n374) );
  scg4d1_hd U1043 ( .A(b_m[20]), .B(n1804), .C(z_m[17]), .D(n1803), .E(a_m[20]), .F(n1571), .G(n1576), .H(z[17]), .Y(n375) );
  scg4d1_hd U1044 ( .A(b_m[19]), .B(n1804), .C(z_m[16]), .D(n1803), .E(a_m[19]), .F(n1571), .G(n1576), .H(z[16]), .Y(n376) );
  scg4d1_hd U1045 ( .A(b_m[18]), .B(n1804), .C(z_m[15]), .D(n1803), .E(a_m[18]), .F(n1571), .G(n1576), .H(z[15]), .Y(n377) );
  scg4d1_hd U1046 ( .A(b_m[17]), .B(n1804), .C(z_m[14]), .D(n1803), .E(a_m[17]), .F(n1571), .G(n1576), .H(z[14]), .Y(n378) );
  scg4d1_hd U1047 ( .A(b_m[16]), .B(n1804), .C(z_m[13]), .D(n1803), .E(a_m[16]), .F(n1571), .G(n1576), .H(z[13]), .Y(n379) );
  scg4d1_hd U1048 ( .A(b_m[15]), .B(n1804), .C(z_m[12]), .D(n1803), .E(a_m[15]), .F(n1571), .G(n1576), .H(z[12]), .Y(n380) );
  scg4d1_hd U1049 ( .A(b_m[14]), .B(n1804), .C(z_m[11]), .D(n1803), .E(a_m[14]), .F(n1802), .G(n1576), .H(z[11]), .Y(n381) );
  scg4d1_hd U1050 ( .A(b_m[13]), .B(n1804), .C(z_m[10]), .D(n1803), .E(a_m[13]), .F(n1802), .G(n1576), .H(z[10]), .Y(n382) );
  scg4d1_hd U1051 ( .A(b_m[12]), .B(n1804), .C(z_m[9]), .D(n1803), .E(a_m[12]), 
        .F(n1802), .G(n1576), .H(z[9]), .Y(n383) );
  scg4d1_hd U1052 ( .A(b_m[11]), .B(n1804), .C(z_m[8]), .D(n1803), .E(a_m[11]), 
        .F(n1802), .G(n1576), .H(z[8]), .Y(n384) );
  scg4d1_hd U1053 ( .A(b_m[10]), .B(n1804), .C(z_m[7]), .D(n1803), .E(a_m[10]), 
        .F(n1802), .G(n1576), .H(z[7]), .Y(n385) );
  scg4d1_hd U1054 ( .A(b_m[9]), .B(n1804), .C(z_m[6]), .D(n1803), .E(a_m[9]), 
        .F(n1802), .G(n1576), .H(z[6]), .Y(n386) );
  scg4d1_hd U1055 ( .A(b_m[8]), .B(n1804), .C(z_m[5]), .D(n1803), .E(a_m[8]), 
        .F(n1571), .G(n1576), .H(z[5]), .Y(n387) );
  scg4d1_hd U1056 ( .A(b_m[7]), .B(n1804), .C(z_m[4]), .D(n1803), .E(a_m[7]), 
        .F(n1571), .G(n2260), .H(z[4]), .Y(n388) );
  scg4d1_hd U1057 ( .A(b_m[6]), .B(n1804), .C(z_m[3]), .D(n1803), .E(a_m[6]), 
        .F(n1571), .G(n1576), .H(z[3]), .Y(n389) );
  scg4d1_hd U1058 ( .A(b_m[5]), .B(n1804), .C(z_m[2]), .D(n1803), .E(a_m[5]), 
        .F(n1571), .G(n1576), .H(z[2]), .Y(n390) );
  scg4d1_hd U1059 ( .A(b_m[4]), .B(n1804), .C(z_m[1]), .D(n1803), .E(a_m[4]), 
        .F(n1571), .G(n1576), .H(z[1]), .Y(n391) );
  scg4d1_hd U1060 ( .A(b_m[3]), .B(n1804), .C(z_m[0]), .D(n1803), .E(a_m[3]), 
        .F(n1802), .G(n1576), .H(z[0]), .Y(n392) );
  ao22d1_hd U1061 ( .A(n1975), .B(sum[0]), .C(sticky), .D(n1805), .Y(n1808) );
  ao22d1_hd U1062 ( .A(n1806), .B(round_bit), .C(n1946), .D(sum[1]), .Y(n1807)
         );
  ivd1_hd U1063 ( .A(round_bit), .Y(n1811) );
  ao22d1_hd U1064 ( .A(n1572), .B(sum[1]), .C(n1946), .D(sum[2]), .Y(n1810) );
  nd3d1_hd U1065 ( .A(n2232), .B(guard), .C(n265), .Y(n1809) );
  oa211d1_hd U1066 ( .A(n1811), .B(n265), .C(n1810), .D(n1809), .Y(n394) );
  nr3d1_hd U1067 ( .A(z_m[0]), .B(sticky), .C(round_bit), .Y(n1812) );
  ao22d1_hd U1068 ( .A(n1572), .B(sum[25]), .C(n1946), .D(sum[26]), .Y(n1816)
         );
  nd3d1_hd U1069 ( .A(z_m[0]), .B(z_m[2]), .C(z_m[1]), .Y(n1920) );
  ivd1_hd U1070 ( .A(n1920), .Y(n1921) );
  nd3d1_hd U1071 ( .A(n1921), .B(z_m[4]), .C(z_m[3]), .Y(n1908) );
  nr3d1_hd U1072 ( .A(n1908), .B(n1913), .C(n1926), .Y(n1893) );
  nd3d1_hd U1073 ( .A(n1893), .B(z_m[8]), .C(z_m[7]), .Y(n1881) );
  nr3d1_hd U1074 ( .A(n1881), .B(n1901), .C(n1886), .Y(n1869) );
  nd3d1_hd U1075 ( .A(n1869), .B(z_m[12]), .C(z_m[11]), .Y(n1857) );
  nr3d1_hd U1076 ( .A(n1857), .B(n1862), .C(n1874), .Y(n1845) );
  nd3d1_hd U1077 ( .A(n1845), .B(z_m[16]), .C(z_m[15]), .Y(n1833) );
  nr3d1_hd U1078 ( .A(n1833), .B(n1838), .C(n1850), .Y(n1970) );
  oa21d1_hd U1079 ( .A(n1970), .B(n2261), .C(n1955), .Y(n1829) );
  ao21d1_hd U1080 ( .A(n1974), .B(n1813), .C(n1829), .Y(n1817) );
  oa21d1_hd U1081 ( .A(z_m[21]), .B(n1934), .C(n1817), .Y(n1957) );
  ivd1_hd U1082 ( .A(z_m[19]), .Y(n1965) );
  nr2d1_hd U1083 ( .A(n1965), .B(n1827), .Y(n1823) );
  oa21d1_hd U1084 ( .A(z_m[22]), .B(n1961), .C(n1959), .Y(n1814) );
  ao22d1_hd U1085 ( .A(z_m[22]), .B(n1957), .C(z_m[21]), .D(n1814), .Y(n1815)
         );
  oa211d1_hd U1086 ( .A(n1967), .B(n1948), .C(n1816), .D(n1815), .Y(n395) );
  ao22d1_hd U1087 ( .A(n1572), .B(sum[24]), .C(sum[25]), .D(n1946), .Y(n1820)
         );
  ao22d1_hd U1088 ( .A(z_m[21]), .B(n1817), .C(n1961), .D(n1826), .Y(n1818) );
  ao21d1_hd U1089 ( .A(z_m[20]), .B(n1952), .C(n1818), .Y(n1819) );
  oa211d1_hd U1090 ( .A(n1968), .B(n1948), .C(n1820), .D(n1819), .Y(n396) );
  ao22d1_hd U1091 ( .A(n1572), .B(sum[23]), .C(n1946), .D(sum[24]), .Y(n1825)
         );
  ao21d1_hd U1092 ( .A(n1958), .B(n1965), .C(n1829), .Y(n1821) );
  oa22d1_hd U1093 ( .A(n1821), .B(n1832), .C(n1965), .D(n1959), .Y(n1822) );
  ao21d1_hd U1094 ( .A(n1823), .B(n1832), .C(n1822), .Y(n1824) );
  oa211d1_hd U1095 ( .A(n1826), .B(n1948), .C(n1825), .D(n1824), .Y(n397) );
  ao22d1_hd U1096 ( .A(n1572), .B(sum[22]), .C(n1946), .D(sum[23]), .Y(n1831)
         );
  oa22d1_hd U1097 ( .A(z_m[19]), .B(n1827), .C(n1959), .D(n1838), .Y(n1828) );
  ao21d1_hd U1098 ( .A(z_m[19]), .B(n1829), .C(n1828), .Y(n1830) );
  oa211d1_hd U1099 ( .A(n1832), .B(n1948), .C(n1831), .D(n1830), .Y(n398) );
  nr2d1_hd U1100 ( .A(n1934), .B(n1833), .Y(n1841) );
  ao21d1_hd U1101 ( .A(n1841), .B(n1838), .C(n1952), .Y(n1837) );
  ao22d1_hd U1102 ( .A(n1572), .B(sum[21]), .C(n1946), .D(sum[22]), .Y(n1836)
         );
  ao21d1_hd U1103 ( .A(n1974), .B(n1833), .C(n1935), .Y(n1839) );
  oa21d1_hd U1104 ( .A(z_m[17]), .B(n1934), .C(n1839), .Y(n1834) );
  ao22d1_hd U1105 ( .A(z_m[19]), .B(n1941), .C(z_m[18]), .D(n1834), .Y(n1835)
         );
  oa211d1_hd U1106 ( .A(n1837), .B(n1850), .C(n1836), .D(n1835), .Y(n399) );
  ao22d1_hd U1107 ( .A(n1572), .B(sum[20]), .C(n1946), .D(sum[21]), .Y(n1843)
         );
  oa22d1_hd U1108 ( .A(n1839), .B(n1850), .C(n1838), .D(n1948), .Y(n1840) );
  ao21d1_hd U1109 ( .A(n1841), .B(n1850), .C(n1840), .Y(n1842) );
  oa211d1_hd U1110 ( .A(n1844), .B(n1959), .C(n1843), .D(n1842), .Y(n400) );
  ao22d1_hd U1111 ( .A(n1572), .B(sum[19]), .C(n1946), .D(sum[20]), .Y(n1849)
         );
  scg20d1_hd U1112 ( .A(n2261), .B(n1845), .C(n1935), .Y(n1853) );
  oa21d1_hd U1113 ( .A(z_m[15]), .B(n1934), .C(n1853), .Y(n1847) );
  oa21d1_hd U1114 ( .A(z_m[16]), .B(n1852), .C(n1959), .Y(n1846) );
  ao22d1_hd U1115 ( .A(z_m[16]), .B(n1847), .C(z_m[15]), .D(n1846), .Y(n1848)
         );
  oa211d1_hd U1116 ( .A(n1850), .B(n1948), .C(n1849), .D(n1848), .Y(n401) );
  ao22d1_hd U1117 ( .A(n1572), .B(sum[18]), .C(n1946), .D(sum[19]), .Y(n1856)
         );
  ao22d1_hd U1118 ( .A(z_m[15]), .B(n1853), .C(n1852), .D(n1851), .Y(n1854) );
  ao21d1_hd U1119 ( .A(z_m[16]), .B(n1941), .C(n1854), .Y(n1855) );
  oa211d1_hd U1120 ( .A(n1862), .B(n1959), .C(n1856), .D(n1855), .Y(n402) );
  nr2d1_hd U1121 ( .A(n1934), .B(n1857), .Y(n1865) );
  ao21d1_hd U1122 ( .A(n1865), .B(n1862), .C(n1952), .Y(n1861) );
  ao22d1_hd U1123 ( .A(n1572), .B(sum[17]), .C(n1946), .D(sum[18]), .Y(n1860)
         );
  ao21d1_hd U1124 ( .A(n1974), .B(n1857), .C(n1935), .Y(n1863) );
  oa21d1_hd U1125 ( .A(z_m[13]), .B(n1934), .C(n1863), .Y(n1858) );
  ao22d1_hd U1126 ( .A(z_m[14]), .B(n1858), .C(z_m[15]), .D(n1941), .Y(n1859)
         );
  oa211d1_hd U1127 ( .A(n1861), .B(n1874), .C(n1860), .D(n1859), .Y(n403) );
  ao22d1_hd U1128 ( .A(n1572), .B(sum[16]), .C(n1946), .D(sum[17]), .Y(n1867)
         );
  oa22d1_hd U1129 ( .A(n1863), .B(n1874), .C(n1862), .D(n1948), .Y(n1864) );
  ao21d1_hd U1130 ( .A(n1865), .B(n1874), .C(n1864), .Y(n1866) );
  oa211d1_hd U1131 ( .A(n1868), .B(n1959), .C(n1867), .D(n1866), .Y(n404) );
  ao22d1_hd U1132 ( .A(n1572), .B(sum[15]), .C(n1946), .D(sum[16]), .Y(n1873)
         );
  scg20d1_hd U1133 ( .A(n2261), .B(n1869), .C(n1935), .Y(n1877) );
  oa21d1_hd U1134 ( .A(z_m[11]), .B(n1934), .C(n1877), .Y(n1871) );
  oa21d1_hd U1135 ( .A(z_m[12]), .B(n1876), .C(n1959), .Y(n1870) );
  ao22d1_hd U1136 ( .A(z_m[12]), .B(n1871), .C(z_m[11]), .D(n1870), .Y(n1872)
         );
  oa211d1_hd U1137 ( .A(n1874), .B(n1948), .C(n1873), .D(n1872), .Y(n405) );
  ao22d1_hd U1138 ( .A(n1572), .B(sum[14]), .C(n1946), .D(sum[15]), .Y(n1880)
         );
  ao22d1_hd U1139 ( .A(z_m[11]), .B(n1877), .C(n1876), .D(n1875), .Y(n1878) );
  ao21d1_hd U1140 ( .A(z_m[12]), .B(n1941), .C(n1878), .Y(n1879) );
  oa211d1_hd U1141 ( .A(n1886), .B(n1959), .C(n1880), .D(n1879), .Y(n406) );
  nr2d1_hd U1142 ( .A(n1934), .B(n1881), .Y(n1889) );
  ao21d1_hd U1143 ( .A(n1889), .B(n1886), .C(n1952), .Y(n1885) );
  ao22d1_hd U1144 ( .A(n1572), .B(sum[13]), .C(n1946), .D(sum[14]), .Y(n1884)
         );
  ao21d1_hd U1145 ( .A(n1974), .B(n1881), .C(n1935), .Y(n1887) );
  oa21d1_hd U1146 ( .A(z_m[9]), .B(n1934), .C(n1887), .Y(n1882) );
  ao22d1_hd U1147 ( .A(z_m[10]), .B(n1882), .C(z_m[11]), .D(n1941), .Y(n1883)
         );
  oa211d1_hd U1148 ( .A(n1885), .B(n1901), .C(n1884), .D(n1883), .Y(n407) );
  ao22d1_hd U1149 ( .A(n1572), .B(sum[12]), .C(n1946), .D(sum[13]), .Y(n1891)
         );
  oa22d1_hd U1150 ( .A(n1887), .B(n1901), .C(n1886), .D(n1948), .Y(n1888) );
  ao21d1_hd U1151 ( .A(n1889), .B(n1901), .C(n1888), .Y(n1890) );
  oa211d1_hd U1152 ( .A(n1892), .B(n1959), .C(n1891), .D(n1890), .Y(n408) );
  ao22d1_hd U1153 ( .A(n1572), .B(sum[11]), .C(n1946), .D(sum[12]), .Y(n1900)
         );
  scg20d1_hd U1154 ( .A(n2261), .B(n1893), .C(n1935), .Y(n1904) );
  oa21d1_hd U1155 ( .A(z_m[7]), .B(n1934), .C(n1904), .Y(n1898) );
  oa21d1_hd U1156 ( .A(z_m[8]), .B(n1903), .C(n1959), .Y(n1894) );
  ao22d1_hd U1157 ( .A(z_m[8]), .B(n1898), .C(z_m[7]), .D(n1894), .Y(n1899) );
  oa211d1_hd U1158 ( .A(n1901), .B(n1948), .C(n1900), .D(n1899), .Y(n409) );
  ao22d1_hd U1159 ( .A(n1572), .B(sum[10]), .C(n1946), .D(sum[11]), .Y(n1907)
         );
  ao22d1_hd U1160 ( .A(z_m[7]), .B(n1904), .C(n1903), .D(n1902), .Y(n1905) );
  ao21d1_hd U1161 ( .A(z_m[8]), .B(n1941), .C(n1905), .Y(n1906) );
  oa211d1_hd U1162 ( .A(n1913), .B(n1959), .C(n1907), .D(n1906), .Y(n410) );
  nr2d1_hd U1163 ( .A(n1934), .B(n1908), .Y(n1916) );
  ao21d1_hd U1164 ( .A(n1916), .B(n1913), .C(n1952), .Y(n1912) );
  ao22d1_hd U1165 ( .A(n1572), .B(sum[9]), .C(n1946), .D(sum[10]), .Y(n1911)
         );
  ao21d1_hd U1166 ( .A(n1974), .B(n1908), .C(n1935), .Y(n1914) );
  oa21d1_hd U1167 ( .A(z_m[5]), .B(n1934), .C(n1914), .Y(n1909) );
  ao22d1_hd U1168 ( .A(z_m[6]), .B(n1909), .C(z_m[7]), .D(n1941), .Y(n1910) );
  oa211d1_hd U1169 ( .A(n1912), .B(n1926), .C(n1911), .D(n1910), .Y(n411) );
  ao22d1_hd U1170 ( .A(n1572), .B(sum[8]), .C(n1946), .D(sum[9]), .Y(n1918) );
  oa22d1_hd U1171 ( .A(n1914), .B(n1926), .C(n1913), .D(n1948), .Y(n1915) );
  ao21d1_hd U1172 ( .A(n1916), .B(n1926), .C(n1915), .Y(n1917) );
  oa211d1_hd U1173 ( .A(n1919), .B(n1959), .C(n1918), .D(n1917), .Y(n412) );
  ao22d1_hd U1174 ( .A(n1572), .B(sum[7]), .C(n1946), .D(sum[8]), .Y(n1925) );
  ao21d1_hd U1175 ( .A(n1974), .B(n1920), .C(n1935), .Y(n1929) );
  oa21d1_hd U1176 ( .A(z_m[3]), .B(n1934), .C(n1929), .Y(n1923) );
  oa21d1_hd U1177 ( .A(z_m[4]), .B(n1928), .C(n1959), .Y(n1922) );
  ao22d1_hd U1178 ( .A(z_m[4]), .B(n1923), .C(z_m[3]), .D(n1922), .Y(n1924) );
  oa211d1_hd U1179 ( .A(n1926), .B(n1948), .C(n1925), .D(n1924), .Y(n413) );
  ao22d1_hd U1180 ( .A(n1572), .B(sum[6]), .C(n1946), .D(sum[7]), .Y(n1932) );
  ao22d1_hd U1181 ( .A(z_m[3]), .B(n1929), .C(n1928), .D(n1927), .Y(n1930) );
  ao21d1_hd U1182 ( .A(z_m[4]), .B(n1941), .C(n1930), .Y(n1931) );
  scg15d1_hd U1183 ( .A(z_m[2]), .B(n1952), .C(n1932), .D(n1931), .Y(n414) );
  nr3d1_hd U1184 ( .A(z_m[2]), .B(n1934), .C(n1956), .Y(n1933) );
  nr2d1_hd U1185 ( .A(n1933), .B(n1952), .Y(n1939) );
  ao22d1_hd U1186 ( .A(n1572), .B(sum[5]), .C(n1946), .D(sum[6]), .Y(n1938) );
  nr2d1_hd U1187 ( .A(z_m[0]), .B(n1934), .Y(n1951) );
  nr2d1_hd U1188 ( .A(n1935), .B(n1951), .Y(n1945) );
  ao22d1_hd U1189 ( .A(z_m[2]), .B(n1936), .C(z_m[3]), .D(n1941), .Y(n1937) );
  oa211d1_hd U1190 ( .A(n1939), .B(n1949), .C(n1938), .D(n1937), .Y(n415) );
  ao22d1_hd U1191 ( .A(n1572), .B(sum[4]), .C(n1946), .D(sum[5]), .Y(n1944) );
  ao22d1_hd U1192 ( .A(z_m[0]), .B(n1942), .C(z_m[2]), .D(n1941), .Y(n1943) );
  oa211d1_hd U1193 ( .A(n1945), .B(n1949), .C(n1944), .D(n1943), .Y(n416) );
  ao22d1_hd U1194 ( .A(n1572), .B(sum[3]), .C(n1946), .D(sum[4]), .Y(n1954) );
  nr2d1_hd U1195 ( .A(n1949), .B(n1948), .Y(n1950) );
  ao211d1_hd U1196 ( .A(n1952), .B(guard), .C(n1951), .D(n1950), .Y(n1953) );
  oa211d1_hd U1197 ( .A(n1956), .B(n1955), .C(n1954), .D(n1953), .Y(n417) );
  ao21d1_hd U1198 ( .A(n1958), .B(n1968), .C(n1957), .Y(n1964) );
  oa21d1_hd U1199 ( .A(n1961), .B(n1960), .C(n1959), .Y(n1962) );
  ao22d1_hd U1200 ( .A(z_m[22]), .B(n1962), .C(n1975), .D(sum[26]), .Y(n1963)
         );
  oa211d1_hd U1201 ( .A(n1964), .B(n1967), .C(n1963), .D(n1972), .Y(n418) );
  nr4d1_hd U1202 ( .A(n1968), .B(n1967), .C(n1966), .D(n1965), .Y(n1969) );
  nd4d1_hd U1203 ( .A(z_m[21]), .B(z_m[20]), .C(n1970), .D(n1969), .Y(n1971)
         );
  nd4d1_hd U1204 ( .A(n1973), .B(n1283), .C(n1972), .D(n1971), .Y(n1987) );
  nr3d1_hd U1205 ( .A(n1975), .B(state[1]), .C(n1974), .Y(n1976) );
  ao22d1_hd U1206 ( .A(a_e[8]), .B(n1569), .C(n1993), .D(C91_DATA2_8), .Y(
        n1977) );
  oa21d1_hd U1207 ( .A(n1978), .B(n1987), .C(n1977), .Y(n419) );
  ao22d1_hd U1208 ( .A(z_e[7]), .B(n1989), .C(n1993), .D(C91_DATA2_7), .Y(
        n1979) );
  oa21d1_hd U1209 ( .A(n2104), .B(n1283), .C(n1979), .Y(n420) );
  ao22d1_hd U1210 ( .A(z_e[6]), .B(n1989), .C(n1993), .D(C91_DATA2_6), .Y(
        n1980) );
  oa21d1_hd U1211 ( .A(n2100), .B(n1283), .C(n1980), .Y(n421) );
  ao22d1_hd U1212 ( .A(z_e[5]), .B(n1989), .C(n1993), .D(C91_DATA2_5), .Y(
        n1981) );
  oa21d1_hd U1213 ( .A(n2119), .B(n1283), .C(n1981), .Y(n422) );
  ao22d1_hd U1214 ( .A(z_e[4]), .B(n1989), .C(n1993), .D(C91_DATA2_4), .Y(
        n1982) );
  oa21d1_hd U1215 ( .A(n2124), .B(n1283), .C(n1982), .Y(n423) );
  ao22d1_hd U1216 ( .A(z_e[3]), .B(n1989), .C(n1993), .D(C91_DATA2_3), .Y(
        n1983) );
  oa21d1_hd U1217 ( .A(n2131), .B(n1283), .C(n1983), .Y(n424) );
  ao22d1_hd U1218 ( .A(z_e[2]), .B(n1989), .C(n1993), .D(C91_DATA2_2), .Y(
        n1984) );
  oa21d1_hd U1219 ( .A(n2140), .B(n1283), .C(n1984), .Y(n425) );
  ao22d1_hd U1220 ( .A(z_e[1]), .B(n1989), .C(n1993), .D(C91_DATA2_1), .Y(
        n1985) );
  oa21d1_hd U1221 ( .A(n2148), .B(n1283), .C(n1985), .Y(n426) );
  ao22d1_hd U1222 ( .A(a_e[0]), .B(n1569), .C(n1993), .D(n1988), .Y(n1986) );
  oa21d1_hd U1223 ( .A(n1988), .B(n1987), .C(n1986), .Y(n427) );
  ao22d1_hd U1224 ( .A(a_e[9]), .B(n1569), .C(z_e[9]), .D(n1989), .Y(n1996) );
  ao22d1_hd U1225 ( .A(z_e[9]), .B(n1896), .C(n1991), .D(n1990), .Y(n1994) );
  oa211d1_hd U1226 ( .A(DP_OP_154J2_137_6175_n2), .B(n1994), .C(n1993), .D(
        n1992), .Y(n1995) );
  ao22d1_hd U1227 ( .A(b_m[25]), .B(n2039), .C(n1577), .D(b[21]), .Y(n1997) );
  oa21d1_hd U1228 ( .A(n1998), .B(n1575), .C(n1997), .Y(n429) );
  ao22d1_hd U1229 ( .A(b_m[24]), .B(n2039), .C(n1578), .D(b[20]), .Y(n1999) );
  oa21d1_hd U1230 ( .A(n2000), .B(n1575), .C(n1999), .Y(n430) );
  ao22d1_hd U1231 ( .A(b_m[23]), .B(n2039), .C(n1579), .D(b[19]), .Y(n2001) );
  oa21d1_hd U1232 ( .A(n2002), .B(n1575), .C(n2001), .Y(n431) );
  ao22d1_hd U1233 ( .A(b_m[22]), .B(n2039), .C(n1578), .D(b[18]), .Y(n2003) );
  oa21d1_hd U1234 ( .A(n2004), .B(n1575), .C(n2003), .Y(n432) );
  ao22d1_hd U1235 ( .A(b_m[21]), .B(n2039), .C(n1578), .D(b[17]), .Y(n2005) );
  oa21d1_hd U1236 ( .A(n2006), .B(n1575), .C(n2005), .Y(n433) );
  ao22d1_hd U1237 ( .A(b_m[20]), .B(n2039), .C(n1578), .D(b[16]), .Y(n2007) );
  oa21d1_hd U1238 ( .A(n2008), .B(n1575), .C(n2007), .Y(n434) );
  ao22d1_hd U1239 ( .A(b_m[19]), .B(n2039), .C(n1578), .D(b[15]), .Y(n2009) );
  oa21d1_hd U1240 ( .A(n2010), .B(n1575), .C(n2009), .Y(n435) );
  ao22d1_hd U1241 ( .A(b_m[18]), .B(n2039), .C(n1578), .D(b[14]), .Y(n2011) );
  oa21d1_hd U1242 ( .A(n2012), .B(n1575), .C(n2011), .Y(n436) );
  ao22d1_hd U1243 ( .A(b_m[17]), .B(n2039), .C(n1578), .D(b[13]), .Y(n2013) );
  oa21d1_hd U1244 ( .A(n2014), .B(n1575), .C(n2013), .Y(n437) );
  ao22d1_hd U1245 ( .A(b_m[16]), .B(n2039), .C(n1578), .D(b[12]), .Y(n2015) );
  oa21d1_hd U1246 ( .A(n2016), .B(n1575), .C(n2015), .Y(n438) );
  ao22d1_hd U1247 ( .A(b_m[15]), .B(n2039), .C(n1578), .D(b[11]), .Y(n2017) );
  oa21d1_hd U1248 ( .A(n2018), .B(n1575), .C(n2017), .Y(n439) );
  ao22d1_hd U1249 ( .A(b_m[14]), .B(n2039), .C(n1578), .D(b[10]), .Y(n2019) );
  oa21d1_hd U1250 ( .A(n2020), .B(n1575), .C(n2019), .Y(n440) );
  ao22d1_hd U1251 ( .A(b_m[13]), .B(n2039), .C(n1578), .D(b[9]), .Y(n2021) );
  oa21d1_hd U1252 ( .A(n2022), .B(n1575), .C(n2021), .Y(n441) );
  ao22d1_hd U1253 ( .A(b_m[12]), .B(n2039), .C(n1578), .D(b[8]), .Y(n2023) );
  oa21d1_hd U1254 ( .A(n2024), .B(n1575), .C(n2023), .Y(n442) );
  ao22d1_hd U1255 ( .A(b_m[11]), .B(n2039), .C(n1578), .D(b[7]), .Y(n2025) );
  oa21d1_hd U1256 ( .A(n2026), .B(n1575), .C(n2025), .Y(n443) );
  ao22d1_hd U1257 ( .A(b_m[10]), .B(n2039), .C(n1578), .D(b[6]), .Y(n2027) );
  oa21d1_hd U1258 ( .A(n2028), .B(n1575), .C(n2027), .Y(n444) );
  ao22d1_hd U1259 ( .A(b_m[9]), .B(n2039), .C(n1578), .D(b[5]), .Y(n2029) );
  oa21d1_hd U1260 ( .A(n2030), .B(n1575), .C(n2029), .Y(n445) );
  ao22d1_hd U1261 ( .A(b_m[8]), .B(n2039), .C(n1578), .D(b[4]), .Y(n2031) );
  oa21d1_hd U1262 ( .A(n2032), .B(n1575), .C(n2031), .Y(n446) );
  ao22d1_hd U1263 ( .A(b_m[7]), .B(n2039), .C(n1578), .D(b[3]), .Y(n2033) );
  oa21d1_hd U1264 ( .A(n2034), .B(n1575), .C(n2033), .Y(n447) );
  ao22d1_hd U1265 ( .A(b_m[6]), .B(n2039), .C(n1578), .D(b[2]), .Y(n2035) );
  oa21d1_hd U1266 ( .A(n2036), .B(n1575), .C(n2035), .Y(n448) );
  ao22d1_hd U1267 ( .A(b_m[5]), .B(n2039), .C(n1578), .D(b[1]), .Y(n2037) );
  oa21d1_hd U1268 ( .A(n2038), .B(n1575), .C(n2037), .Y(n449) );
  ao22d1_hd U1269 ( .A(b_m[4]), .B(n2039), .C(n1578), .D(b[0]), .Y(n2040) );
  oa21d1_hd U1270 ( .A(n2041), .B(n1575), .C(n2040), .Y(n450) );
  oa22d1_hd U1271 ( .A(n2042), .B(n1575), .C(n2041), .D(n2252), .Y(n451) );
  oa22d1_hd U1272 ( .A(n2043), .B(n1575), .C(n2042), .D(n2252), .Y(n452) );
  oa22d1_hd U1273 ( .A(n1579), .B(n2044), .C(n2043), .D(n2252), .Y(n453) );
  ao22d1_hd U1274 ( .A(a_m[25]), .B(n2087), .C(n1578), .D(a[21]), .Y(n2045) );
  oa21d1_hd U1275 ( .A(n2046), .B(n1573), .C(n2045), .Y(n454) );
  ao22d1_hd U1276 ( .A(a_m[24]), .B(n2087), .C(n1578), .D(a[20]), .Y(n2047) );
  oa21d1_hd U1277 ( .A(n2048), .B(n1573), .C(n2047), .Y(n455) );
  ao22d1_hd U1278 ( .A(a_m[23]), .B(n2087), .C(n1578), .D(a[19]), .Y(n2049) );
  oa21d1_hd U1279 ( .A(n2050), .B(n1573), .C(n2049), .Y(n456) );
  ao22d1_hd U1280 ( .A(a_m[22]), .B(n2087), .C(n1578), .D(a[18]), .Y(n2051) );
  oa21d1_hd U1281 ( .A(n2052), .B(n1573), .C(n2051), .Y(n457) );
  ao22d1_hd U1282 ( .A(a_m[21]), .B(n2087), .C(n1578), .D(a[17]), .Y(n2053) );
  oa21d1_hd U1283 ( .A(n2054), .B(n1573), .C(n2053), .Y(n458) );
  ao22d1_hd U1284 ( .A(a_m[20]), .B(n2087), .C(n1579), .D(a[16]), .Y(n2055) );
  oa21d1_hd U1285 ( .A(n2056), .B(n1573), .C(n2055), .Y(n459) );
  ao22d1_hd U1286 ( .A(a_m[19]), .B(n2087), .C(n1578), .D(a[15]), .Y(n2057) );
  oa21d1_hd U1287 ( .A(n2058), .B(n1573), .C(n2057), .Y(n460) );
  ao22d1_hd U1288 ( .A(a_m[18]), .B(n2087), .C(n1578), .D(a[14]), .Y(n2059) );
  oa21d1_hd U1289 ( .A(n2060), .B(n1573), .C(n2059), .Y(n461) );
  ao22d1_hd U1290 ( .A(a_m[17]), .B(n2087), .C(n1579), .D(a[13]), .Y(n2061) );
  oa21d1_hd U1291 ( .A(n2062), .B(n1573), .C(n2061), .Y(n462) );
  ao22d1_hd U1292 ( .A(a_m[16]), .B(n2087), .C(n1578), .D(a[12]), .Y(n2063) );
  oa21d1_hd U1293 ( .A(n2064), .B(n1573), .C(n2063), .Y(n463) );
  ao22d1_hd U1294 ( .A(a_m[15]), .B(n2087), .C(n1579), .D(a[11]), .Y(n2065) );
  oa21d1_hd U1295 ( .A(n2066), .B(n1573), .C(n2065), .Y(n464) );
  ao22d1_hd U1296 ( .A(a_m[14]), .B(n2087), .C(n1577), .D(a[10]), .Y(n2067) );
  oa21d1_hd U1297 ( .A(n2068), .B(n1573), .C(n2067), .Y(n465) );
  ao22d1_hd U1298 ( .A(a_m[13]), .B(n2087), .C(n1577), .D(a[9]), .Y(n2069) );
  oa21d1_hd U1299 ( .A(n2070), .B(n1573), .C(n2069), .Y(n466) );
  ao22d1_hd U1300 ( .A(a_m[12]), .B(n2087), .C(n1577), .D(a[8]), .Y(n2071) );
  oa21d1_hd U1301 ( .A(n2072), .B(n1573), .C(n2071), .Y(n467) );
  ao22d1_hd U1302 ( .A(a_m[11]), .B(n2087), .C(n1577), .D(a[7]), .Y(n2073) );
  oa21d1_hd U1303 ( .A(n2074), .B(n1573), .C(n2073), .Y(n468) );
  ao22d1_hd U1304 ( .A(a_m[10]), .B(n2087), .C(n1577), .D(a[6]), .Y(n2075) );
  oa21d1_hd U1305 ( .A(n2076), .B(n1573), .C(n2075), .Y(n469) );
  ao22d1_hd U1306 ( .A(a_m[9]), .B(n2087), .C(n1577), .D(a[5]), .Y(n2077) );
  oa21d1_hd U1307 ( .A(n2078), .B(n1573), .C(n2077), .Y(n470) );
  ao22d1_hd U1308 ( .A(a_m[8]), .B(n2087), .C(n1577), .D(a[4]), .Y(n2079) );
  oa21d1_hd U1309 ( .A(n2080), .B(n1573), .C(n2079), .Y(n471) );
  ao22d1_hd U1310 ( .A(a_m[7]), .B(n2087), .C(n1577), .D(a[3]), .Y(n2081) );
  oa21d1_hd U1311 ( .A(n2082), .B(n1573), .C(n2081), .Y(n472) );
  ao22d1_hd U1312 ( .A(a_m[6]), .B(n2087), .C(n1578), .D(a[2]), .Y(n2083) );
  oa21d1_hd U1313 ( .A(n2084), .B(n1573), .C(n2083), .Y(n473) );
  ao22d1_hd U1314 ( .A(a_m[5]), .B(n2087), .C(n1577), .D(a[1]), .Y(n2085) );
  oa21d1_hd U1315 ( .A(n2086), .B(n1573), .C(n2085), .Y(n474) );
  ao22d1_hd U1316 ( .A(a_m[4]), .B(n2087), .C(n1577), .D(a[0]), .Y(n2088) );
  oa21d1_hd U1317 ( .A(n2089), .B(n1573), .C(n2088), .Y(n475) );
  oa22d1_hd U1318 ( .A(n2090), .B(n1573), .C(n2089), .D(n2094), .Y(n476) );
  oa22d1_hd U1319 ( .A(n2091), .B(n1573), .C(n2090), .D(n2094), .Y(n477) );
  oa22d1_hd U1320 ( .A(n1579), .B(n2092), .C(n2091), .D(n2094), .Y(n478) );
  ao22d1_hd U1321 ( .A(a_m[25]), .B(n1574), .C(n1577), .D(a[22]), .Y(n2093) );
  oa21d1_hd U1322 ( .A(n2095), .B(n2094), .C(n2093), .Y(n479) );
  nr2d1_hd U1323 ( .A(n2148), .B(n2147), .Y(n2136) );
  nr2d1_hd U1324 ( .A(n2131), .B(n2130), .Y(n2121) );
  ao21d1_hd U1325 ( .A(n2189), .B(n2099), .C(n2154), .Y(n2120) );
  oa21d1_hd U1326 ( .A(n2100), .B(n2119), .C(n2189), .Y(n2098) );
  ao21d1_hd U1327 ( .A(n2139), .B(n2104), .C(n2106), .Y(n2156) );
  ivd1_hd U1328 ( .A(a[25]), .Y(n2138) );
  nr2d1_hd U1329 ( .A(n2150), .B(n2138), .Y(n2137) );
  ivd1_hd U1330 ( .A(a[27]), .Y(n2123) );
  nr2d1_hd U1331 ( .A(n2133), .B(n2123), .Y(n2122) );
  ivd1_hd U1332 ( .A(a[29]), .Y(n2109) );
  nr2d1_hd U1333 ( .A(n2116), .B(n2109), .Y(n2103) );
  nr2d1_hd U1334 ( .A(n2103), .B(n1897), .Y(n2111) );
  nr2d1_hd U1335 ( .A(n2157), .B(n2099), .Y(n2115) );
  nr2d1_hd U1336 ( .A(n2100), .B(n2114), .Y(n2105) );
  nd3d1_hd U1337 ( .A(a_e[7]), .B(n2105), .C(n2102), .Y(n2101) );
  oa211d1_hd U1338 ( .A(n2156), .B(n2102), .C(n2158), .D(n2101), .Y(n480) );
  ao22d1_hd U1339 ( .A(a_e[7]), .B(n2106), .C(n2105), .D(n2104), .Y(n2107) );
  oa211d1_hd U1340 ( .A(n1897), .B(n2108), .C(n2107), .D(n2158), .Y(n481) );
  oa21d1_hd U1341 ( .A(a_e[5]), .B(n2157), .C(n2120), .Y(n2112) );
  ao22d1_hd U1342 ( .A(a_e[6]), .B(n2112), .C(n2111), .D(n2110), .Y(n2113) );
  oa211d1_hd U1343 ( .A(a_e[6]), .B(n2114), .C(n2113), .D(n2143), .Y(n482) );
  ao21d1_hd U1344 ( .A(n2115), .B(n2119), .C(n2159), .Y(n2118) );
  oa211d1_hd U1345 ( .A(n2122), .B(a[28]), .C(n1579), .D(n2116), .Y(n2117) );
  oa211d1_hd U1346 ( .A(n2120), .B(n2119), .C(n2118), .D(n2117), .Y(n483) );
  ao211d1_hd U1347 ( .A(n2133), .B(n2123), .C(n2122), .D(n1897), .Y(n2126) );
  ao21d1_hd U1348 ( .A(n2189), .B(n2130), .C(n2154), .Y(n2132) );
  ao21d1_hd U1349 ( .A(n2132), .B(n2129), .C(n2124), .Y(n2125) );
  nr2d1_hd U1350 ( .A(n2126), .B(n2125), .Y(n2127) );
  oa211d1_hd U1351 ( .A(a_e[4]), .B(n2128), .C(n2127), .D(n2143), .Y(n484) );
  oa22d1_hd U1352 ( .A(n2132), .B(n2131), .C(n2130), .D(n2129), .Y(n2135) );
  oa211d1_hd U1353 ( .A(n2137), .B(a[26]), .C(n1579), .D(n2133), .Y(n2134) );
  scg13d1_hd U1354 ( .A(n2135), .B(n2159), .C(n2134), .Y(n485) );
  ao211d1_hd U1355 ( .A(n2150), .B(n2138), .C(n2137), .D(n1897), .Y(n2142) );
  nr2d1_hd U1356 ( .A(a_e[0]), .B(n2157), .Y(n2153) );
  nr2d1_hd U1357 ( .A(n2154), .B(n2153), .Y(n2149) );
  ao21d1_hd U1358 ( .A(n2149), .B(n2146), .C(n2140), .Y(n2141) );
  nr2d1_hd U1359 ( .A(n2142), .B(n2141), .Y(n2144) );
  oa211d1_hd U1360 ( .A(a_e[2]), .B(n2145), .C(n2144), .D(n2143), .Y(n486) );
  oa22d1_hd U1361 ( .A(n2149), .B(n2148), .C(n2147), .D(n2146), .Y(n2152) );
  oa211d1_hd U1362 ( .A(a[23]), .B(a[24]), .C(n1579), .D(n2150), .Y(n2151) );
  scg13d1_hd U1363 ( .A(n2152), .B(n2159), .C(n2151), .Y(n487) );
  ao21d1_hd U1364 ( .A(n2154), .B(a_e[0]), .C(n2153), .Y(n2155) );
  oa21d1_hd U1365 ( .A(a[23]), .B(n1897), .C(n2155), .Y(n488) );
  oa21d1_hd U1366 ( .A(a_e[8]), .B(n2157), .C(n2156), .Y(n2160) );
  scg17d1_hd U1367 ( .A(a_e[9]), .B(n2160), .C(n2159), .D(n2158), .Y(n489) );
  nr2d1_hd U1368 ( .A(n2215), .B(n2214), .Y(n2204) );
  nr2d1_hd U1369 ( .A(n2164), .B(n2198), .Y(n2194) );
  ao21d1_hd U1370 ( .A(n2165), .B(n2189), .C(n2221), .Y(n2188) );
  oa21d1_hd U1371 ( .A(n2167), .B(n2187), .C(n2189), .Y(n2166) );
  ao21d1_hd U1372 ( .A(n2205), .B(n2171), .C(n2173), .Y(n2254) );
  ivd1_hd U1373 ( .A(b[25]), .Y(n2207) );
  nr2d1_hd U1374 ( .A(n2217), .B(n2207), .Y(n2206) );
  ivd1_hd U1375 ( .A(b[27]), .Y(n2191) );
  nr2d1_hd U1376 ( .A(n2201), .B(n2191), .Y(n2190) );
  ivd1_hd U1377 ( .A(b[29]), .Y(n2177) );
  nr2d1_hd U1378 ( .A(n2184), .B(n2177), .Y(n2170) );
  nr2d1_hd U1379 ( .A(n2170), .B(n1897), .Y(n2180) );
  nr2bd1_hd U1380 ( .AN(n2194), .B(n2197), .Y(n2183) );
  nr2d1_hd U1381 ( .A(n2167), .B(n2182), .Y(n2172) );
  nd3d1_hd U1382 ( .A(b_e[7]), .B(n2172), .C(n2169), .Y(n2168) );
  oa211d1_hd U1383 ( .A(n2254), .B(n2169), .C(n2256), .D(n2168), .Y(n490) );
  ao22d1_hd U1384 ( .A(b_e[7]), .B(n2173), .C(n2172), .D(n2171), .Y(n2174) );
  oa211d1_hd U1385 ( .A(n2176), .B(n2175), .C(n2174), .D(n2256), .Y(n491) );
  oa21d1_hd U1386 ( .A(b_e[5]), .B(n2255), .C(n2188), .Y(n2178) );
  ao22d1_hd U1387 ( .A(n2180), .B(n2179), .C(b_e[6]), .D(n2178), .Y(n2181) );
  oa211d1_hd U1388 ( .A(b_e[6]), .B(n2182), .C(n2181), .D(n2210), .Y(n492) );
  ao21d1_hd U1389 ( .A(n2183), .B(n2187), .C(n2257), .Y(n2186) );
  oa211d1_hd U1390 ( .A(n2190), .B(b[28]), .C(n1579), .D(n2184), .Y(n2185) );
  oa211d1_hd U1391 ( .A(n2188), .B(n2187), .C(n2186), .D(n2185), .Y(n493) );
  scg6d1_hd U1392 ( .A(n2198), .B(n2189), .C(n2221), .Y(n2200) );
  ao211d1_hd U1393 ( .A(n2201), .B(n2191), .C(n2190), .D(n1897), .Y(n2192) );
  ao211d1_hd U1394 ( .A(b_e[4]), .B(n2200), .C(n2257), .D(n2192), .Y(n2196) );
  nd3d1_hd U1395 ( .A(n2205), .B(n2194), .C(n2193), .Y(n2195) );
  oa211d1_hd U1396 ( .A(b_e[3]), .B(n2197), .C(n2196), .D(n2195), .Y(n494) );
  nr3d1_hd U1397 ( .A(b_e[3]), .B(n2255), .C(n2198), .Y(n2199) );
  ao211d1_hd U1398 ( .A(b_e[3]), .B(n2200), .C(n2257), .D(n2199), .Y(n2203) );
  oa211d1_hd U1399 ( .A(n2206), .B(b[26]), .C(n1579), .D(n2201), .Y(n2202) );
  nr2d1_hd U1400 ( .A(b_e[0]), .B(n2255), .Y(n2220) );
  nr2d1_hd U1401 ( .A(n2221), .B(n2220), .Y(n2216) );
  ao211d1_hd U1402 ( .A(n2217), .B(n2207), .C(n2206), .D(n1897), .Y(n2208) );
  ao21d1_hd U1403 ( .A(n2209), .B(b_e[2]), .C(n2208), .Y(n2211) );
  oa211d1_hd U1404 ( .A(b_e[2]), .B(n2212), .C(n2211), .D(n2210), .Y(n496) );
  oa22d1_hd U1405 ( .A(n2216), .B(n2215), .C(n2214), .D(n2213), .Y(n2219) );
  oa211d1_hd U1406 ( .A(b[23]), .B(b[24]), .C(n1579), .D(n2217), .Y(n2218) );
  scg13d1_hd U1407 ( .A(n2219), .B(n2257), .C(n2218), .Y(n497) );
  ao21d1_hd U1408 ( .A(n2221), .B(b_e[0]), .C(n2220), .Y(n2222) );
  oa21d1_hd U1409 ( .A(b[23]), .B(n1897), .C(n2222), .Y(n498) );
  scg21d1_hd U1410 ( .A(n2223), .B(o_AB_ACK), .C(i_RST), .D(n1570), .Y(n499)
         );
  oa211d1_hd U1411 ( .A(state[3]), .B(n2228), .C(n2227), .D(n2226), .Y(n2242)
         );
  nd3d1_hd U1412 ( .A(n1580), .B(o_Z_STB), .C(i_Z_ACK), .Y(n2266) );
  nd4d1_hd U1413 ( .A(N41), .B(n2261), .C(n2266), .D(n1283), .Y(n2229) );
  nr3d1_hd U1414 ( .A(n27), .B(n2242), .C(n2229), .Y(n2234) );
  ao22d1_hd U1415 ( .A(n2232), .B(n2231), .C(n1896), .D(n2230), .Y(n2233) );
  oa211d1_hd U1416 ( .A(n2236), .B(n2235), .C(n2234), .D(n2233), .Y(n2262) );
  ivd1_hd U1417 ( .A(n2262), .Y(n2239) );
  nr2d1_hd U1418 ( .A(n2237), .B(n2247), .Y(n2238) );
  ao22d1_hd U1419 ( .A(state[2]), .B(n2239), .C(N41), .D(n2238), .Y(n2240) );
  oa21d1_hd U1420 ( .A(n2241), .B(n2264), .C(n2240), .Y(n500) );
  nr2d1_hd U1421 ( .A(n1896), .B(n2242), .Y(n2244) );
  oa22d1_hd U1422 ( .A(n2244), .B(n2264), .C(n2243), .D(n2262), .Y(n501) );
  oa211d1_hd U1423 ( .A(n2247), .B(state[0]), .C(n2246), .D(n2245), .Y(n2248)
         );
  ivd1_hd U1424 ( .A(n2248), .Y(n2250) );
  oa22d1_hd U1425 ( .A(n2250), .B(n2264), .C(n2249), .D(n2262), .Y(n502) );
  ao22d1_hd U1426 ( .A(b_m[25]), .B(n2161), .C(n1577), .D(b[22]), .Y(n2251) );
  oa21d1_hd U1427 ( .A(n2253), .B(n2252), .C(n2251), .Y(n503) );
  oa21d1_hd U1428 ( .A(b_e[8]), .B(n2255), .C(n2254), .Y(n2258) );
  scg17d1_hd U1429 ( .A(b_e[9]), .B(n2258), .C(n2257), .D(n2256), .Y(n504) );
  oa22d1_hd U1430 ( .A(n2265), .B(n2264), .C(n2263), .D(n2262), .Y(n505) );
  ivd1_hd U1431 ( .A(n2266), .Y(n2267) );
  scg21d1_hd U1432 ( .A(n1580), .B(o_Z_STB), .C(i_RST), .D(n2267), .Y(n506) );
endmodule


module float_adder_0 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3, C91_DATA2_4,
         C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8, n1, n2, n27, n265,
         n266, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n509, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23,
         C2_Z_22, C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16,
         C2_Z_15, C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_43J2_124_6938_n58, DP_OP_43J2_124_6938_n57,
         DP_OP_43J2_124_6938_n56, DP_OP_43J2_124_6938_n55,
         DP_OP_43J2_124_6938_n54, DP_OP_43J2_124_6938_n53,
         DP_OP_43J2_124_6938_n52, DP_OP_43J2_124_6938_n51,
         DP_OP_43J2_124_6938_n50, DP_OP_43J2_124_6938_n49,
         DP_OP_43J2_124_6938_n48, DP_OP_43J2_124_6938_n47,
         DP_OP_43J2_124_6938_n46, DP_OP_43J2_124_6938_n45,
         DP_OP_43J2_124_6938_n44, DP_OP_43J2_124_6938_n43,
         DP_OP_43J2_124_6938_n42, DP_OP_43J2_124_6938_n41,
         DP_OP_43J2_124_6938_n40, DP_OP_43J2_124_6938_n39,
         DP_OP_43J2_124_6938_n38, DP_OP_43J2_124_6938_n37,
         DP_OP_43J2_124_6938_n36, DP_OP_43J2_124_6938_n35,
         DP_OP_43J2_124_6938_n34, DP_OP_43J2_124_6938_n33,
         DP_OP_43J2_124_6938_n32, DP_OP_43J2_124_6938_n27,
         DP_OP_43J2_124_6938_n26, DP_OP_43J2_124_6938_n25,
         DP_OP_43J2_124_6938_n24, DP_OP_43J2_124_6938_n23,
         DP_OP_43J2_124_6938_n22, DP_OP_43J2_124_6938_n21,
         DP_OP_43J2_124_6938_n20, DP_OP_43J2_124_6938_n19,
         DP_OP_43J2_124_6938_n18, DP_OP_43J2_124_6938_n17,
         DP_OP_43J2_124_6938_n16, DP_OP_43J2_124_6938_n15,
         DP_OP_43J2_124_6938_n14, DP_OP_43J2_124_6938_n13,
         DP_OP_43J2_124_6938_n12, DP_OP_43J2_124_6938_n11,
         DP_OP_43J2_124_6938_n10, DP_OP_43J2_124_6938_n9,
         DP_OP_43J2_124_6938_n8, DP_OP_43J2_124_6938_n7,
         DP_OP_43J2_124_6938_n6, DP_OP_43J2_124_6938_n5,
         DP_OP_43J2_124_6938_n4, DP_OP_43J2_124_6938_n3,
         DP_OP_43J2_124_6938_n2, DP_OP_43J2_124_6938_n1,
         DP_OP_154J2_137_6175_n9, DP_OP_154J2_137_6175_n8,
         DP_OP_154J2_137_6175_n7, DP_OP_154J2_137_6175_n6,
         DP_OP_154J2_137_6175_n5, DP_OP_154J2_137_6175_n4,
         DP_OP_154J2_137_6175_n3, DP_OP_154J2_137_6175_n2, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J2_137_6175_U10 ( .A(n2269), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J2_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J2_137_6175_U9 ( .A(n2269), .B(z_e[2]), .CI(
        DP_OP_154J2_137_6175_n9), .CO(DP_OP_154J2_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J2_137_6175_U8 ( .A(n2269), .B(z_e[3]), .CI(
        DP_OP_154J2_137_6175_n8), .CO(DP_OP_154J2_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J2_137_6175_U7 ( .A(n2269), .B(z_e[4]), .CI(
        DP_OP_154J2_137_6175_n7), .CO(DP_OP_154J2_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J2_137_6175_U6 ( .A(n2269), .B(z_e[5]), .CI(
        DP_OP_154J2_137_6175_n6), .CO(DP_OP_154J2_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J2_137_6175_U5 ( .A(n2269), .B(z_e[6]), .CI(
        DP_OP_154J2_137_6175_n5), .CO(DP_OP_154J2_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J2_137_6175_U4 ( .A(n2269), .B(z_e[7]), .CI(
        DP_OP_154J2_137_6175_n4), .CO(DP_OP_154J2_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J2_137_6175_U3 ( .A(n2269), .B(z_e[8]), .CI(
        DP_OP_154J2_137_6175_n3), .CO(DP_OP_154J2_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1580), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n509), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n509), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1580), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1580), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1580), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1580), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1580), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n1580), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n1580), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n1580), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n1580), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n1580), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n1580), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n1580), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n1580), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1580), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1580), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1580), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1580), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1580), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n509), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n509), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n509), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n509), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1580), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1580), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n1580), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1580), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1580), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1580), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n1570), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n1570), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n1570), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n1570), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n1569), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n1569), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n1570), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n1570), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n1570), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n1570), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n1570), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n1570), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n1570), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n1570), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n1570), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n1570), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n1570), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n1570), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n1570), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n1570), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n1570), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n1570), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n1570), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n1570), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n1570), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n1570), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n1570), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n1570), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n1570), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n1570), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n1570), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n1570), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n1570), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n1570), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n1570), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n1570), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n1570), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n1570), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n1570), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n1570), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n1570), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n1570), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n1570), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n1570), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n1570), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n1570), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n1570), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n1570), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n1570), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n1570), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n1570), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n1570), .CK(i_CLK), .Q(b[22]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n1569), .CK(i_CLK), .Q(sum[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n1569), .CK(i_CLK), .Q(sum[2]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n1569), .CK(i_CLK), .Q(sum[26]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n1569), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n1569), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n1569), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n1569), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n1569), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n1569), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n1569), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n1569), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n1569), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n1569), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n1569), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n1569), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n1569), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n1569), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n1569), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n1569), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n1569), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n1569), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n1569), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n1569), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n1569), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n1569), .CK(i_CLK), .Q(sum[25]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n1569), .CK(i_CLK), .Q(sum[1]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n1570), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n1570), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n1570), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n1570), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n1569), .CK(i_CLK), .Q(sum[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n1570), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n1570), .CK(i_CLK), .Q(b[28]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n1570), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n1570), .CK(i_CLK), .Q(b[25]) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n1570), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n1570), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n1570), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n1570), .CK(i_CLK), .Q(b[26]) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n1570), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n1570), .CK(i_CLK), .Q(b[23]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n265), .CK(i_CLK), .Q(guard) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1577), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1577), .CK(i_CLK), .Q(a_s) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n2270), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n2270), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J2_124_6938_U28 ( .A(C2_Z_0), .B(n2271), .CI(
        DP_OP_43J2_124_6938_n58), .CO(DP_OP_43J2_124_6938_n27), .S(N310) );
  fad1_hd DP_OP_43J2_124_6938_U27 ( .A(DP_OP_43J2_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J2_124_6938_n27), .CO(DP_OP_43J2_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J2_124_6938_U26 ( .A(DP_OP_43J2_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J2_124_6938_n26), .CO(DP_OP_43J2_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J2_124_6938_U25 ( .A(DP_OP_43J2_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J2_124_6938_n25), .CO(DP_OP_43J2_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J2_124_6938_U24 ( .A(DP_OP_43J2_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J2_124_6938_n24), .CO(DP_OP_43J2_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J2_124_6938_U23 ( .A(DP_OP_43J2_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J2_124_6938_n23), .CO(DP_OP_43J2_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J2_124_6938_U2 ( .A(DP_OP_43J2_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J2_124_6938_n2), .CO(DP_OP_43J2_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J2_124_6938_U3 ( .A(DP_OP_43J2_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J2_124_6938_n3), .CO(DP_OP_43J2_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J2_124_6938_U4 ( .A(DP_OP_43J2_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J2_124_6938_n4), .CO(DP_OP_43J2_124_6938_n3), .S(N334) );
  fad1_hd DP_OP_43J2_124_6938_U5 ( .A(DP_OP_43J2_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J2_124_6938_n5), .CO(DP_OP_43J2_124_6938_n4), .S(N333) );
  fad1_hd DP_OP_43J2_124_6938_U6 ( .A(DP_OP_43J2_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J2_124_6938_n6), .CO(DP_OP_43J2_124_6938_n5), .S(N332) );
  fad1_hd DP_OP_43J2_124_6938_U7 ( .A(DP_OP_43J2_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J2_124_6938_n7), .CO(DP_OP_43J2_124_6938_n6), .S(N331) );
  fad1_hd DP_OP_43J2_124_6938_U8 ( .A(DP_OP_43J2_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J2_124_6938_n8), .CO(DP_OP_43J2_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J2_124_6938_U9 ( .A(DP_OP_43J2_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J2_124_6938_n9), .CO(DP_OP_43J2_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J2_124_6938_U10 ( .A(DP_OP_43J2_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J2_124_6938_n10), .CO(DP_OP_43J2_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J2_124_6938_U11 ( .A(DP_OP_43J2_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J2_124_6938_n11), .CO(DP_OP_43J2_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J2_124_6938_U12 ( .A(DP_OP_43J2_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J2_124_6938_n12), .CO(DP_OP_43J2_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J2_124_6938_U13 ( .A(DP_OP_43J2_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J2_124_6938_n13), .CO(DP_OP_43J2_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J2_124_6938_U14 ( .A(DP_OP_43J2_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J2_124_6938_n14), .CO(DP_OP_43J2_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J2_124_6938_U15 ( .A(DP_OP_43J2_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J2_124_6938_n15), .CO(DP_OP_43J2_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J2_124_6938_U16 ( .A(DP_OP_43J2_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J2_124_6938_n16), .CO(DP_OP_43J2_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J2_124_6938_U17 ( .A(DP_OP_43J2_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J2_124_6938_n17), .CO(DP_OP_43J2_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J2_124_6938_U18 ( .A(DP_OP_43J2_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J2_124_6938_n18), .CO(DP_OP_43J2_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J2_124_6938_U19 ( .A(DP_OP_43J2_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J2_124_6938_n19), .CO(DP_OP_43J2_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J2_124_6938_U20 ( .A(DP_OP_43J2_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J2_124_6938_n20), .CO(DP_OP_43J2_124_6938_n19), .S(N318)
         );
  fad1_hd DP_OP_43J2_124_6938_U21 ( .A(DP_OP_43J2_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J2_124_6938_n21), .CO(DP_OP_43J2_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J2_124_6938_U22 ( .A(DP_OP_43J2_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J2_124_6938_n22), .CO(DP_OP_43J2_124_6938_n21), .S(N316)
         );
  fd1qd1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK) );
  nr2d1_hd U523 ( .A(n1991), .B(n1935), .Y(n1952) );
  clknd2d1_hd U524 ( .A(b_m[5]), .B(n2084), .Y(n1587) );
  clknd2d1_hd U525 ( .A(n1595), .B(n1594), .Y(n1596) );
  clknd2d1_hd U526 ( .A(b_m[18]), .B(n1611), .Y(n1612) );
  clknd2d1_hd U527 ( .A(b_m[8]), .B(n2078), .Y(n1592) );
  clknd2d1_hd U528 ( .A(n1590), .B(b_m[7]), .Y(n1591) );
  clknd2d1_hd U529 ( .A(b_m[12]), .B(n2070), .Y(n1600) );
  clknd2d1_hd U530 ( .A(b_m[11]), .B(n1598), .Y(n1599) );
  clknd2d1_hd U531 ( .A(b_m[17]), .B(n2060), .Y(n1610) );
  clknd2d1_hd U532 ( .A(b_e[8]), .B(n2102), .Y(n1697) );
  clknd2d1_hd U533 ( .A(n1680), .B(n1679), .Y(n1688) );
  clknd2d1_hd U534 ( .A(b_e[6]), .B(n2100), .Y(n1679) );
  clknd2d1_hd U535 ( .A(a_e[9]), .B(n1683), .Y(n1700) );
  clknd2d1_hd U536 ( .A(b_m[19]), .B(n2056), .Y(n1613) );
  clknd2d1_hd U537 ( .A(n1700), .B(n1699), .Y(n1701) );
  clknd2d1_hd U538 ( .A(a_e[8]), .B(n2169), .Y(n1694) );
  clknd2d1_hd U539 ( .A(n2189), .B(n1701), .Y(n2235) );
  clknd2d1_hd U540 ( .A(n1705), .B(n1727), .Y(n2231) );
  clknd2d1_hd U541 ( .A(n1712), .B(n2097), .Y(n1715) );
  clknd2d1_hd U542 ( .A(n1703), .B(z_e[1]), .Y(n1727) );
  clknd2d1_hd U543 ( .A(n1717), .B(n1715), .Y(n1719) );
  clknd2d1_hd U544 ( .A(n1750), .B(n1792), .Y(n1716) );
  clknd2d1_hd U545 ( .A(n2163), .B(n1711), .Y(n1717) );
  clknd2d1_hd U546 ( .A(a_e[4]), .B(n2121), .Y(n2099) );
  clknd2d1_hd U547 ( .A(state[0]), .B(n2243), .Y(n2228) );
  clknd2d1_hd U548 ( .A(n1974), .B(guard), .Y(n1966) );
  clknd2d1_hd U549 ( .A(n1575), .B(n2189), .Y(n2252) );
  clknd2d1_hd U550 ( .A(n1718), .B(n2263), .Y(n1707) );
  clknd2d1_hd U551 ( .A(n1573), .B(n2189), .Y(n2094) );
  clknd2d1_hd U552 ( .A(n2188), .B(n2166), .Y(n2173) );
  clknd2d1_hd U553 ( .A(n2249), .B(n2243), .Y(n2246) );
  clknd2d1_hd U554 ( .A(n2205), .B(n2215), .Y(n2213) );
  clknd2d1_hd U555 ( .A(b_e[2]), .B(n2204), .Y(n2198) );
  clknd2d1_hd U556 ( .A(a_e[2]), .B(n2136), .Y(n2130) );
  clknd2d1_hd U557 ( .A(n2139), .B(n2131), .Y(n2129) );
  clknd2d1_hd U558 ( .A(n2139), .B(n2148), .Y(n2146) );
  clknd2d1_hd U559 ( .A(n2120), .B(n2098), .Y(n2106) );
  clknd2d1_hd U560 ( .A(n2180), .B(n2176), .Y(n2256) );
  clknd2d1_hd U561 ( .A(b_e[5]), .B(n2183), .Y(n2182) );
  clknd2d1_hd U562 ( .A(n2194), .B(b_e[4]), .Y(n2165) );
  clknd2d1_hd U563 ( .A(n2190), .B(b[28]), .Y(n2184) );
  clknd2d1_hd U564 ( .A(state[2]), .B(n2263), .Y(n2247) );
  clknd2d1_hd U565 ( .A(N41), .B(n2262), .Y(n2264) );
  clknd2d1_hd U566 ( .A(n1958), .B(n1949), .Y(n1940) );
  clknd2d1_hd U567 ( .A(n1945), .B(n1940), .Y(n1936) );
  clknd2d1_hd U568 ( .A(n1958), .B(n1921), .Y(n1928) );
  clknd2d1_hd U569 ( .A(z_m[21]), .B(n1967), .Y(n1960) );
  clknd2d1_hd U570 ( .A(n1975), .B(sum[27]), .Y(n1972) );
  clknd2d1_hd U571 ( .A(n1958), .B(n1893), .Y(n1903) );
  clknd2d1_hd U572 ( .A(n1958), .B(n1869), .Y(n1876) );
  clknd2d1_hd U573 ( .A(n1958), .B(n1970), .Y(n1827) );
  clknd2d1_hd U574 ( .A(n1958), .B(n1845), .Y(n1852) );
  clknd2d1_hd U575 ( .A(z_m[20]), .B(n1823), .Y(n1961) );
  clknd2d1_hd U576 ( .A(z_m[19]), .B(z_m[20]), .Y(n1813) );
  clknd2d1_hd U577 ( .A(n2193), .B(n2124), .Y(n1758) );
  clknd2d1_hd U578 ( .A(n2167), .B(n2100), .Y(n1743) );
  clknd2d1_hd U579 ( .A(b_e[0]), .B(a_e[0]), .Y(n1786) );
  clknd2d1_hd U580 ( .A(n1751), .B(n1750), .Y(n1779) );
  clknd2d1_hd U581 ( .A(n1778), .B(n1773), .Y(n1772) );
  clknd2d1_hd U582 ( .A(n1764), .B(n1760), .Y(n1759) );
  clknd2d1_hd U583 ( .A(b_e[7]), .B(a_e[7]), .Y(n1738) );
  clknd2d1_hd U584 ( .A(n1749), .B(n1745), .Y(n1744) );
  clknd2d1_hd U585 ( .A(n1796), .B(n1735), .Y(n1790) );
  clknd2d1_hd U586 ( .A(n1726), .B(n1725), .Y(n1729) );
  clknd2d1_hd U587 ( .A(state[1]), .B(n2249), .Y(n2225) );
  clknd2d1_hd U588 ( .A(state[3]), .B(n1718), .Y(n2224) );
  clknd2d1_hd U589 ( .A(a[23]), .B(a[24]), .Y(n2150) );
  clknd2d1_hd U590 ( .A(n2137), .B(a[26]), .Y(n2133) );
  clknd2d1_hd U591 ( .A(b[23]), .B(b[24]), .Y(n2217) );
  clknd2d1_hd U592 ( .A(n2216), .B(n2213), .Y(n2209) );
  clknd2d1_hd U593 ( .A(a_e[5]), .B(n2115), .Y(n2114) );
  clknd2d1_hd U594 ( .A(n2122), .B(a[28]), .Y(n2116) );
  clknd2d1_hd U595 ( .A(b_e[4]), .B(n2205), .Y(n2197) );
  clknd2d1_hd U596 ( .A(n2206), .B(b[26]), .Y(n2201) );
  clknd2d1_hd U597 ( .A(n1579), .B(n2170), .Y(n2175) );
  clknd2d1_hd U598 ( .A(n2203), .B(n2202), .Y(n495) );
  clknd2d1_hd U599 ( .A(a[30]), .B(n2103), .Y(n2108) );
  clknd2d1_hd U600 ( .A(n2184), .B(n2177), .Y(n2179) );
  clknd2d1_hd U601 ( .A(n1959), .B(n1940), .Y(n1942) );
  clknd2d1_hd U602 ( .A(n1996), .B(n1995), .Y(n428) );
  clknd2d1_hd U603 ( .A(DP_OP_154J2_137_6175_n2), .B(n1994), .Y(n1992) );
  clknd2d1_hd U604 ( .A(n1973), .B(n1805), .Y(n265) );
  clknd2d1_hd U605 ( .A(n1808), .B(n1807), .Y(n393) );
  clknd2d1_hd U606 ( .A(n1789), .B(n1741), .Y(n362) );
  clknd2d1_hd U607 ( .A(n2139), .B(n2136), .Y(n2145) );
  clknd2d1_hd U608 ( .A(n2139), .B(n2121), .Y(n2128) );
  clknd2d1_hd U609 ( .A(n2205), .B(n2204), .Y(n2212) );
  clknd2d1_hd U610 ( .A(n2116), .B(n2109), .Y(n2110) );
  ivd4_hd U611 ( .A(n1656), .Y(n1568) );
  ivd3_hd U612 ( .A(n2272), .Y(n1569) );
  oa22d2_hd U613 ( .A(n1657), .B(n1709), .C(a_s), .D(b_s), .Y(n1791) );
  xo2d1_hd U614 ( .A(n2271), .B(DP_OP_43J2_124_6938_n1), .Y(N337) );
  ad2d4_hd U615 ( .A(n2271), .B(n1626), .Y(n1656) );
  oa21d1_hd U616 ( .A(n1623), .B(n1622), .C(n1621), .Y(n1624) );
  ao21d1_hd U617 ( .A(a_m[23]), .B(n2000), .C(n1620), .Y(n1623) );
  nid1_hd U618 ( .A(n1802), .Y(n1571) );
  nid6_hd U619 ( .A(n27), .Y(n1570) );
  ivd2_hd U620 ( .A(n1791), .Y(n2271) );
  ad3d1_hd U621 ( .A(n2223), .B(i_AB_STB), .C(o_AB_ACK), .Y(n27) );
  or2d2_hd U622 ( .A(n1707), .B(n2228), .Y(n2268) );
  ivd1_hd U623 ( .A(b_m[23]), .Y(n2000) );
  nr2d4_hd U624 ( .A(n1656), .B(n1791), .Y(n1654) );
  scg9d1_hd U625 ( .A(n2241), .B(n1701), .C(n2268), .Y(n2161) );
  ad3d1_hd U626 ( .A(n2261), .B(n1576), .C(n2259), .Y(n2265) );
  scg2d1_hd U627 ( .A(b_e[9]), .B(n1698), .C(n1697), .D(n1696), .Y(n1699) );
  ivd2_hd U628 ( .A(n1779), .Y(n1804) );
  ivd2_hd U629 ( .A(n1972), .Y(n1946) );
  or4d1_hd U630 ( .A(z_m[23]), .B(z_e[0]), .C(n1728), .D(n1727), .Y(n1735) );
  or4d1_hd U631 ( .A(n1678), .B(a_e[9]), .C(a_e[0]), .D(a_e[8]), .Y(n1792) );
  or2d1_hd U632 ( .A(n2246), .B(n2247), .Y(n2272) );
  ivd1_hd U633 ( .A(b_m[2]), .Y(n2042) );
  ivd1_hd U634 ( .A(b_m[1]), .Y(n2043) );
  or2d1_hd U635 ( .A(b_e[2]), .B(a_e[2]), .Y(n1771) );
  nr2d2_hd U636 ( .A(n1797), .B(n2227), .Y(n1803) );
  ivd2_hd U637 ( .A(n1952), .Y(n1959) );
  nr2ad1_hd U638 ( .A(n1976), .B(n1989), .Y(n1993) );
  nr2ad1_hd U639 ( .A(n2259), .B(n1935), .Y(n1941) );
  nr2ad1_hd U640 ( .A(n2225), .B(n2247), .Y(n2269) );
  ivd1_hd U641 ( .A(b_m[0]), .Y(n2044) );
  oa22ad1_hd U642 ( .A(n1589), .B(a_m[6]), .C(n1588), .D(b_m[6]), .Y(n1590) );
  ivd1_hd U643 ( .A(b_m[3]), .Y(n2041) );
  ivd1_hd U644 ( .A(b_m[4]), .Y(n2038) );
  ao22d1_hd U645 ( .A(a_m[26]), .B(n2253), .C(n1625), .D(n1624), .Y(n1626) );
  ivd1_hd U646 ( .A(a_m[3]), .Y(n2089) );
  ivd1_hd U647 ( .A(a_m[5]), .Y(n2084) );
  ivd1_hd U648 ( .A(b_m[5]), .Y(n2036) );
  nid2_hd U649 ( .A(n2260), .Y(n1576) );
  ivd1_hd U650 ( .A(n1958), .Y(n1934) );
  ivd1_hd U651 ( .A(n1987), .Y(n1989) );
  ivd1_hd U652 ( .A(n2096), .Y(n1574) );
  oa21d1_hd U653 ( .A(a_m[21]), .B(n2004), .C(n1617), .Y(n1618) );
  ivd1_hd U654 ( .A(a_m[4]), .Y(n2086) );
  ivd1_hd U655 ( .A(n1787), .Y(n1800) );
  ivd1_hd U656 ( .A(n2268), .Y(n1577) );
  nr2d1_hd U657 ( .A(n2261), .B(n1935), .Y(n1958) );
  ivd1_hd U658 ( .A(n1974), .Y(n2261) );
  nid2_hd U659 ( .A(n1947), .Y(n1572) );
  ivd1_hd U660 ( .A(n1941), .Y(n1948) );
  nr2d1_hd U661 ( .A(n2224), .B(n2246), .Y(n1974) );
  ivd1_hd U662 ( .A(n2269), .Y(n1991) );
  ivd2_hd U663 ( .A(n2161), .Y(n1575) );
  ivd2_hd U664 ( .A(n1574), .Y(n1573) );
  ivd1_hd U665 ( .A(n2270), .Y(n2226) );
  ivd1_hd U666 ( .A(n2241), .Y(n2189) );
  nd2bd1_hd U667 ( .AN(n1707), .B(n2237), .Y(n2241) );
  ivd1_hd U668 ( .A(b_m[24]), .Y(n1998) );
  ivd1_hd U669 ( .A(a_m[16]), .Y(n2062) );
  ivd1_hd U670 ( .A(b_m[10]), .Y(n2026) );
  ivd1_hd U671 ( .A(b_m[13]), .Y(n2020) );
  ivd1_hd U672 ( .A(a_m[15]), .Y(n2064) );
  ivd1_hd U673 ( .A(b_m[14]), .Y(n2018) );
  ivd1_hd U674 ( .A(a_m[17]), .Y(n2060) );
  ivd1_hd U675 ( .A(b_m[17]), .Y(n2012) );
  ivd1_hd U676 ( .A(b_m[21]), .Y(n2004) );
  nid2_hd U677 ( .A(n509), .Y(n1580) );
  nr3d1_hd U678 ( .A(n1751), .B(n1717), .C(n1716), .Y(n1802) );
  ivd1_hd U679 ( .A(n1715), .Y(n1751) );
  ivd2_hd U680 ( .A(n2252), .Y(n2039) );
  scg20d2_hd U681 ( .A(n1812), .B(n1966), .C(n265), .Y(n1935) );
  ivd1_hd U682 ( .A(n1975), .Y(n1805) );
  ivd2_hd U683 ( .A(n2268), .Y(n1578) );
  ivd2_hd U684 ( .A(n2094), .Y(n2087) );
  nr2d1_hd U685 ( .A(n2228), .B(n2247), .Y(n1975) );
  nd2bd1_hd U686 ( .AN(n2247), .B(n2237), .Y(n2259) );
  ivd1_hd U687 ( .A(n2205), .Y(n2255) );
  nr2d1_hd U688 ( .A(n2221), .B(n2241), .Y(n2205) );
  ao21d1_hd U689 ( .A(n2163), .B(n2162), .C(n1575), .Y(n2221) );
  ivd1_hd U690 ( .A(n2268), .Y(n1579) );
  ivd1_hd U691 ( .A(n2139), .Y(n2157) );
  nr2d1_hd U692 ( .A(n2154), .B(n2241), .Y(n2139) );
  ao21d1_hd U693 ( .A(n2097), .B(n2162), .C(n1573), .Y(n2154) );
  scg16d1_hd U694 ( .A(n2236), .B(n2235), .C(n2268), .Y(n2096) );
  ivd1_hd U695 ( .A(b_e[1]), .Y(n2215) );
  nr2d1_hd U696 ( .A(n1719), .B(n1716), .Y(n2162) );
  nr2d1_hd U697 ( .A(n1707), .B(n2225), .Y(n2270) );
  ivd1_hd U698 ( .A(b_e[6]), .Y(n2167) );
  ivd1_hd U699 ( .A(a_e[8]), .Y(n2102) );
  ivd1_hd U700 ( .A(a_e[5]), .Y(n2119) );
  ivd1_hd U701 ( .A(a_e[6]), .Y(n2100) );
  nr2d1_hd U702 ( .A(n2249), .B(n2243), .Y(n2237) );
  ivd1_hd U703 ( .A(state[0]), .Y(n2249) );
  ivd1_hd U704 ( .A(state[1]), .Y(n2243) );
  ivd1_hd U705 ( .A(state[3]), .Y(n2263) );
  ivd1_hd U706 ( .A(b_m[25]), .Y(n1628) );
  ivd1_hd U707 ( .A(b_m[19]), .Y(n2008) );
  ivd1_hd U708 ( .A(b_m[20]), .Y(n2006) );
  ivd1_hd U709 ( .A(a_m[20]), .Y(n2054) );
  ivd1_hd U710 ( .A(b_m[22]), .Y(n2002) );
  ivd1_hd U711 ( .A(a_m[22]), .Y(n2050) );
  ivd1_hd U712 ( .A(a_m[25]), .Y(n1668) );
  ivd1_hd U713 ( .A(b_m[26]), .Y(n2253) );
  ivd1_hd U714 ( .A(n2162), .Y(n2245) );
  nr2d1_hd U715 ( .A(n2225), .B(n2224), .Y(n509) );
  ivd1_hd U716 ( .A(n1796), .Y(n2227) );
  ivd1_hd U717 ( .A(z_m[1]), .Y(n1949) );
  ao21d1_hd U718 ( .A(n1796), .B(n1797), .C(n1734), .Y(n1789) );
  ivd1_hd U719 ( .A(n1710), .Y(n1793) );
  nr2d1_hd U720 ( .A(n2228), .B(n2224), .Y(n1796) );
  ivd1_hd U721 ( .A(z_m[20]), .Y(n1832) );
  ivd1_hd U722 ( .A(z_m[21]), .Y(n1826) );
  ivd1_hd U723 ( .A(n1935), .Y(n1955) );
  ivd1_hd U724 ( .A(z_m[22]), .Y(n1968) );
  ivd1_hd U725 ( .A(z_m[17]), .Y(n1850) );
  ivd1_hd U726 ( .A(z_m[18]), .Y(n1838) );
  ivd1_hd U727 ( .A(z_m[13]), .Y(n1874) );
  ivd1_hd U728 ( .A(z_m[14]), .Y(n1862) );
  ivd1_hd U729 ( .A(z_m[10]), .Y(n1886) );
  ivd1_hd U730 ( .A(z_m[9]), .Y(n1901) );
  ivd1_hd U731 ( .A(z_m[5]), .Y(n1926) );
  ivd1_hd U732 ( .A(z_m[6]), .Y(n1913) );
  ivd1_hd U733 ( .A(z_m[23]), .Y(n1967) );
  ivd1_hd U734 ( .A(z_e[0]), .Y(n1988) );
  ivd1_hd U735 ( .A(z_e[7]), .Y(n1733) );
  ivd1_hd U736 ( .A(z_e[8]), .Y(n1978) );
  ivd1_hd U737 ( .A(n2257), .Y(n2210) );
  nr2d1_hd U738 ( .A(n2226), .B(n2221), .Y(n2257) );
  ivd1_hd U739 ( .A(b[30]), .Y(n2176) );
  ivd1_hd U740 ( .A(n2159), .Y(n2143) );
  nr2d1_hd U741 ( .A(n2226), .B(n2154), .Y(n2159) );
  ivd1_hd U742 ( .A(a_e[7]), .Y(n2104) );
  ivd1_hd U743 ( .A(a_e[4]), .Y(n2124) );
  ivd1_hd U744 ( .A(a_e[2]), .Y(n2140) );
  ivd1_hd U745 ( .A(b_e[7]), .Y(n2171) );
  nr3d1_hd U746 ( .A(n1676), .B(n1675), .C(n1674), .Y(n1712) );
  ivd1_hd U747 ( .A(b_e[9]), .Y(n1683) );
  ivd1_hd U748 ( .A(b_e[0]), .Y(n2214) );
  ivd1_hd U749 ( .A(b_e[5]), .Y(n2187) );
  ivd1_hd U750 ( .A(b_e[8]), .Y(n2169) );
  ivd1_hd U751 ( .A(a_e[0]), .Y(n2147) );
  ivd1_hd U752 ( .A(a_e[1]), .Y(n2148) );
  ivd1_hd U753 ( .A(a_e[3]), .Y(n2131) );
  ivd1_hd U754 ( .A(state[2]), .Y(n1718) );
  ivd1_hd U755 ( .A(a_m[1]), .Y(n2091) );
  ivd1_hd U756 ( .A(a_m[2]), .Y(n2090) );
  ivd1_hd U757 ( .A(a_m[6]), .Y(n2082) );
  ivd1_hd U758 ( .A(b_m[6]), .Y(n2034) );
  ivd1_hd U759 ( .A(a_m[7]), .Y(n2080) );
  ivd1_hd U760 ( .A(b_m[7]), .Y(n2032) );
  ivd1_hd U761 ( .A(a_m[11]), .Y(n2072) );
  ivd1_hd U762 ( .A(b_m[11]), .Y(n2024) );
  ivd1_hd U763 ( .A(a_m[13]), .Y(n2068) );
  ivd1_hd U764 ( .A(a_m[14]), .Y(n2066) );
  ivd1_hd U765 ( .A(a_m[18]), .Y(n2058) );
  ivd1_hd U766 ( .A(b_m[18]), .Y(n2010) );
  ivd1_hd U767 ( .A(a_m[21]), .Y(n2052) );
  ivd1_hd U768 ( .A(a_m[23]), .Y(n2048) );
  ivd1_hd U769 ( .A(a_m[24]), .Y(n2046) );
  ivd1_hd U770 ( .A(a_m[19]), .Y(n2056) );
  ivd1_hd U771 ( .A(b_m[15]), .Y(n2016) );
  ivd1_hd U772 ( .A(b_m[16]), .Y(n2014) );
  ivd1_hd U773 ( .A(a_m[12]), .Y(n2070) );
  ivd1_hd U774 ( .A(a_m[8]), .Y(n2078) );
  ivd1_hd U775 ( .A(b_m[8]), .Y(n2030) );
  ivd1_hd U776 ( .A(b_m[9]), .Y(n2028) );
  ivd1_hd U777 ( .A(a_m[10]), .Y(n2074) );
  ivd1_hd U778 ( .A(a_m[9]), .Y(n2076) );
  ivd1_hd U779 ( .A(b_m[12]), .Y(n2022) );
  ivd1_hd U780 ( .A(a_m[26]), .Y(n2095) );
  ivd1_hd U781 ( .A(a_s), .Y(n1709) );
  ivd1_hd U782 ( .A(b_s), .Y(n1657) );
  ivd1_hd U783 ( .A(z_m[0]), .Y(n1956) );
  nr2d1_hd U784 ( .A(n1576), .B(n2226), .Y(n1787) );
  nd2bd1_hd U785 ( .AN(a[30]), .B(n2111), .Y(n2158) );
  ivd1_hd U786 ( .A(a_e[9]), .Y(n1698) );
  nr2d1_hd U787 ( .A(sum[27]), .B(n1805), .Y(n1947) );
  ao22d1_hd U788 ( .A(b_m[25]), .B(n1668), .C(b_m[26]), .D(n2095), .Y(n1625)
         );
  ao22d1_hd U789 ( .A(a_m[21]), .B(n2004), .C(a_m[22]), .D(n2002), .Y(n1619)
         );
  ao22d1_hd U790 ( .A(a_m[20]), .B(n2006), .C(a_m[19]), .D(n2008), .Y(n1616)
         );
  nr2d1_hd U791 ( .A(b_m[15]), .B(n2064), .Y(n1606) );
  ao22d1_hd U792 ( .A(a_m[13]), .B(n2020), .C(a_m[12]), .D(n2022), .Y(n1604)
         );
  ao22d1_hd U793 ( .A(b_m[9]), .B(n2076), .C(b_m[10]), .D(n2074), .Y(n1597) );
  ao22d1_hd U794 ( .A(a_m[9]), .B(n2028), .C(a_m[8]), .D(n2030), .Y(n1595) );
  ao211d1_hd U795 ( .A(a_m[1]), .B(n2043), .C(a_m[0]), .D(n2044), .Y(n1582) );
  oa22d1_hd U796 ( .A(a_m[1]), .B(n2043), .C(a_m[2]), .D(n2042), .Y(n1581) );
  oa22d1_hd U797 ( .A(b_m[3]), .B(n2089), .C(n1582), .D(n1581), .Y(n1583) );
  ao21d1_hd U798 ( .A(a_m[2]), .B(n2042), .C(n1583), .Y(n1585) );
  oa22d1_hd U799 ( .A(a_m[4]), .B(n2038), .C(a_m[3]), .D(n2041), .Y(n1584) );
  oa22d1_hd U800 ( .A(n1585), .B(n1584), .C(b_m[4]), .D(n2086), .Y(n1586) );
  ao22d1_hd U801 ( .A(a_m[5]), .B(n2036), .C(n1587), .D(n1586), .Y(n1588) );
  nr2d1_hd U802 ( .A(n1588), .B(b_m[6]), .Y(n1589) );
  nr2d1_hd U803 ( .A(n1590), .B(b_m[7]), .Y(n1593) );
  oa211d1_hd U804 ( .A(a_m[7]), .B(n1593), .C(n1592), .D(n1591), .Y(n1594) );
  ao22d1_hd U805 ( .A(a_m[10]), .B(n2026), .C(n1597), .D(n1596), .Y(n1598) );
  nr2d1_hd U806 ( .A(b_m[11]), .B(n1598), .Y(n1601) );
  oa211d1_hd U807 ( .A(a_m[11]), .B(n1601), .C(n1600), .D(n1599), .Y(n1603) );
  oa22d1_hd U808 ( .A(a_m[13]), .B(n2020), .C(a_m[14]), .D(n2018), .Y(n1602)
         );
  ao21d1_hd U809 ( .A(n1604), .B(n1603), .C(n1602), .Y(n1605) );
  ao211d1_hd U810 ( .A(a_m[14]), .B(n2018), .C(n1606), .D(n1605), .Y(n1608) );
  oa22d1_hd U811 ( .A(a_m[16]), .B(n2014), .C(a_m[15]), .D(n2016), .Y(n1607)
         );
  oa22d1_hd U812 ( .A(n1608), .B(n1607), .C(b_m[16]), .D(n2062), .Y(n1609) );
  ao22d1_hd U813 ( .A(a_m[17]), .B(n2012), .C(n1610), .D(n1609), .Y(n1611) );
  nr2d1_hd U814 ( .A(b_m[18]), .B(n1611), .Y(n1614) );
  oa211d1_hd U815 ( .A(a_m[18]), .B(n1614), .C(n1613), .D(n1612), .Y(n1615) );
  ao22d1_hd U816 ( .A(b_m[20]), .B(n2054), .C(n1616), .D(n1615), .Y(n1617) );
  ao22d1_hd U817 ( .A(b_m[22]), .B(n2050), .C(n1619), .D(n1618), .Y(n1620) );
  oa22d1_hd U818 ( .A(a_m[23]), .B(n2000), .C(a_m[24]), .D(n1998), .Y(n1622)
         );
  ao22d1_hd U819 ( .A(a_m[24]), .B(n1998), .C(a_m[25]), .D(n1628), .Y(n1621)
         );
  ivd1_hd U820 ( .A(a_m[0]), .Y(n2092) );
  ao22d1_hd U821 ( .A(n1656), .B(n2044), .C(n2092), .D(n1568), .Y(C2_Z_0) );
  ao22d1_hd U822 ( .A(n1656), .B(n2043), .C(n2091), .D(n1568), .Y(C2_Z_1) );
  ao22d1_hd U823 ( .A(n1656), .B(n2026), .C(n2074), .D(n1568), .Y(C2_Z_10) );
  ao22d1_hd U824 ( .A(n1656), .B(n2024), .C(n2072), .D(n1568), .Y(C2_Z_11) );
  ao22d1_hd U825 ( .A(n1656), .B(n2022), .C(n2070), .D(n1568), .Y(C2_Z_12) );
  ao22d1_hd U826 ( .A(n1656), .B(n2020), .C(n2068), .D(n1568), .Y(C2_Z_13) );
  ao22d1_hd U827 ( .A(n1656), .B(n2018), .C(n2066), .D(n1568), .Y(C2_Z_14) );
  ao22d1_hd U828 ( .A(n1656), .B(n2016), .C(n2064), .D(n1568), .Y(C2_Z_15) );
  ao22d1_hd U829 ( .A(n1656), .B(n2014), .C(n2062), .D(n1568), .Y(C2_Z_16) );
  ao22d1_hd U830 ( .A(n1656), .B(n2012), .C(n2060), .D(n1568), .Y(C2_Z_17) );
  ao22d1_hd U831 ( .A(n1656), .B(n2010), .C(n2058), .D(n1568), .Y(C2_Z_18) );
  ao22d1_hd U832 ( .A(n1656), .B(n2008), .C(n2056), .D(n1568), .Y(C2_Z_19) );
  ao22d1_hd U833 ( .A(n1656), .B(n2042), .C(n2090), .D(n1568), .Y(C2_Z_2) );
  ao22d1_hd U834 ( .A(n1656), .B(n2006), .C(n2054), .D(n1568), .Y(C2_Z_20) );
  ao22d1_hd U835 ( .A(n1656), .B(n2004), .C(n2052), .D(n1568), .Y(C2_Z_21) );
  ao22d1_hd U836 ( .A(n1656), .B(n2002), .C(n2050), .D(n1568), .Y(C2_Z_22) );
  ao22d1_hd U837 ( .A(n1656), .B(n2000), .C(n2048), .D(n1568), .Y(C2_Z_23) );
  ao22d1_hd U838 ( .A(n1656), .B(n1998), .C(n2046), .D(n1568), .Y(C2_Z_24) );
  ao22d1_hd U839 ( .A(n1656), .B(n1628), .C(n1668), .D(n1568), .Y(C2_Z_25) );
  oa21d1_hd U840 ( .A(n2253), .B(n1791), .C(n2095), .Y(C2_Z_26) );
  ao22d1_hd U841 ( .A(n1656), .B(n2041), .C(n2089), .D(n1568), .Y(C2_Z_3) );
  ao22d1_hd U842 ( .A(n1656), .B(n2038), .C(n2086), .D(n1568), .Y(C2_Z_4) );
  ao22d1_hd U843 ( .A(n1656), .B(n2036), .C(n2084), .D(n1568), .Y(C2_Z_5) );
  ao22d1_hd U844 ( .A(n1656), .B(n2034), .C(n2082), .D(n1568), .Y(C2_Z_6) );
  ao22d1_hd U845 ( .A(n1656), .B(n2032), .C(n2080), .D(n1568), .Y(C2_Z_7) );
  ao22d1_hd U846 ( .A(n1656), .B(n2030), .C(n2078), .D(n1568), .Y(C2_Z_8) );
  ao22d1_hd U847 ( .A(n1656), .B(n2028), .C(n2076), .D(n1568), .Y(C2_Z_9) );
  nr2d1_hd U848 ( .A(n2253), .B(n2095), .Y(n1627) );
  ao22d1_hd U849 ( .A(n2271), .B(n1627), .C(n2253), .D(n1791), .Y(
        DP_OP_43J2_124_6938_n32) );
  ao22d1_hd U850 ( .A(b_m[25]), .B(n1791), .C(n1654), .D(n1628), .Y(n1629) );
  oa21d1_hd U851 ( .A(a_m[25]), .B(n1568), .C(n1629), .Y(
        DP_OP_43J2_124_6938_n33) );
  ao22d1_hd U852 ( .A(b_m[24]), .B(n1791), .C(n1654), .D(n1998), .Y(n1630) );
  oa21d1_hd U853 ( .A(a_m[24]), .B(n1568), .C(n1630), .Y(
        DP_OP_43J2_124_6938_n34) );
  ao22d1_hd U854 ( .A(b_m[23]), .B(n1791), .C(n1654), .D(n2000), .Y(n1631) );
  oa21d1_hd U855 ( .A(a_m[23]), .B(n1568), .C(n1631), .Y(
        DP_OP_43J2_124_6938_n35) );
  ao22d1_hd U856 ( .A(n1656), .B(n2050), .C(n1654), .D(n2002), .Y(n1632) );
  oa21d1_hd U857 ( .A(n2271), .B(n2002), .C(n1632), .Y(DP_OP_43J2_124_6938_n36) );
  ao22d1_hd U858 ( .A(b_m[21]), .B(n1791), .C(n1654), .D(n2004), .Y(n1633) );
  oa21d1_hd U859 ( .A(a_m[21]), .B(n1568), .C(n1633), .Y(
        DP_OP_43J2_124_6938_n37) );
  ao22d1_hd U860 ( .A(n1656), .B(n2054), .C(n1654), .D(n2006), .Y(n1634) );
  oa21d1_hd U861 ( .A(n2271), .B(n2006), .C(n1634), .Y(DP_OP_43J2_124_6938_n38) );
  ao22d1_hd U862 ( .A(n1656), .B(n2056), .C(n1654), .D(n2008), .Y(n1635) );
  oa21d1_hd U863 ( .A(n2271), .B(n2008), .C(n1635), .Y(DP_OP_43J2_124_6938_n39) );
  ao22d1_hd U864 ( .A(b_m[18]), .B(n1791), .C(n1654), .D(n2010), .Y(n1636) );
  oa21d1_hd U865 ( .A(a_m[18]), .B(n1568), .C(n1636), .Y(
        DP_OP_43J2_124_6938_n40) );
  ao22d1_hd U866 ( .A(n1656), .B(n2060), .C(n1654), .D(n2012), .Y(n1637) );
  oa21d1_hd U867 ( .A(n2271), .B(n2012), .C(n1637), .Y(DP_OP_43J2_124_6938_n41) );
  ao22d1_hd U868 ( .A(n1656), .B(n2062), .C(n1654), .D(n2014), .Y(n1638) );
  oa21d1_hd U869 ( .A(n2271), .B(n2014), .C(n1638), .Y(DP_OP_43J2_124_6938_n42) );
  ao22d1_hd U870 ( .A(n1656), .B(n2064), .C(n1654), .D(n2016), .Y(n1639) );
  oa21d1_hd U871 ( .A(n2271), .B(n2016), .C(n1639), .Y(DP_OP_43J2_124_6938_n43) );
  ao22d1_hd U872 ( .A(b_m[14]), .B(n1791), .C(n1654), .D(n2018), .Y(n1640) );
  oa21d1_hd U873 ( .A(a_m[14]), .B(n1568), .C(n1640), .Y(
        DP_OP_43J2_124_6938_n44) );
  ao22d1_hd U874 ( .A(b_m[13]), .B(n1791), .C(n1654), .D(n2020), .Y(n1641) );
  oa21d1_hd U875 ( .A(a_m[13]), .B(n1568), .C(n1641), .Y(
        DP_OP_43J2_124_6938_n45) );
  ao22d1_hd U876 ( .A(n1656), .B(n2070), .C(n1654), .D(n2022), .Y(n1642) );
  oa21d1_hd U877 ( .A(n2271), .B(n2022), .C(n1642), .Y(DP_OP_43J2_124_6938_n46) );
  ao22d1_hd U878 ( .A(b_m[11]), .B(n1791), .C(n1654), .D(n2024), .Y(n1643) );
  oa21d1_hd U879 ( .A(a_m[11]), .B(n1568), .C(n1643), .Y(
        DP_OP_43J2_124_6938_n47) );
  ao22d1_hd U880 ( .A(n1656), .B(n2074), .C(n1654), .D(n2026), .Y(n1644) );
  oa21d1_hd U881 ( .A(n2271), .B(n2026), .C(n1644), .Y(DP_OP_43J2_124_6938_n48) );
  ao22d1_hd U882 ( .A(n1656), .B(n2076), .C(n1654), .D(n2028), .Y(n1645) );
  oa21d1_hd U883 ( .A(n2271), .B(n2028), .C(n1645), .Y(DP_OP_43J2_124_6938_n49) );
  ao22d1_hd U884 ( .A(n1656), .B(n2078), .C(n1654), .D(n2030), .Y(n1646) );
  oa21d1_hd U885 ( .A(n2271), .B(n2030), .C(n1646), .Y(DP_OP_43J2_124_6938_n50) );
  ao22d1_hd U886 ( .A(b_m[7]), .B(n1791), .C(n1654), .D(n2032), .Y(n1647) );
  oa21d1_hd U887 ( .A(a_m[7]), .B(n1568), .C(n1647), .Y(
        DP_OP_43J2_124_6938_n51) );
  ao22d1_hd U888 ( .A(b_m[6]), .B(n1791), .C(n1654), .D(n2034), .Y(n1648) );
  oa21d1_hd U889 ( .A(a_m[6]), .B(n1568), .C(n1648), .Y(
        DP_OP_43J2_124_6938_n52) );
  ao22d1_hd U890 ( .A(n1656), .B(n2084), .C(n1654), .D(n2036), .Y(n1649) );
  oa21d1_hd U891 ( .A(n2271), .B(n2036), .C(n1649), .Y(DP_OP_43J2_124_6938_n53) );
  ao22d1_hd U892 ( .A(n1656), .B(n2086), .C(n1654), .D(n2038), .Y(n1650) );
  oa21d1_hd U893 ( .A(n2271), .B(n2038), .C(n1650), .Y(DP_OP_43J2_124_6938_n54) );
  ao22d1_hd U894 ( .A(n1656), .B(n2089), .C(n1654), .D(n2041), .Y(n1651) );
  oa21d1_hd U895 ( .A(n2271), .B(n2041), .C(n1651), .Y(DP_OP_43J2_124_6938_n55) );
  ao22d1_hd U896 ( .A(b_m[2]), .B(n1791), .C(n1654), .D(n2042), .Y(n1652) );
  oa21d1_hd U897 ( .A(a_m[2]), .B(n1568), .C(n1652), .Y(
        DP_OP_43J2_124_6938_n56) );
  ao22d1_hd U898 ( .A(b_m[1]), .B(n1791), .C(n1654), .D(n2043), .Y(n1653) );
  oa21d1_hd U899 ( .A(a_m[1]), .B(n1568), .C(n1653), .Y(
        DP_OP_43J2_124_6938_n57) );
  ao22d1_hd U900 ( .A(b_m[0]), .B(n1791), .C(n1654), .D(n2044), .Y(n1655) );
  oa21d1_hd U901 ( .A(a_m[0]), .B(n1568), .C(n1655), .Y(
        DP_OP_43J2_124_6938_n58) );
  ao22d1_hd U902 ( .A(n1656), .B(n1657), .C(n1709), .D(n1568), .Y(N338) );
  nr4d1_hd U903 ( .A(a_e[1]), .B(a_e[2]), .C(a_e[3]), .D(a_e[4]), .Y(n1658) );
  nd4d1_hd U904 ( .A(a_e[7]), .B(n1658), .C(n2100), .D(n2119), .Y(n1678) );
  nr4d1_hd U905 ( .A(n1678), .B(n2147), .C(n1698), .D(n2102), .Y(n2097) );
  nr4d1_hd U906 ( .A(b_e[2]), .B(b_e[1]), .C(b_e[3]), .D(b_e[4]), .Y(n1659) );
  nd4d1_hd U907 ( .A(b_e[7]), .B(n1659), .C(n2187), .D(n2167), .Y(n1677) );
  nr4d1_hd U908 ( .A(n2169), .B(n1677), .C(n2214), .D(n1683), .Y(n2163) );
  nd4d1_hd U909 ( .A(n2036), .B(n2038), .C(n2028), .D(n2016), .Y(n1667) );
  nr4d1_hd U910 ( .A(b_m[0]), .B(b_m[1]), .C(b_m[2]), .D(b_m[3]), .Y(n1660) );
  nd4d1_hd U911 ( .A(n1660), .B(n2014), .C(n2034), .D(n2020), .Y(n1666) );
  nr4d1_hd U912 ( .A(b_m[25]), .B(b_m[23]), .C(b_m[22]), .D(b_m[26]), .Y(n1664) );
  nr4d1_hd U913 ( .A(b_m[18]), .B(b_m[11]), .C(b_m[14]), .D(b_m[24]), .Y(n1663) );
  nr4d1_hd U914 ( .A(b_m[8]), .B(b_m[7]), .C(b_m[10]), .D(b_m[12]), .Y(n1662)
         );
  nr4d1_hd U915 ( .A(b_m[17]), .B(b_m[19]), .C(b_m[20]), .D(b_m[21]), .Y(n1661) );
  nd4d1_hd U916 ( .A(n1664), .B(n1663), .C(n1662), .D(n1661), .Y(n1665) );
  nr3d1_hd U917 ( .A(n1667), .B(n1666), .C(n1665), .Y(n1711) );
  nd4d1_hd U918 ( .A(n2060), .B(n2078), .C(n2052), .D(n2046), .Y(n1676) );
  nr4d1_hd U919 ( .A(a_m[18]), .B(a_m[12]), .C(a_m[20]), .D(a_m[26]), .Y(n1669) );
  nd4d1_hd U920 ( .A(n1669), .B(n2048), .C(n2050), .D(n1668), .Y(n1675) );
  nr4d1_hd U921 ( .A(a_m[11]), .B(a_m[6]), .C(a_m[9]), .D(a_m[10]), .Y(n1673)
         );
  nr4d1_hd U922 ( .A(a_m[13]), .B(a_m[14]), .C(a_m[15]), .D(a_m[19]), .Y(n1672) );
  nr4d1_hd U923 ( .A(a_m[16]), .B(a_m[5]), .C(a_m[4]), .D(a_m[7]), .Y(n1671)
         );
  nr4d1_hd U924 ( .A(a_m[0]), .B(a_m[1]), .C(a_m[2]), .D(a_m[3]), .Y(n1670) );
  nd4d1_hd U925 ( .A(n1673), .B(n1672), .C(n1671), .D(n1670), .Y(n1674) );
  nr4d1_hd U926 ( .A(b_e[8]), .B(b_e[0]), .C(b_e[9]), .D(n1677), .Y(n1710) );
  nr2d1_hd U927 ( .A(n1710), .B(n2226), .Y(n1750) );
  ao22d1_hd U928 ( .A(b_e[2]), .B(n2140), .C(b_e[3]), .D(n2131), .Y(n1685) );
  nr2d1_hd U929 ( .A(a_e[1]), .B(n2215), .Y(n1681) );
  ao22d1_hd U930 ( .A(b_e[4]), .B(n2124), .C(b_e[5]), .D(n2119), .Y(n1680) );
  ao211d1_hd U931 ( .A(b_e[0]), .B(n2147), .C(n1681), .D(n1688), .Y(n1682) );
  oa211d1_hd U932 ( .A(a_e[7]), .B(n2171), .C(n1685), .D(n1682), .Y(n1684) );
  nd3bd1_hd U933 ( .AN(n1684), .B(n1697), .C(n1700), .Y(n2236) );
  ao211d1_hd U934 ( .A(b_e[6]), .B(n2100), .C(b_e[5]), .D(n2119), .Y(n1692) );
  ivd1_hd U935 ( .A(b_e[4]), .Y(n2193) );
  ivd1_hd U936 ( .A(b_e[3]), .Y(n2164) );
  ao22d1_hd U937 ( .A(a_e[4]), .B(n2193), .C(a_e[3]), .D(n2164), .Y(n1690) );
  ao211d1_hd U938 ( .A(b_e[1]), .B(n2148), .C(b_e[0]), .D(n2147), .Y(n1687) );
  oa22d1_hd U939 ( .A(b_e[1]), .B(n2148), .C(b_e[2]), .D(n2140), .Y(n1686) );
  oa21d1_hd U940 ( .A(n1687), .B(n1686), .C(n1685), .Y(n1689) );
  ao21d1_hd U941 ( .A(n1690), .B(n1689), .C(n1688), .Y(n1691) );
  ao211d1_hd U942 ( .A(a_e[6]), .B(n2167), .C(n1692), .D(n1691), .Y(n1695) );
  scg6d1_hd U943 ( .A(b_e[7]), .B(n1695), .C(n2104), .Y(n1693) );
  oa211d1_hd U944 ( .A(b_e[7]), .B(n1695), .C(n1694), .D(n1693), .Y(n1696) );
  oa21d1_hd U945 ( .A(n2097), .B(n2245), .C(n1574), .Y(n1) );
  oa21d1_hd U946 ( .A(n2163), .B(n2245), .C(n2161), .Y(n2) );
  nr2d1_hd U947 ( .A(n1733), .B(n1978), .Y(n1703) );
  nr4d1_hd U948 ( .A(z_e[2]), .B(z_e[3]), .C(z_e[4]), .D(z_e[5]), .Y(n1702) );
  ivd1_hd U949 ( .A(z_e[6]), .Y(n1745) );
  nd3d1_hd U950 ( .A(z_e[9]), .B(n1702), .C(n1745), .Y(n1728) );
  ivd1_hd U951 ( .A(z_e[9]), .Y(n1990) );
  ao21d1_hd U952 ( .A(n1703), .B(n1728), .C(n1990), .Y(n1705) );
  nr2d1_hd U953 ( .A(n2259), .B(n2231), .Y(n1806) );
  nr2d1_hd U954 ( .A(n1727), .B(n1988), .Y(n1704) );
  scg16d1_hd U955 ( .A(n1705), .B(n1704), .C(n1967), .Y(n2230) );
  nr2d1_hd U956 ( .A(n2230), .B(n1991), .Y(n1706) );
  nr2d1_hd U957 ( .A(n1806), .B(n1706), .Y(n1973) );
  ivd1_hd U958 ( .A(n2259), .Y(n2232) );
  scg4d1_hd U959 ( .A(n2232), .B(z_m[0]), .C(n2269), .D(round_bit), .E(n1572), 
        .F(sum[2]), .G(sum[3]), .H(n1946), .Y(n266) );
  nr2d1_hd U960 ( .A(n1707), .B(n2246), .Y(n2223) );
  nr2d1_hd U961 ( .A(a_s), .B(n1717), .Y(n1708) );
  oa21d1_hd U962 ( .A(n1715), .B(n1708), .C(n1793), .Y(n1714) );
  nr3d1_hd U963 ( .A(n1710), .B(n1792), .C(n1709), .Y(n1713) );
  oa22d1_hd U964 ( .A(n1712), .B(n1792), .C(n1711), .D(n1793), .Y(n1794) );
  ao211d1_hd U965 ( .A(b_s), .B(n1714), .C(n1713), .D(n1794), .Y(n1732) );
  ao21d1_hd U966 ( .A(n1792), .B(n1793), .C(n2226), .Y(n1734) );
  ao211d1_hd U967 ( .A(n2270), .B(n1719), .C(n1734), .D(n1796), .Y(n2260) );
  ao22d1_hd U968 ( .A(a_s), .B(n1571), .C(n1576), .D(z[31]), .Y(n1731) );
  ivd1_hd U969 ( .A(z_m[4]), .Y(n1919) );
  ivd1_hd U970 ( .A(z_m[3]), .Y(n1927) );
  nd4d1_hd U971 ( .A(n1949), .B(n1919), .C(n1927), .D(n1913), .Y(n1720) );
  nr4d1_hd U972 ( .A(z_m[0]), .B(z_m[19]), .C(z_m[2]), .D(n1720), .Y(n1726) );
  ivd1_hd U973 ( .A(z_m[12]), .Y(n1868) );
  ivd1_hd U974 ( .A(z_m[11]), .Y(n1875) );
  nd4d1_hd U975 ( .A(n1886), .B(n1868), .C(n1875), .D(n1862), .Y(n1724) );
  ivd1_hd U976 ( .A(z_m[8]), .Y(n1892) );
  ivd1_hd U977 ( .A(z_m[7]), .Y(n1902) );
  nd4d1_hd U978 ( .A(n1926), .B(n1892), .C(n1902), .D(n1901), .Y(n1723) );
  nd4d1_hd U979 ( .A(n1968), .B(n1826), .C(n1832), .D(n1850), .Y(n1722) );
  ivd1_hd U980 ( .A(z_m[16]), .Y(n1844) );
  ivd1_hd U981 ( .A(z_m[15]), .Y(n1851) );
  nd4d1_hd U982 ( .A(n1874), .B(n1844), .C(n1851), .D(n1838), .Y(n1721) );
  nr4d1_hd U983 ( .A(n1724), .B(n1723), .C(n1722), .D(n1721), .Y(n1725) );
  oa211d1_hd U984 ( .A(n1729), .B(n1735), .C(n1796), .D(z_s), .Y(n1730) );
  oa211d1_hd U985 ( .A(n1732), .B(n2226), .C(n1731), .D(n1730), .Y(n361) );
  ao21d1_hd U986 ( .A(n1733), .B(n1978), .C(z_e[9]), .Y(n1797) );
  nr2d1_hd U987 ( .A(z_e[1]), .B(z_e[0]), .Y(n1778) );
  ivd1_hd U988 ( .A(z_e[2]), .Y(n1773) );
  nr2d1_hd U989 ( .A(z_e[3]), .B(n1772), .Y(n1764) );
  ivd1_hd U990 ( .A(z_e[4]), .Y(n1760) );
  nr2d1_hd U991 ( .A(z_e[5]), .B(n1759), .Y(n1749) );
  nr2d1_hd U992 ( .A(z_e[7]), .B(n1744), .Y(n1736) );
  ao211d1_hd U993 ( .A(z_e[7]), .B(n1744), .C(n1790), .D(n1736), .Y(n1740) );
  nd3d1_hd U994 ( .A(n2215), .B(n2148), .C(n1786), .Y(n1780) );
  nr2d1_hd U995 ( .A(n1780), .B(n1771), .Y(n1770) );
  nd3d1_hd U996 ( .A(n1770), .B(n2164), .C(n2131), .Y(n1765) );
  nr2d1_hd U997 ( .A(n1765), .B(n1758), .Y(n1757) );
  nd3d1_hd U998 ( .A(n1757), .B(n2187), .C(n2119), .Y(n1752) );
  nr2d1_hd U999 ( .A(n1752), .B(n1743), .Y(n1742) );
  nr2d1_hd U1000 ( .A(n1742), .B(n1738), .Y(n1737) );
  ao211d1_hd U1001 ( .A(n1742), .B(n1738), .C(n1800), .D(n1737), .Y(n1739) );
  ao211d1_hd U1002 ( .A(n1576), .B(z[30]), .C(n1740), .D(n1739), .Y(n1741) );
  ao21d1_hd U1003 ( .A(n1752), .B(n1743), .C(n1742), .Y(n1748) );
  ivd1_hd U1004 ( .A(n1790), .Y(n1775) );
  oa21d1_hd U1005 ( .A(n1749), .B(n1745), .C(n1744), .Y(n1746) );
  ao22d1_hd U1006 ( .A(n1576), .B(z[29]), .C(n1775), .D(n1746), .Y(n1747) );
  oa211d1_hd U1007 ( .A(n1748), .B(n1800), .C(n1789), .D(n1747), .Y(n363) );
  ao21d1_hd U1008 ( .A(z_e[5]), .B(n1759), .C(n1749), .Y(n1756) );
  ao22d1_hd U1009 ( .A(b_e[5]), .B(n1804), .C(a_e[5]), .D(n1787), .Y(n1753) );
  oa22d1_hd U1010 ( .A(n1757), .B(n1753), .C(n1800), .D(n1752), .Y(n1754) );
  ao21d1_hd U1011 ( .A(n1576), .B(z[28]), .C(n1754), .Y(n1755) );
  oa211d1_hd U1012 ( .A(n1756), .B(n1790), .C(n1789), .D(n1755), .Y(n364) );
  ao21d1_hd U1013 ( .A(n1765), .B(n1758), .C(n1757), .Y(n1763) );
  oa21d1_hd U1014 ( .A(n1764), .B(n1760), .C(n1759), .Y(n1761) );
  ao22d1_hd U1015 ( .A(n1576), .B(z[27]), .C(n1775), .D(n1761), .Y(n1762) );
  oa211d1_hd U1016 ( .A(n1763), .B(n1800), .C(n1789), .D(n1762), .Y(n365) );
  ao21d1_hd U1017 ( .A(z_e[3]), .B(n1772), .C(n1764), .Y(n1769) );
  ao22d1_hd U1018 ( .A(b_e[3]), .B(n1804), .C(a_e[3]), .D(n1787), .Y(n1766) );
  oa22d1_hd U1019 ( .A(n1770), .B(n1766), .C(n1800), .D(n1765), .Y(n1767) );
  ao21d1_hd U1020 ( .A(n1576), .B(z[26]), .C(n1767), .Y(n1768) );
  oa211d1_hd U1021 ( .A(n1769), .B(n1790), .C(n1789), .D(n1768), .Y(n366) );
  ao21d1_hd U1022 ( .A(n1780), .B(n1771), .C(n1770), .Y(n1777) );
  oa21d1_hd U1023 ( .A(n1778), .B(n1773), .C(n1772), .Y(n1774) );
  ao22d1_hd U1024 ( .A(n1576), .B(z[25]), .C(n1775), .D(n1774), .Y(n1776) );
  oa211d1_hd U1025 ( .A(n1777), .B(n1800), .C(n1789), .D(n1776), .Y(n367) );
  ao21d1_hd U1026 ( .A(z_e[0]), .B(z_e[1]), .C(n1778), .Y(n1785) );
  nr3d1_hd U1027 ( .A(n2215), .B(n1786), .C(n1779), .Y(n1783) );
  nd2bd1_hd U1028 ( .AN(n1786), .B(a_e[1]), .Y(n1781) );
  ao21d1_hd U1029 ( .A(n1781), .B(n1780), .C(n1800), .Y(n1782) );
  ao211d1_hd U1030 ( .A(n1576), .B(z[24]), .C(n1783), .D(n1782), .Y(n1784) );
  oa211d1_hd U1031 ( .A(n1785), .B(n1790), .C(n1789), .D(n1784), .Y(n368) );
  ao22d1_hd U1032 ( .A(n1576), .B(z[23]), .C(n1787), .D(n1786), .Y(n1788) );
  oa211d1_hd U1033 ( .A(z_e[0]), .B(n1790), .C(n1789), .D(n1788), .Y(n369) );
  nr3d1_hd U1034 ( .A(n1793), .B(n1792), .C(n1791), .Y(n1795) );
  nr2d1_hd U1035 ( .A(n1795), .B(n1794), .Y(n1801) );
  ao22d1_hd U1036 ( .A(b_m[25]), .B(n1804), .C(z_m[22]), .D(n1803), .Y(n1799)
         );
  ao22d1_hd U1037 ( .A(a_m[25]), .B(n1571), .C(n1576), .D(z[22]), .Y(n1798) );
  oa211d1_hd U1038 ( .A(n1801), .B(n1800), .C(n1799), .D(n1798), .Y(n370) );
  scg4d1_hd U1039 ( .A(b_m[24]), .B(n1804), .C(z_m[21]), .D(n1803), .E(a_m[24]), .F(n1571), .G(n1576), .H(z[21]), .Y(n371) );
  scg4d1_hd U1040 ( .A(b_m[23]), .B(n1804), .C(z_m[20]), .D(n1803), .E(a_m[23]), .F(n1571), .G(n1576), .H(z[20]), .Y(n372) );
  scg4d1_hd U1041 ( .A(b_m[22]), .B(n1804), .C(z_m[19]), .D(n1803), .E(a_m[22]), .F(n1571), .G(n1576), .H(z[19]), .Y(n373) );
  scg4d1_hd U1042 ( .A(b_m[21]), .B(n1804), .C(z_m[18]), .D(n1803), .E(a_m[21]), .F(n1571), .G(n1576), .H(z[18]), .Y(n374) );
  scg4d1_hd U1043 ( .A(b_m[20]), .B(n1804), .C(z_m[17]), .D(n1803), .E(a_m[20]), .F(n1571), .G(n1576), .H(z[17]), .Y(n375) );
  scg4d1_hd U1044 ( .A(b_m[19]), .B(n1804), .C(z_m[16]), .D(n1803), .E(a_m[19]), .F(n1571), .G(n1576), .H(z[16]), .Y(n376) );
  scg4d1_hd U1045 ( .A(b_m[18]), .B(n1804), .C(z_m[15]), .D(n1803), .E(a_m[18]), .F(n1571), .G(n1576), .H(z[15]), .Y(n377) );
  scg4d1_hd U1046 ( .A(b_m[17]), .B(n1804), .C(z_m[14]), .D(n1803), .E(a_m[17]), .F(n1571), .G(n1576), .H(z[14]), .Y(n378) );
  scg4d1_hd U1047 ( .A(b_m[16]), .B(n1804), .C(z_m[13]), .D(n1803), .E(a_m[16]), .F(n1571), .G(n1576), .H(z[13]), .Y(n379) );
  scg4d1_hd U1048 ( .A(b_m[15]), .B(n1804), .C(z_m[12]), .D(n1803), .E(a_m[15]), .F(n1571), .G(n1576), .H(z[12]), .Y(n380) );
  scg4d1_hd U1049 ( .A(b_m[14]), .B(n1804), .C(z_m[11]), .D(n1803), .E(a_m[14]), .F(n1802), .G(n1576), .H(z[11]), .Y(n381) );
  scg4d1_hd U1050 ( .A(b_m[13]), .B(n1804), .C(z_m[10]), .D(n1803), .E(a_m[13]), .F(n1802), .G(n1576), .H(z[10]), .Y(n382) );
  scg4d1_hd U1051 ( .A(b_m[12]), .B(n1804), .C(z_m[9]), .D(n1803), .E(a_m[12]), 
        .F(n1802), .G(n1576), .H(z[9]), .Y(n383) );
  scg4d1_hd U1052 ( .A(b_m[11]), .B(n1804), .C(z_m[8]), .D(n1803), .E(a_m[11]), 
        .F(n1802), .G(n1576), .H(z[8]), .Y(n384) );
  scg4d1_hd U1053 ( .A(b_m[10]), .B(n1804), .C(z_m[7]), .D(n1803), .E(a_m[10]), 
        .F(n1802), .G(n1576), .H(z[7]), .Y(n385) );
  scg4d1_hd U1054 ( .A(b_m[9]), .B(n1804), .C(z_m[6]), .D(n1803), .E(a_m[9]), 
        .F(n1802), .G(n1576), .H(z[6]), .Y(n386) );
  scg4d1_hd U1055 ( .A(b_m[8]), .B(n1804), .C(z_m[5]), .D(n1803), .E(a_m[8]), 
        .F(n1571), .G(n1576), .H(z[5]), .Y(n387) );
  scg4d1_hd U1056 ( .A(b_m[7]), .B(n1804), .C(z_m[4]), .D(n1803), .E(a_m[7]), 
        .F(n1571), .G(n2260), .H(z[4]), .Y(n388) );
  scg4d1_hd U1057 ( .A(b_m[6]), .B(n1804), .C(z_m[3]), .D(n1803), .E(a_m[6]), 
        .F(n1571), .G(n1576), .H(z[3]), .Y(n389) );
  scg4d1_hd U1058 ( .A(b_m[5]), .B(n1804), .C(z_m[2]), .D(n1803), .E(a_m[5]), 
        .F(n1571), .G(n1576), .H(z[2]), .Y(n390) );
  scg4d1_hd U1059 ( .A(b_m[4]), .B(n1804), .C(z_m[1]), .D(n1803), .E(a_m[4]), 
        .F(n1571), .G(n1576), .H(z[1]), .Y(n391) );
  scg4d1_hd U1060 ( .A(b_m[3]), .B(n1804), .C(z_m[0]), .D(n1803), .E(a_m[3]), 
        .F(n1802), .G(n1576), .H(z[0]), .Y(n392) );
  ao22d1_hd U1061 ( .A(n1975), .B(sum[0]), .C(sticky), .D(n1805), .Y(n1808) );
  ao22d1_hd U1062 ( .A(n1806), .B(round_bit), .C(n1946), .D(sum[1]), .Y(n1807)
         );
  ivd1_hd U1063 ( .A(round_bit), .Y(n1811) );
  ao22d1_hd U1064 ( .A(n1572), .B(sum[1]), .C(n1946), .D(sum[2]), .Y(n1810) );
  nd3d1_hd U1065 ( .A(n2232), .B(guard), .C(n265), .Y(n1809) );
  oa211d1_hd U1066 ( .A(n1811), .B(n265), .C(n1810), .D(n1809), .Y(n394) );
  nr3d1_hd U1067 ( .A(z_m[0]), .B(sticky), .C(round_bit), .Y(n1812) );
  ao22d1_hd U1068 ( .A(n1572), .B(sum[25]), .C(n1946), .D(sum[26]), .Y(n1816)
         );
  nd3d1_hd U1069 ( .A(z_m[0]), .B(z_m[2]), .C(z_m[1]), .Y(n1920) );
  ivd1_hd U1070 ( .A(n1920), .Y(n1921) );
  nd3d1_hd U1071 ( .A(n1921), .B(z_m[4]), .C(z_m[3]), .Y(n1908) );
  nr3d1_hd U1072 ( .A(n1908), .B(n1913), .C(n1926), .Y(n1893) );
  nd3d1_hd U1073 ( .A(n1893), .B(z_m[8]), .C(z_m[7]), .Y(n1881) );
  nr3d1_hd U1074 ( .A(n1881), .B(n1901), .C(n1886), .Y(n1869) );
  nd3d1_hd U1075 ( .A(n1869), .B(z_m[12]), .C(z_m[11]), .Y(n1857) );
  nr3d1_hd U1076 ( .A(n1857), .B(n1862), .C(n1874), .Y(n1845) );
  nd3d1_hd U1077 ( .A(n1845), .B(z_m[16]), .C(z_m[15]), .Y(n1833) );
  nr3d1_hd U1078 ( .A(n1833), .B(n1838), .C(n1850), .Y(n1970) );
  oa21d1_hd U1079 ( .A(n1970), .B(n2261), .C(n1955), .Y(n1829) );
  ao21d1_hd U1080 ( .A(n1974), .B(n1813), .C(n1829), .Y(n1817) );
  oa21d1_hd U1081 ( .A(z_m[21]), .B(n1934), .C(n1817), .Y(n1957) );
  ivd1_hd U1082 ( .A(z_m[19]), .Y(n1965) );
  nr2d1_hd U1083 ( .A(n1965), .B(n1827), .Y(n1823) );
  oa21d1_hd U1084 ( .A(z_m[22]), .B(n1961), .C(n1959), .Y(n1814) );
  ao22d1_hd U1085 ( .A(z_m[22]), .B(n1957), .C(z_m[21]), .D(n1814), .Y(n1815)
         );
  oa211d1_hd U1086 ( .A(n1967), .B(n1948), .C(n1816), .D(n1815), .Y(n395) );
  ao22d1_hd U1087 ( .A(n1572), .B(sum[24]), .C(sum[25]), .D(n1946), .Y(n1820)
         );
  ao22d1_hd U1088 ( .A(z_m[21]), .B(n1817), .C(n1961), .D(n1826), .Y(n1818) );
  ao21d1_hd U1089 ( .A(z_m[20]), .B(n1952), .C(n1818), .Y(n1819) );
  oa211d1_hd U1090 ( .A(n1968), .B(n1948), .C(n1820), .D(n1819), .Y(n396) );
  ao22d1_hd U1091 ( .A(n1572), .B(sum[23]), .C(n1946), .D(sum[24]), .Y(n1825)
         );
  ao21d1_hd U1092 ( .A(n1958), .B(n1965), .C(n1829), .Y(n1821) );
  oa22d1_hd U1093 ( .A(n1821), .B(n1832), .C(n1965), .D(n1959), .Y(n1822) );
  ao21d1_hd U1094 ( .A(n1823), .B(n1832), .C(n1822), .Y(n1824) );
  oa211d1_hd U1095 ( .A(n1826), .B(n1948), .C(n1825), .D(n1824), .Y(n397) );
  ao22d1_hd U1096 ( .A(n1572), .B(sum[22]), .C(n1946), .D(sum[23]), .Y(n1831)
         );
  oa22d1_hd U1097 ( .A(z_m[19]), .B(n1827), .C(n1959), .D(n1838), .Y(n1828) );
  ao21d1_hd U1098 ( .A(z_m[19]), .B(n1829), .C(n1828), .Y(n1830) );
  oa211d1_hd U1099 ( .A(n1832), .B(n1948), .C(n1831), .D(n1830), .Y(n398) );
  nr2d1_hd U1100 ( .A(n1934), .B(n1833), .Y(n1841) );
  ao21d1_hd U1101 ( .A(n1841), .B(n1838), .C(n1952), .Y(n1837) );
  ao22d1_hd U1102 ( .A(n1572), .B(sum[21]), .C(n1946), .D(sum[22]), .Y(n1836)
         );
  ao21d1_hd U1103 ( .A(n1974), .B(n1833), .C(n1935), .Y(n1839) );
  oa21d1_hd U1104 ( .A(z_m[17]), .B(n1934), .C(n1839), .Y(n1834) );
  ao22d1_hd U1105 ( .A(z_m[19]), .B(n1941), .C(z_m[18]), .D(n1834), .Y(n1835)
         );
  oa211d1_hd U1106 ( .A(n1837), .B(n1850), .C(n1836), .D(n1835), .Y(n399) );
  ao22d1_hd U1107 ( .A(n1572), .B(sum[20]), .C(n1946), .D(sum[21]), .Y(n1843)
         );
  oa22d1_hd U1108 ( .A(n1839), .B(n1850), .C(n1838), .D(n1948), .Y(n1840) );
  ao21d1_hd U1109 ( .A(n1841), .B(n1850), .C(n1840), .Y(n1842) );
  oa211d1_hd U1110 ( .A(n1844), .B(n1959), .C(n1843), .D(n1842), .Y(n400) );
  ao22d1_hd U1111 ( .A(n1572), .B(sum[19]), .C(n1946), .D(sum[20]), .Y(n1849)
         );
  scg20d1_hd U1112 ( .A(n2261), .B(n1845), .C(n1935), .Y(n1853) );
  oa21d1_hd U1113 ( .A(z_m[15]), .B(n1934), .C(n1853), .Y(n1847) );
  oa21d1_hd U1114 ( .A(z_m[16]), .B(n1852), .C(n1959), .Y(n1846) );
  ao22d1_hd U1115 ( .A(z_m[16]), .B(n1847), .C(z_m[15]), .D(n1846), .Y(n1848)
         );
  oa211d1_hd U1116 ( .A(n1850), .B(n1948), .C(n1849), .D(n1848), .Y(n401) );
  ao22d1_hd U1117 ( .A(n1572), .B(sum[18]), .C(n1946), .D(sum[19]), .Y(n1856)
         );
  ao22d1_hd U1118 ( .A(z_m[15]), .B(n1853), .C(n1852), .D(n1851), .Y(n1854) );
  ao21d1_hd U1119 ( .A(z_m[16]), .B(n1941), .C(n1854), .Y(n1855) );
  oa211d1_hd U1120 ( .A(n1862), .B(n1959), .C(n1856), .D(n1855), .Y(n402) );
  nr2d1_hd U1121 ( .A(n1934), .B(n1857), .Y(n1865) );
  ao21d1_hd U1122 ( .A(n1865), .B(n1862), .C(n1952), .Y(n1861) );
  ao22d1_hd U1123 ( .A(n1572), .B(sum[17]), .C(n1946), .D(sum[18]), .Y(n1860)
         );
  ao21d1_hd U1124 ( .A(n1974), .B(n1857), .C(n1935), .Y(n1863) );
  oa21d1_hd U1125 ( .A(z_m[13]), .B(n1934), .C(n1863), .Y(n1858) );
  ao22d1_hd U1126 ( .A(z_m[14]), .B(n1858), .C(z_m[15]), .D(n1941), .Y(n1859)
         );
  oa211d1_hd U1127 ( .A(n1861), .B(n1874), .C(n1860), .D(n1859), .Y(n403) );
  ao22d1_hd U1128 ( .A(n1572), .B(sum[16]), .C(n1946), .D(sum[17]), .Y(n1867)
         );
  oa22d1_hd U1129 ( .A(n1863), .B(n1874), .C(n1862), .D(n1948), .Y(n1864) );
  ao21d1_hd U1130 ( .A(n1865), .B(n1874), .C(n1864), .Y(n1866) );
  oa211d1_hd U1131 ( .A(n1868), .B(n1959), .C(n1867), .D(n1866), .Y(n404) );
  ao22d1_hd U1132 ( .A(n1572), .B(sum[15]), .C(n1946), .D(sum[16]), .Y(n1873)
         );
  scg20d1_hd U1133 ( .A(n2261), .B(n1869), .C(n1935), .Y(n1877) );
  oa21d1_hd U1134 ( .A(z_m[11]), .B(n1934), .C(n1877), .Y(n1871) );
  oa21d1_hd U1135 ( .A(z_m[12]), .B(n1876), .C(n1959), .Y(n1870) );
  ao22d1_hd U1136 ( .A(z_m[12]), .B(n1871), .C(z_m[11]), .D(n1870), .Y(n1872)
         );
  oa211d1_hd U1137 ( .A(n1874), .B(n1948), .C(n1873), .D(n1872), .Y(n405) );
  ao22d1_hd U1138 ( .A(n1572), .B(sum[14]), .C(n1946), .D(sum[15]), .Y(n1880)
         );
  ao22d1_hd U1139 ( .A(z_m[11]), .B(n1877), .C(n1876), .D(n1875), .Y(n1878) );
  ao21d1_hd U1140 ( .A(z_m[12]), .B(n1941), .C(n1878), .Y(n1879) );
  oa211d1_hd U1141 ( .A(n1886), .B(n1959), .C(n1880), .D(n1879), .Y(n406) );
  nr2d1_hd U1142 ( .A(n1934), .B(n1881), .Y(n1889) );
  ao21d1_hd U1143 ( .A(n1889), .B(n1886), .C(n1952), .Y(n1885) );
  ao22d1_hd U1144 ( .A(n1572), .B(sum[13]), .C(n1946), .D(sum[14]), .Y(n1884)
         );
  ao21d1_hd U1145 ( .A(n1974), .B(n1881), .C(n1935), .Y(n1887) );
  oa21d1_hd U1146 ( .A(z_m[9]), .B(n1934), .C(n1887), .Y(n1882) );
  ao22d1_hd U1147 ( .A(z_m[10]), .B(n1882), .C(z_m[11]), .D(n1941), .Y(n1883)
         );
  oa211d1_hd U1148 ( .A(n1885), .B(n1901), .C(n1884), .D(n1883), .Y(n407) );
  ao22d1_hd U1149 ( .A(n1572), .B(sum[12]), .C(n1946), .D(sum[13]), .Y(n1891)
         );
  oa22d1_hd U1150 ( .A(n1887), .B(n1901), .C(n1886), .D(n1948), .Y(n1888) );
  ao21d1_hd U1151 ( .A(n1889), .B(n1901), .C(n1888), .Y(n1890) );
  oa211d1_hd U1152 ( .A(n1892), .B(n1959), .C(n1891), .D(n1890), .Y(n408) );
  ao22d1_hd U1153 ( .A(n1572), .B(sum[11]), .C(n1946), .D(sum[12]), .Y(n1900)
         );
  scg20d1_hd U1154 ( .A(n2261), .B(n1893), .C(n1935), .Y(n1904) );
  oa21d1_hd U1155 ( .A(z_m[7]), .B(n1934), .C(n1904), .Y(n1898) );
  oa21d1_hd U1156 ( .A(z_m[8]), .B(n1903), .C(n1959), .Y(n1894) );
  ao22d1_hd U1157 ( .A(z_m[8]), .B(n1898), .C(z_m[7]), .D(n1894), .Y(n1899) );
  oa211d1_hd U1158 ( .A(n1901), .B(n1948), .C(n1900), .D(n1899), .Y(n409) );
  ao22d1_hd U1159 ( .A(n1572), .B(sum[10]), .C(n1946), .D(sum[11]), .Y(n1907)
         );
  ao22d1_hd U1160 ( .A(z_m[7]), .B(n1904), .C(n1903), .D(n1902), .Y(n1905) );
  ao21d1_hd U1161 ( .A(z_m[8]), .B(n1941), .C(n1905), .Y(n1906) );
  oa211d1_hd U1162 ( .A(n1913), .B(n1959), .C(n1907), .D(n1906), .Y(n410) );
  nr2d1_hd U1163 ( .A(n1934), .B(n1908), .Y(n1916) );
  ao21d1_hd U1164 ( .A(n1916), .B(n1913), .C(n1952), .Y(n1912) );
  ao22d1_hd U1165 ( .A(n1572), .B(sum[9]), .C(n1946), .D(sum[10]), .Y(n1911)
         );
  ao21d1_hd U1166 ( .A(n1974), .B(n1908), .C(n1935), .Y(n1914) );
  oa21d1_hd U1167 ( .A(z_m[5]), .B(n1934), .C(n1914), .Y(n1909) );
  ao22d1_hd U1168 ( .A(z_m[6]), .B(n1909), .C(z_m[7]), .D(n1941), .Y(n1910) );
  oa211d1_hd U1169 ( .A(n1912), .B(n1926), .C(n1911), .D(n1910), .Y(n411) );
  ao22d1_hd U1170 ( .A(n1572), .B(sum[8]), .C(n1946), .D(sum[9]), .Y(n1918) );
  oa22d1_hd U1171 ( .A(n1914), .B(n1926), .C(n1913), .D(n1948), .Y(n1915) );
  ao21d1_hd U1172 ( .A(n1916), .B(n1926), .C(n1915), .Y(n1917) );
  oa211d1_hd U1173 ( .A(n1919), .B(n1959), .C(n1918), .D(n1917), .Y(n412) );
  ao22d1_hd U1174 ( .A(n1572), .B(sum[7]), .C(n1946), .D(sum[8]), .Y(n1925) );
  ao21d1_hd U1175 ( .A(n1974), .B(n1920), .C(n1935), .Y(n1929) );
  oa21d1_hd U1176 ( .A(z_m[3]), .B(n1934), .C(n1929), .Y(n1923) );
  oa21d1_hd U1177 ( .A(z_m[4]), .B(n1928), .C(n1959), .Y(n1922) );
  ao22d1_hd U1178 ( .A(z_m[4]), .B(n1923), .C(z_m[3]), .D(n1922), .Y(n1924) );
  oa211d1_hd U1179 ( .A(n1926), .B(n1948), .C(n1925), .D(n1924), .Y(n413) );
  ao22d1_hd U1180 ( .A(n1572), .B(sum[6]), .C(n1946), .D(sum[7]), .Y(n1932) );
  ao22d1_hd U1181 ( .A(z_m[3]), .B(n1929), .C(n1928), .D(n1927), .Y(n1930) );
  ao21d1_hd U1182 ( .A(z_m[4]), .B(n1941), .C(n1930), .Y(n1931) );
  scg15d1_hd U1183 ( .A(z_m[2]), .B(n1952), .C(n1932), .D(n1931), .Y(n414) );
  nr3d1_hd U1184 ( .A(z_m[2]), .B(n1934), .C(n1956), .Y(n1933) );
  nr2d1_hd U1185 ( .A(n1933), .B(n1952), .Y(n1939) );
  ao22d1_hd U1186 ( .A(n1572), .B(sum[5]), .C(n1946), .D(sum[6]), .Y(n1938) );
  nr2d1_hd U1187 ( .A(z_m[0]), .B(n1934), .Y(n1951) );
  nr2d1_hd U1188 ( .A(n1935), .B(n1951), .Y(n1945) );
  ao22d1_hd U1189 ( .A(z_m[2]), .B(n1936), .C(z_m[3]), .D(n1941), .Y(n1937) );
  oa211d1_hd U1190 ( .A(n1939), .B(n1949), .C(n1938), .D(n1937), .Y(n415) );
  ao22d1_hd U1191 ( .A(n1572), .B(sum[4]), .C(n1946), .D(sum[5]), .Y(n1944) );
  ao22d1_hd U1192 ( .A(z_m[0]), .B(n1942), .C(z_m[2]), .D(n1941), .Y(n1943) );
  oa211d1_hd U1193 ( .A(n1945), .B(n1949), .C(n1944), .D(n1943), .Y(n416) );
  ao22d1_hd U1194 ( .A(n1572), .B(sum[3]), .C(n1946), .D(sum[4]), .Y(n1954) );
  nr2d1_hd U1195 ( .A(n1949), .B(n1948), .Y(n1950) );
  ao211d1_hd U1196 ( .A(n1952), .B(guard), .C(n1951), .D(n1950), .Y(n1953) );
  oa211d1_hd U1197 ( .A(n1956), .B(n1955), .C(n1954), .D(n1953), .Y(n417) );
  ao21d1_hd U1198 ( .A(n1958), .B(n1968), .C(n1957), .Y(n1964) );
  oa21d1_hd U1199 ( .A(n1961), .B(n1960), .C(n1959), .Y(n1962) );
  ao22d1_hd U1200 ( .A(z_m[22]), .B(n1962), .C(n1975), .D(sum[26]), .Y(n1963)
         );
  oa211d1_hd U1201 ( .A(n1964), .B(n1967), .C(n1963), .D(n1972), .Y(n418) );
  nr4d1_hd U1202 ( .A(n1968), .B(n1967), .C(n1966), .D(n1965), .Y(n1969) );
  nd4d1_hd U1203 ( .A(z_m[21]), .B(z_m[20]), .C(n1970), .D(n1969), .Y(n1971)
         );
  nd4d1_hd U1204 ( .A(n1973), .B(n2272), .C(n1972), .D(n1971), .Y(n1987) );
  nr3d1_hd U1205 ( .A(n1975), .B(state[1]), .C(n1974), .Y(n1976) );
  ao22d1_hd U1206 ( .A(a_e[8]), .B(n1569), .C(n1993), .D(C91_DATA2_8), .Y(
        n1977) );
  oa21d1_hd U1207 ( .A(n1978), .B(n1987), .C(n1977), .Y(n419) );
  ao22d1_hd U1208 ( .A(z_e[7]), .B(n1989), .C(n1993), .D(C91_DATA2_7), .Y(
        n1979) );
  oa21d1_hd U1209 ( .A(n2104), .B(n2272), .C(n1979), .Y(n420) );
  ao22d1_hd U1210 ( .A(z_e[6]), .B(n1989), .C(n1993), .D(C91_DATA2_6), .Y(
        n1980) );
  oa21d1_hd U1211 ( .A(n2100), .B(n2272), .C(n1980), .Y(n421) );
  ao22d1_hd U1212 ( .A(z_e[5]), .B(n1989), .C(n1993), .D(C91_DATA2_5), .Y(
        n1981) );
  oa21d1_hd U1213 ( .A(n2119), .B(n2272), .C(n1981), .Y(n422) );
  ao22d1_hd U1214 ( .A(z_e[4]), .B(n1989), .C(n1993), .D(C91_DATA2_4), .Y(
        n1982) );
  oa21d1_hd U1215 ( .A(n2124), .B(n2272), .C(n1982), .Y(n423) );
  ao22d1_hd U1216 ( .A(z_e[3]), .B(n1989), .C(n1993), .D(C91_DATA2_3), .Y(
        n1983) );
  oa21d1_hd U1217 ( .A(n2131), .B(n2272), .C(n1983), .Y(n424) );
  ao22d1_hd U1218 ( .A(z_e[2]), .B(n1989), .C(n1993), .D(C91_DATA2_2), .Y(
        n1984) );
  oa21d1_hd U1219 ( .A(n2140), .B(n2272), .C(n1984), .Y(n425) );
  ao22d1_hd U1220 ( .A(z_e[1]), .B(n1989), .C(n1993), .D(C91_DATA2_1), .Y(
        n1985) );
  oa21d1_hd U1221 ( .A(n2148), .B(n2272), .C(n1985), .Y(n426) );
  ao22d1_hd U1222 ( .A(a_e[0]), .B(n1569), .C(n1993), .D(n1988), .Y(n1986) );
  oa21d1_hd U1223 ( .A(n1988), .B(n1987), .C(n1986), .Y(n427) );
  ao22d1_hd U1224 ( .A(a_e[9]), .B(n1569), .C(z_e[9]), .D(n1989), .Y(n1996) );
  ao22d1_hd U1225 ( .A(z_e[9]), .B(n2269), .C(n1991), .D(n1990), .Y(n1994) );
  oa211d1_hd U1226 ( .A(DP_OP_154J2_137_6175_n2), .B(n1994), .C(n1993), .D(
        n1992), .Y(n1995) );
  ao22d1_hd U1227 ( .A(b_m[25]), .B(n2039), .C(n1577), .D(b[21]), .Y(n1997) );
  oa21d1_hd U1228 ( .A(n1998), .B(n1575), .C(n1997), .Y(n429) );
  ao22d1_hd U1229 ( .A(b_m[24]), .B(n2039), .C(n1578), .D(b[20]), .Y(n1999) );
  oa21d1_hd U1230 ( .A(n2000), .B(n1575), .C(n1999), .Y(n430) );
  ao22d1_hd U1231 ( .A(b_m[23]), .B(n2039), .C(n1579), .D(b[19]), .Y(n2001) );
  oa21d1_hd U1232 ( .A(n2002), .B(n1575), .C(n2001), .Y(n431) );
  ao22d1_hd U1233 ( .A(b_m[22]), .B(n2039), .C(n1578), .D(b[18]), .Y(n2003) );
  oa21d1_hd U1234 ( .A(n2004), .B(n1575), .C(n2003), .Y(n432) );
  ao22d1_hd U1235 ( .A(b_m[21]), .B(n2039), .C(n1578), .D(b[17]), .Y(n2005) );
  oa21d1_hd U1236 ( .A(n2006), .B(n1575), .C(n2005), .Y(n433) );
  ao22d1_hd U1237 ( .A(b_m[20]), .B(n2039), .C(n1578), .D(b[16]), .Y(n2007) );
  oa21d1_hd U1238 ( .A(n2008), .B(n1575), .C(n2007), .Y(n434) );
  ao22d1_hd U1239 ( .A(b_m[19]), .B(n2039), .C(n1578), .D(b[15]), .Y(n2009) );
  oa21d1_hd U1240 ( .A(n2010), .B(n1575), .C(n2009), .Y(n435) );
  ao22d1_hd U1241 ( .A(b_m[18]), .B(n2039), .C(n1578), .D(b[14]), .Y(n2011) );
  oa21d1_hd U1242 ( .A(n2012), .B(n1575), .C(n2011), .Y(n436) );
  ao22d1_hd U1243 ( .A(b_m[17]), .B(n2039), .C(n1578), .D(b[13]), .Y(n2013) );
  oa21d1_hd U1244 ( .A(n2014), .B(n1575), .C(n2013), .Y(n437) );
  ao22d1_hd U1245 ( .A(b_m[16]), .B(n2039), .C(n1578), .D(b[12]), .Y(n2015) );
  oa21d1_hd U1246 ( .A(n2016), .B(n1575), .C(n2015), .Y(n438) );
  ao22d1_hd U1247 ( .A(b_m[15]), .B(n2039), .C(n1578), .D(b[11]), .Y(n2017) );
  oa21d1_hd U1248 ( .A(n2018), .B(n1575), .C(n2017), .Y(n439) );
  ao22d1_hd U1249 ( .A(b_m[14]), .B(n2039), .C(n1578), .D(b[10]), .Y(n2019) );
  oa21d1_hd U1250 ( .A(n2020), .B(n1575), .C(n2019), .Y(n440) );
  ao22d1_hd U1251 ( .A(b_m[13]), .B(n2039), .C(n1578), .D(b[9]), .Y(n2021) );
  oa21d1_hd U1252 ( .A(n2022), .B(n1575), .C(n2021), .Y(n441) );
  ao22d1_hd U1253 ( .A(b_m[12]), .B(n2039), .C(n1578), .D(b[8]), .Y(n2023) );
  oa21d1_hd U1254 ( .A(n2024), .B(n1575), .C(n2023), .Y(n442) );
  ao22d1_hd U1255 ( .A(b_m[11]), .B(n2039), .C(n1578), .D(b[7]), .Y(n2025) );
  oa21d1_hd U1256 ( .A(n2026), .B(n1575), .C(n2025), .Y(n443) );
  ao22d1_hd U1257 ( .A(b_m[10]), .B(n2039), .C(n1578), .D(b[6]), .Y(n2027) );
  oa21d1_hd U1258 ( .A(n2028), .B(n1575), .C(n2027), .Y(n444) );
  ao22d1_hd U1259 ( .A(b_m[9]), .B(n2039), .C(n1578), .D(b[5]), .Y(n2029) );
  oa21d1_hd U1260 ( .A(n2030), .B(n1575), .C(n2029), .Y(n445) );
  ao22d1_hd U1261 ( .A(b_m[8]), .B(n2039), .C(n1578), .D(b[4]), .Y(n2031) );
  oa21d1_hd U1262 ( .A(n2032), .B(n1575), .C(n2031), .Y(n446) );
  ao22d1_hd U1263 ( .A(b_m[7]), .B(n2039), .C(n1578), .D(b[3]), .Y(n2033) );
  oa21d1_hd U1264 ( .A(n2034), .B(n1575), .C(n2033), .Y(n447) );
  ao22d1_hd U1265 ( .A(b_m[6]), .B(n2039), .C(n1578), .D(b[2]), .Y(n2035) );
  oa21d1_hd U1266 ( .A(n2036), .B(n1575), .C(n2035), .Y(n448) );
  ao22d1_hd U1267 ( .A(b_m[5]), .B(n2039), .C(n1578), .D(b[1]), .Y(n2037) );
  oa21d1_hd U1268 ( .A(n2038), .B(n1575), .C(n2037), .Y(n449) );
  ao22d1_hd U1269 ( .A(b_m[4]), .B(n2039), .C(n1578), .D(b[0]), .Y(n2040) );
  oa21d1_hd U1270 ( .A(n2041), .B(n1575), .C(n2040), .Y(n450) );
  oa22d1_hd U1271 ( .A(n2042), .B(n1575), .C(n2041), .D(n2252), .Y(n451) );
  oa22d1_hd U1272 ( .A(n2043), .B(n1575), .C(n2042), .D(n2252), .Y(n452) );
  oa22d1_hd U1273 ( .A(n1579), .B(n2044), .C(n2043), .D(n2252), .Y(n453) );
  ao22d1_hd U1274 ( .A(a_m[25]), .B(n2087), .C(n1578), .D(a[21]), .Y(n2045) );
  oa21d1_hd U1275 ( .A(n2046), .B(n1573), .C(n2045), .Y(n454) );
  ao22d1_hd U1276 ( .A(a_m[24]), .B(n2087), .C(n1578), .D(a[20]), .Y(n2047) );
  oa21d1_hd U1277 ( .A(n2048), .B(n1573), .C(n2047), .Y(n455) );
  ao22d1_hd U1278 ( .A(a_m[23]), .B(n2087), .C(n1578), .D(a[19]), .Y(n2049) );
  oa21d1_hd U1279 ( .A(n2050), .B(n1573), .C(n2049), .Y(n456) );
  ao22d1_hd U1280 ( .A(a_m[22]), .B(n2087), .C(n1578), .D(a[18]), .Y(n2051) );
  oa21d1_hd U1281 ( .A(n2052), .B(n1573), .C(n2051), .Y(n457) );
  ao22d1_hd U1282 ( .A(a_m[21]), .B(n2087), .C(n1578), .D(a[17]), .Y(n2053) );
  oa21d1_hd U1283 ( .A(n2054), .B(n1573), .C(n2053), .Y(n458) );
  ao22d1_hd U1284 ( .A(a_m[20]), .B(n2087), .C(n1579), .D(a[16]), .Y(n2055) );
  oa21d1_hd U1285 ( .A(n2056), .B(n1573), .C(n2055), .Y(n459) );
  ao22d1_hd U1286 ( .A(a_m[19]), .B(n2087), .C(n1578), .D(a[15]), .Y(n2057) );
  oa21d1_hd U1287 ( .A(n2058), .B(n1573), .C(n2057), .Y(n460) );
  ao22d1_hd U1288 ( .A(a_m[18]), .B(n2087), .C(n1578), .D(a[14]), .Y(n2059) );
  oa21d1_hd U1289 ( .A(n2060), .B(n1573), .C(n2059), .Y(n461) );
  ao22d1_hd U1290 ( .A(a_m[17]), .B(n2087), .C(n1579), .D(a[13]), .Y(n2061) );
  oa21d1_hd U1291 ( .A(n2062), .B(n1573), .C(n2061), .Y(n462) );
  ao22d1_hd U1292 ( .A(a_m[16]), .B(n2087), .C(n1578), .D(a[12]), .Y(n2063) );
  oa21d1_hd U1293 ( .A(n2064), .B(n1573), .C(n2063), .Y(n463) );
  ao22d1_hd U1294 ( .A(a_m[15]), .B(n2087), .C(n1579), .D(a[11]), .Y(n2065) );
  oa21d1_hd U1295 ( .A(n2066), .B(n1573), .C(n2065), .Y(n464) );
  ao22d1_hd U1296 ( .A(a_m[14]), .B(n2087), .C(n1577), .D(a[10]), .Y(n2067) );
  oa21d1_hd U1297 ( .A(n2068), .B(n1573), .C(n2067), .Y(n465) );
  ao22d1_hd U1298 ( .A(a_m[13]), .B(n2087), .C(n1577), .D(a[9]), .Y(n2069) );
  oa21d1_hd U1299 ( .A(n2070), .B(n1573), .C(n2069), .Y(n466) );
  ao22d1_hd U1300 ( .A(a_m[12]), .B(n2087), .C(n1577), .D(a[8]), .Y(n2071) );
  oa21d1_hd U1301 ( .A(n2072), .B(n1573), .C(n2071), .Y(n467) );
  ao22d1_hd U1302 ( .A(a_m[11]), .B(n2087), .C(n1577), .D(a[7]), .Y(n2073) );
  oa21d1_hd U1303 ( .A(n2074), .B(n1573), .C(n2073), .Y(n468) );
  ao22d1_hd U1304 ( .A(a_m[10]), .B(n2087), .C(n1577), .D(a[6]), .Y(n2075) );
  oa21d1_hd U1305 ( .A(n2076), .B(n1573), .C(n2075), .Y(n469) );
  ao22d1_hd U1306 ( .A(a_m[9]), .B(n2087), .C(n1577), .D(a[5]), .Y(n2077) );
  oa21d1_hd U1307 ( .A(n2078), .B(n1573), .C(n2077), .Y(n470) );
  ao22d1_hd U1308 ( .A(a_m[8]), .B(n2087), .C(n1577), .D(a[4]), .Y(n2079) );
  oa21d1_hd U1309 ( .A(n2080), .B(n1573), .C(n2079), .Y(n471) );
  ao22d1_hd U1310 ( .A(a_m[7]), .B(n2087), .C(n1577), .D(a[3]), .Y(n2081) );
  oa21d1_hd U1311 ( .A(n2082), .B(n1573), .C(n2081), .Y(n472) );
  ao22d1_hd U1312 ( .A(a_m[6]), .B(n2087), .C(n1578), .D(a[2]), .Y(n2083) );
  oa21d1_hd U1313 ( .A(n2084), .B(n1573), .C(n2083), .Y(n473) );
  ao22d1_hd U1314 ( .A(a_m[5]), .B(n2087), .C(n1577), .D(a[1]), .Y(n2085) );
  oa21d1_hd U1315 ( .A(n2086), .B(n1573), .C(n2085), .Y(n474) );
  ao22d1_hd U1316 ( .A(a_m[4]), .B(n2087), .C(n1577), .D(a[0]), .Y(n2088) );
  oa21d1_hd U1317 ( .A(n2089), .B(n1573), .C(n2088), .Y(n475) );
  oa22d1_hd U1318 ( .A(n2090), .B(n1573), .C(n2089), .D(n2094), .Y(n476) );
  oa22d1_hd U1319 ( .A(n2091), .B(n1573), .C(n2090), .D(n2094), .Y(n477) );
  oa22d1_hd U1320 ( .A(n1579), .B(n2092), .C(n2091), .D(n2094), .Y(n478) );
  ao22d1_hd U1321 ( .A(a_m[25]), .B(n1574), .C(n1577), .D(a[22]), .Y(n2093) );
  oa21d1_hd U1322 ( .A(n2095), .B(n2094), .C(n2093), .Y(n479) );
  nr2d1_hd U1323 ( .A(n2148), .B(n2147), .Y(n2136) );
  nr2d1_hd U1324 ( .A(n2131), .B(n2130), .Y(n2121) );
  ao21d1_hd U1325 ( .A(n2189), .B(n2099), .C(n2154), .Y(n2120) );
  oa21d1_hd U1326 ( .A(n2100), .B(n2119), .C(n2189), .Y(n2098) );
  ao21d1_hd U1327 ( .A(n2139), .B(n2104), .C(n2106), .Y(n2156) );
  ivd1_hd U1328 ( .A(a[25]), .Y(n2138) );
  nr2d1_hd U1329 ( .A(n2150), .B(n2138), .Y(n2137) );
  ivd1_hd U1330 ( .A(a[27]), .Y(n2123) );
  nr2d1_hd U1331 ( .A(n2133), .B(n2123), .Y(n2122) );
  ivd1_hd U1332 ( .A(a[29]), .Y(n2109) );
  nr2d1_hd U1333 ( .A(n2116), .B(n2109), .Y(n2103) );
  nr2d1_hd U1334 ( .A(n2103), .B(n2268), .Y(n2111) );
  nr2d1_hd U1335 ( .A(n2157), .B(n2099), .Y(n2115) );
  nr2d1_hd U1336 ( .A(n2100), .B(n2114), .Y(n2105) );
  nd3d1_hd U1337 ( .A(a_e[7]), .B(n2105), .C(n2102), .Y(n2101) );
  oa211d1_hd U1338 ( .A(n2156), .B(n2102), .C(n2158), .D(n2101), .Y(n480) );
  ao22d1_hd U1339 ( .A(a_e[7]), .B(n2106), .C(n2105), .D(n2104), .Y(n2107) );
  oa211d1_hd U1340 ( .A(n2268), .B(n2108), .C(n2107), .D(n2158), .Y(n481) );
  oa21d1_hd U1341 ( .A(a_e[5]), .B(n2157), .C(n2120), .Y(n2112) );
  ao22d1_hd U1342 ( .A(a_e[6]), .B(n2112), .C(n2111), .D(n2110), .Y(n2113) );
  oa211d1_hd U1343 ( .A(a_e[6]), .B(n2114), .C(n2113), .D(n2143), .Y(n482) );
  ao21d1_hd U1344 ( .A(n2115), .B(n2119), .C(n2159), .Y(n2118) );
  oa211d1_hd U1345 ( .A(n2122), .B(a[28]), .C(n1579), .D(n2116), .Y(n2117) );
  oa211d1_hd U1346 ( .A(n2120), .B(n2119), .C(n2118), .D(n2117), .Y(n483) );
  ao211d1_hd U1347 ( .A(n2133), .B(n2123), .C(n2122), .D(n2268), .Y(n2126) );
  ao21d1_hd U1348 ( .A(n2189), .B(n2130), .C(n2154), .Y(n2132) );
  ao21d1_hd U1349 ( .A(n2132), .B(n2129), .C(n2124), .Y(n2125) );
  nr2d1_hd U1350 ( .A(n2126), .B(n2125), .Y(n2127) );
  oa211d1_hd U1351 ( .A(a_e[4]), .B(n2128), .C(n2127), .D(n2143), .Y(n484) );
  oa22d1_hd U1352 ( .A(n2132), .B(n2131), .C(n2130), .D(n2129), .Y(n2135) );
  oa211d1_hd U1353 ( .A(n2137), .B(a[26]), .C(n1579), .D(n2133), .Y(n2134) );
  scg13d1_hd U1354 ( .A(n2135), .B(n2159), .C(n2134), .Y(n485) );
  ao211d1_hd U1355 ( .A(n2150), .B(n2138), .C(n2137), .D(n2268), .Y(n2142) );
  nr2d1_hd U1356 ( .A(a_e[0]), .B(n2157), .Y(n2153) );
  nr2d1_hd U1357 ( .A(n2154), .B(n2153), .Y(n2149) );
  ao21d1_hd U1358 ( .A(n2149), .B(n2146), .C(n2140), .Y(n2141) );
  nr2d1_hd U1359 ( .A(n2142), .B(n2141), .Y(n2144) );
  oa211d1_hd U1360 ( .A(a_e[2]), .B(n2145), .C(n2144), .D(n2143), .Y(n486) );
  oa22d1_hd U1361 ( .A(n2149), .B(n2148), .C(n2147), .D(n2146), .Y(n2152) );
  oa211d1_hd U1362 ( .A(a[23]), .B(a[24]), .C(n1579), .D(n2150), .Y(n2151) );
  scg13d1_hd U1363 ( .A(n2152), .B(n2159), .C(n2151), .Y(n487) );
  ao21d1_hd U1364 ( .A(n2154), .B(a_e[0]), .C(n2153), .Y(n2155) );
  oa21d1_hd U1365 ( .A(a[23]), .B(n2268), .C(n2155), .Y(n488) );
  oa21d1_hd U1366 ( .A(a_e[8]), .B(n2157), .C(n2156), .Y(n2160) );
  scg17d1_hd U1367 ( .A(a_e[9]), .B(n2160), .C(n2159), .D(n2158), .Y(n489) );
  nr2d1_hd U1368 ( .A(n2215), .B(n2214), .Y(n2204) );
  nr2d1_hd U1369 ( .A(n2164), .B(n2198), .Y(n2194) );
  ao21d1_hd U1370 ( .A(n2165), .B(n2189), .C(n2221), .Y(n2188) );
  oa21d1_hd U1371 ( .A(n2167), .B(n2187), .C(n2189), .Y(n2166) );
  ao21d1_hd U1372 ( .A(n2205), .B(n2171), .C(n2173), .Y(n2254) );
  ivd1_hd U1373 ( .A(b[25]), .Y(n2207) );
  nr2d1_hd U1374 ( .A(n2217), .B(n2207), .Y(n2206) );
  ivd1_hd U1375 ( .A(b[27]), .Y(n2191) );
  nr2d1_hd U1376 ( .A(n2201), .B(n2191), .Y(n2190) );
  ivd1_hd U1377 ( .A(b[29]), .Y(n2177) );
  nr2d1_hd U1378 ( .A(n2184), .B(n2177), .Y(n2170) );
  nr2d1_hd U1379 ( .A(n2170), .B(n2268), .Y(n2180) );
  nr2bd1_hd U1380 ( .AN(n2194), .B(n2197), .Y(n2183) );
  nr2d1_hd U1381 ( .A(n2167), .B(n2182), .Y(n2172) );
  nd3d1_hd U1382 ( .A(b_e[7]), .B(n2172), .C(n2169), .Y(n2168) );
  oa211d1_hd U1383 ( .A(n2254), .B(n2169), .C(n2256), .D(n2168), .Y(n490) );
  ao22d1_hd U1384 ( .A(b_e[7]), .B(n2173), .C(n2172), .D(n2171), .Y(n2174) );
  oa211d1_hd U1385 ( .A(n2176), .B(n2175), .C(n2174), .D(n2256), .Y(n491) );
  oa21d1_hd U1386 ( .A(b_e[5]), .B(n2255), .C(n2188), .Y(n2178) );
  ao22d1_hd U1387 ( .A(n2180), .B(n2179), .C(b_e[6]), .D(n2178), .Y(n2181) );
  oa211d1_hd U1388 ( .A(b_e[6]), .B(n2182), .C(n2181), .D(n2210), .Y(n492) );
  ao21d1_hd U1389 ( .A(n2183), .B(n2187), .C(n2257), .Y(n2186) );
  oa211d1_hd U1390 ( .A(n2190), .B(b[28]), .C(n1579), .D(n2184), .Y(n2185) );
  oa211d1_hd U1391 ( .A(n2188), .B(n2187), .C(n2186), .D(n2185), .Y(n493) );
  scg6d1_hd U1392 ( .A(n2198), .B(n2189), .C(n2221), .Y(n2200) );
  ao211d1_hd U1393 ( .A(n2201), .B(n2191), .C(n2190), .D(n2268), .Y(n2192) );
  ao211d1_hd U1394 ( .A(b_e[4]), .B(n2200), .C(n2257), .D(n2192), .Y(n2196) );
  nd3d1_hd U1395 ( .A(n2205), .B(n2194), .C(n2193), .Y(n2195) );
  oa211d1_hd U1396 ( .A(b_e[3]), .B(n2197), .C(n2196), .D(n2195), .Y(n494) );
  nr3d1_hd U1397 ( .A(b_e[3]), .B(n2255), .C(n2198), .Y(n2199) );
  ao211d1_hd U1398 ( .A(b_e[3]), .B(n2200), .C(n2257), .D(n2199), .Y(n2203) );
  oa211d1_hd U1399 ( .A(n2206), .B(b[26]), .C(n1579), .D(n2201), .Y(n2202) );
  nr2d1_hd U1400 ( .A(b_e[0]), .B(n2255), .Y(n2220) );
  nr2d1_hd U1401 ( .A(n2221), .B(n2220), .Y(n2216) );
  ao211d1_hd U1402 ( .A(n2217), .B(n2207), .C(n2206), .D(n2268), .Y(n2208) );
  ao21d1_hd U1403 ( .A(n2209), .B(b_e[2]), .C(n2208), .Y(n2211) );
  oa211d1_hd U1404 ( .A(b_e[2]), .B(n2212), .C(n2211), .D(n2210), .Y(n496) );
  oa22d1_hd U1405 ( .A(n2216), .B(n2215), .C(n2214), .D(n2213), .Y(n2219) );
  oa211d1_hd U1406 ( .A(b[23]), .B(b[24]), .C(n1579), .D(n2217), .Y(n2218) );
  scg13d1_hd U1407 ( .A(n2219), .B(n2257), .C(n2218), .Y(n497) );
  ao21d1_hd U1408 ( .A(n2221), .B(b_e[0]), .C(n2220), .Y(n2222) );
  oa21d1_hd U1409 ( .A(b[23]), .B(n2268), .C(n2222), .Y(n498) );
  scg21d1_hd U1410 ( .A(n2223), .B(o_AB_ACK), .C(i_RST), .D(n1570), .Y(n499)
         );
  oa211d1_hd U1411 ( .A(state[3]), .B(n2228), .C(n2227), .D(n2226), .Y(n2242)
         );
  nd3d1_hd U1412 ( .A(n1580), .B(o_Z_STB), .C(i_Z_ACK), .Y(n2266) );
  nd4d1_hd U1413 ( .A(N41), .B(n2261), .C(n2266), .D(n2272), .Y(n2229) );
  nr3d1_hd U1414 ( .A(n27), .B(n2242), .C(n2229), .Y(n2234) );
  ao22d1_hd U1415 ( .A(n2232), .B(n2231), .C(n2269), .D(n2230), .Y(n2233) );
  oa211d1_hd U1416 ( .A(n2236), .B(n2235), .C(n2234), .D(n2233), .Y(n2262) );
  ivd1_hd U1417 ( .A(n2262), .Y(n2239) );
  nr2d1_hd U1418 ( .A(n2237), .B(n2247), .Y(n2238) );
  ao22d1_hd U1419 ( .A(state[2]), .B(n2239), .C(N41), .D(n2238), .Y(n2240) );
  oa21d1_hd U1420 ( .A(n2241), .B(n2264), .C(n2240), .Y(n500) );
  nr2d1_hd U1421 ( .A(n2269), .B(n2242), .Y(n2244) );
  oa22d1_hd U1422 ( .A(n2244), .B(n2264), .C(n2243), .D(n2262), .Y(n501) );
  oa211d1_hd U1423 ( .A(n2247), .B(state[0]), .C(n2246), .D(n2245), .Y(n2248)
         );
  ivd1_hd U1424 ( .A(n2248), .Y(n2250) );
  oa22d1_hd U1425 ( .A(n2250), .B(n2264), .C(n2249), .D(n2262), .Y(n502) );
  ao22d1_hd U1426 ( .A(b_m[25]), .B(n2161), .C(n1577), .D(b[22]), .Y(n2251) );
  oa21d1_hd U1427 ( .A(n2253), .B(n2252), .C(n2251), .Y(n503) );
  oa21d1_hd U1428 ( .A(b_e[8]), .B(n2255), .C(n2254), .Y(n2258) );
  scg17d1_hd U1429 ( .A(b_e[9]), .B(n2258), .C(n2257), .D(n2256), .Y(n504) );
  oa22d1_hd U1430 ( .A(n2265), .B(n2264), .C(n2263), .D(n2262), .Y(n505) );
  ivd1_hd U1431 ( .A(n2266), .Y(n2267) );
  scg21d1_hd U1432 ( .A(n1580), .B(o_Z_STB), .C(i_RST), .D(n2267), .Y(n506) );
endmodule


module iir_notch ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   w_add_1_AB_ACK, w_add_2_AB_ACK, w_add_1_Z_STB, w_add_2_Z_STB,
         r_add_1_AB_STB, r_add_1_Z_ACK, r_add_2_AB_STB, r_add_2_Z_ACK,
         w_mult_1_Z_STB, w_mult_2_Z_STB, w_mult_3_Z_STB, w_mult_1_AB_ACK,
         w_mult_2_AB_ACK, w_mult_3_AB_ACK, r_mult_1_AB_STB, r_mult_1_Z_ACK,
         n_2_net_, r_mult_2_AB_STB, r_mult_2_Z_ACK, n_3_net_, r_mult_3_AB_STB,
         r_mult_3_Z_ACK, n_4_net_, N23, r_pstate_0_, r_counter_1_, N739, N1343,
         N1383, N1396, N1401, N1402, N1403, n4, n5, n7, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n506, n542, n548, n557, n558,
         n559, n567, n568, n572, n573, n574, n576, n578, n580, n582, n584,
         n586, n588, n590, n592, n594, n596, n598, n600, n602, n604, n606,
         n608, n610, n612, n614, n616, n618, n620, n622, n624, n626, n628,
         n630, n632, n634, n647, n651, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n791, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079;
  wire   [31:0] r_add_1_A;
  wire   [31:0] r_add_1_B;
  wire   [31:0] w_add_1_Z;
  wire   [31:0] r_add_2_A;
  wire   [31:0] r_add_2_B;
  wire   [31:0] w_add_2_Z;
  wire   [31:0] r_mult_1_A;
  wire   [31:0] r_mult_1_B;
  wire   [31:0] w_mult_1_Z;
  wire   [31:0] r_mult_2_A;
  wire   [31:0] r_mult_2_B;
  wire   [31:0] w_mult_2_Z;
  wire   [31:0] r_mult_3_A;
  wire   [31:0] r_mult_3_B;
  wire   [31:0] w_mult_3_Z;
  wire   [159:0] r_x_data;
  wire   [127:0] r_y_data;

  float_adder_1 add_1 ( .i_A(r_add_1_A), .i_B(r_add_1_B), .i_AB_STB(
        r_add_1_AB_STB), .o_AB_ACK(w_add_1_AB_ACK), .o_Z(w_add_1_Z), .o_Z_STB(
        w_add_1_Z_STB), .i_Z_ACK(r_add_1_Z_ACK), .i_CLK(i_CLK), .i_RST(N23) );
  float_adder_0 add_2 ( .i_A(r_add_2_A), .i_B(r_add_2_B), .i_AB_STB(
        r_add_2_AB_STB), .o_AB_ACK(w_add_2_AB_ACK), .o_Z(w_add_2_Z), .o_Z_STB(
        w_add_2_Z_STB), .i_Z_ACK(r_add_2_Z_ACK), .i_CLK(i_CLK), .i_RST(N23) );
  float_multiplier mult_1 ( .i_A(r_mult_1_A), .i_B(r_mult_1_B), .i_AB_STB(
        r_mult_1_AB_STB), .o_AB_ACK(w_mult_1_AB_ACK), .o_Z(w_mult_1_Z), 
        .o_Z_STB(w_mult_1_Z_STB), .i_Z_ACK(r_mult_1_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(n_2_net_) );
  float_multiplier mult_2 ( .i_A(r_mult_2_A), .i_B(r_mult_2_B), .i_AB_STB(
        r_mult_2_AB_STB), .o_AB_ACK(w_mult_2_AB_ACK), .o_Z(w_mult_2_Z), 
        .o_Z_STB(w_mult_2_Z_STB), .i_Z_ACK(r_mult_2_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(n_3_net_) );
  float_multiplier mult_3 ( .i_A(r_mult_3_A), .i_B(r_mult_3_B), .i_AB_STB(
        r_mult_3_AB_STB), .o_AB_ACK(w_mult_3_AB_ACK), .o_Z(w_mult_3_Z), 
        .o_Z_STB(w_mult_3_Z_STB), .i_Z_ACK(r_mult_3_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(n_4_net_) );
  ivd1_hd I_10 ( .A(i_RSTN), .Y(n_4_net_) );
  ivd1_hd I_9 ( .A(i_RSTN), .Y(n_3_net_) );
  ivd1_hd I_8 ( .A(i_RSTN), .Y(n_2_net_) );
  scg4d1_hd U592 ( .A(n557), .B(r_add_2_A[31]), .C(n834), .D(r_x_data[63]), 
        .E(n558), .F(w_mult_2_Z[31]), .G(w_add_2_Z[31]), .H(n856), .Y(n692) );
  scg4d1_hd U593 ( .A(n557), .B(r_add_2_A[30]), .C(w_mult_2_Z[30]), .D(n558), 
        .E(r_x_data[62]), .F(n834), .G(n856), .H(w_add_2_Z[30]), .Y(n693) );
  scg4d1_hd U594 ( .A(n557), .B(r_add_2_A[29]), .C(w_mult_2_Z[29]), .D(n558), 
        .E(r_x_data[61]), .F(n834), .G(n856), .H(w_add_2_Z[29]), .Y(n694) );
  scg4d1_hd U595 ( .A(n557), .B(r_add_2_A[28]), .C(w_mult_2_Z[28]), .D(n558), 
        .E(r_x_data[60]), .F(n830), .G(n856), .H(w_add_2_Z[28]), .Y(n695) );
  scg4d1_hd U596 ( .A(n557), .B(r_add_2_A[27]), .C(w_mult_2_Z[27]), .D(n558), 
        .E(r_x_data[59]), .F(n830), .G(n856), .H(w_add_2_Z[27]), .Y(n696) );
  scg4d1_hd U597 ( .A(n557), .B(r_add_2_A[26]), .C(w_mult_2_Z[26]), .D(n558), 
        .E(r_x_data[58]), .F(n830), .G(n856), .H(w_add_2_Z[26]), .Y(n697) );
  scg4d1_hd U598 ( .A(n557), .B(r_add_2_A[25]), .C(w_mult_2_Z[25]), .D(n558), 
        .E(r_x_data[57]), .F(n832), .G(n856), .H(w_add_2_Z[25]), .Y(n698) );
  scg4d1_hd U599 ( .A(n557), .B(r_add_2_A[24]), .C(w_mult_2_Z[24]), .D(n558), 
        .E(r_x_data[56]), .F(n832), .G(n856), .H(w_add_2_Z[24]), .Y(n699) );
  scg4d1_hd U600 ( .A(n557), .B(r_add_2_A[23]), .C(w_mult_2_Z[23]), .D(n558), 
        .E(r_x_data[55]), .F(n830), .G(n856), .H(w_add_2_Z[23]), .Y(n700) );
  scg4d1_hd U601 ( .A(n557), .B(r_add_2_A[22]), .C(w_mult_2_Z[22]), .D(n558), 
        .E(r_x_data[54]), .F(n834), .G(n856), .H(w_add_2_Z[22]), .Y(n701) );
  scg4d1_hd U602 ( .A(n557), .B(r_add_2_A[21]), .C(w_mult_2_Z[21]), .D(n558), 
        .E(r_x_data[53]), .F(n834), .G(n856), .H(w_add_2_Z[21]), .Y(n702) );
  scg4d1_hd U603 ( .A(n557), .B(r_add_2_A[20]), .C(w_mult_2_Z[20]), .D(n558), 
        .E(r_x_data[52]), .F(n832), .G(n559), .H(w_add_2_Z[20]), .Y(n703) );
  scg4d1_hd U604 ( .A(n557), .B(r_add_2_A[19]), .C(w_mult_2_Z[19]), .D(n558), 
        .E(r_x_data[51]), .F(n832), .G(n559), .H(w_add_2_Z[19]), .Y(n704) );
  scg4d1_hd U605 ( .A(n557), .B(r_add_2_A[18]), .C(w_mult_2_Z[18]), .D(n558), 
        .E(r_x_data[50]), .F(n834), .G(n559), .H(w_add_2_Z[18]), .Y(n705) );
  scg4d1_hd U606 ( .A(n557), .B(r_add_2_A[17]), .C(w_mult_2_Z[17]), .D(n558), 
        .E(r_x_data[49]), .F(n832), .G(n559), .H(w_add_2_Z[17]), .Y(n706) );
  scg4d1_hd U607 ( .A(n557), .B(r_add_2_A[16]), .C(w_mult_2_Z[16]), .D(n558), 
        .E(r_x_data[48]), .F(n834), .G(n559), .H(w_add_2_Z[16]), .Y(n707) );
  scg4d1_hd U608 ( .A(n557), .B(r_add_2_A[15]), .C(w_mult_2_Z[15]), .D(n558), 
        .E(r_x_data[47]), .F(n832), .G(n559), .H(w_add_2_Z[15]), .Y(n708) );
  scg4d1_hd U609 ( .A(n557), .B(r_add_2_A[14]), .C(w_mult_2_Z[14]), .D(n558), 
        .E(r_x_data[46]), .F(n832), .G(n559), .H(w_add_2_Z[14]), .Y(n709) );
  scg4d1_hd U610 ( .A(n557), .B(r_add_2_A[13]), .C(w_mult_2_Z[13]), .D(n558), 
        .E(r_x_data[45]), .F(n830), .G(n559), .H(w_add_2_Z[13]), .Y(n710) );
  scg4d1_hd U611 ( .A(n557), .B(r_add_2_A[12]), .C(w_mult_2_Z[12]), .D(n558), 
        .E(r_x_data[44]), .F(n830), .G(n856), .H(w_add_2_Z[12]), .Y(n711) );
  scg4d1_hd U612 ( .A(n557), .B(r_add_2_A[11]), .C(w_mult_2_Z[11]), .D(n558), 
        .E(r_x_data[43]), .F(n834), .G(n559), .H(w_add_2_Z[11]), .Y(n712) );
  scg4d1_hd U613 ( .A(n557), .B(r_add_2_A[10]), .C(w_mult_2_Z[10]), .D(n558), 
        .E(r_x_data[42]), .F(n832), .G(n856), .H(w_add_2_Z[10]), .Y(n713) );
  scg4d1_hd U614 ( .A(n557), .B(r_add_2_A[9]), .C(w_mult_2_Z[9]), .D(n558), 
        .E(r_x_data[41]), .F(n832), .G(n559), .H(w_add_2_Z[9]), .Y(n714) );
  scg4d1_hd U615 ( .A(n557), .B(r_add_2_A[8]), .C(w_mult_2_Z[8]), .D(n558), 
        .E(r_x_data[40]), .F(n834), .G(n856), .H(w_add_2_Z[8]), .Y(n715) );
  scg4d1_hd U616 ( .A(n557), .B(r_add_2_A[7]), .C(w_mult_2_Z[7]), .D(n558), 
        .E(r_x_data[39]), .F(n832), .G(n559), .H(w_add_2_Z[7]), .Y(n716) );
  scg4d1_hd U617 ( .A(n557), .B(r_add_2_A[6]), .C(w_mult_2_Z[6]), .D(n558), 
        .E(r_x_data[38]), .F(n834), .G(n559), .H(w_add_2_Z[6]), .Y(n717) );
  scg4d1_hd U618 ( .A(n557), .B(r_add_2_A[5]), .C(w_mult_2_Z[5]), .D(n558), 
        .E(r_x_data[37]), .F(n830), .G(n856), .H(w_add_2_Z[5]), .Y(n718) );
  scg4d1_hd U619 ( .A(n557), .B(r_add_2_A[4]), .C(w_mult_2_Z[4]), .D(n558), 
        .E(r_x_data[36]), .F(n834), .G(n559), .H(w_add_2_Z[4]), .Y(n719) );
  scg4d1_hd U620 ( .A(n557), .B(r_add_2_A[3]), .C(w_mult_2_Z[3]), .D(n558), 
        .E(r_x_data[35]), .F(n830), .G(n559), .H(w_add_2_Z[3]), .Y(n720) );
  scg4d1_hd U621 ( .A(n557), .B(r_add_2_A[2]), .C(w_mult_2_Z[2]), .D(n558), 
        .E(r_x_data[34]), .F(n832), .G(n559), .H(w_add_2_Z[2]), .Y(n721) );
  scg4d1_hd U622 ( .A(n557), .B(r_add_2_A[1]), .C(w_mult_2_Z[1]), .D(n558), 
        .E(r_x_data[33]), .F(n834), .G(n559), .H(w_add_2_Z[1]), .Y(n722) );
  scg4d1_hd U623 ( .A(n557), .B(r_add_2_A[0]), .C(w_mult_2_Z[0]), .D(n558), 
        .E(r_x_data[32]), .F(n834), .G(n559), .H(w_add_2_Z[0]), .Y(n723) );
  scg4d1_hd U637 ( .A(n557), .B(r_add_2_B[21]), .C(w_mult_2_Z[21]), .D(n855), 
        .E(r_x_data[117]), .F(n832), .G(w_mult_3_Z[21]), .H(n854), .Y(n734) );
  scg4d1_hd U638 ( .A(n557), .B(r_add_2_B[20]), .C(w_mult_2_Z[20]), .D(n855), 
        .E(r_x_data[116]), .F(n834), .G(w_mult_3_Z[20]), .H(n568), .Y(n735) );
  scg4d1_hd U639 ( .A(n557), .B(r_add_2_B[19]), .C(w_mult_2_Z[19]), .D(n855), 
        .E(r_x_data[115]), .F(n832), .G(w_mult_3_Z[19]), .H(n854), .Y(n736) );
  scg4d1_hd U643 ( .A(n557), .B(r_add_2_B[15]), .C(w_mult_2_Z[15]), .D(n855), 
        .E(r_x_data[111]), .F(n832), .G(w_mult_3_Z[15]), .H(n854), .Y(n740) );
  ao22d1_hd U661 ( .A(w_mult_2_Z[30]), .B(n853), .C(w_mult_1_Z[30]), .D(n852), 
        .Y(n572) );
  ao22d1_hd U664 ( .A(w_mult_2_Z[29]), .B(n853), .C(w_mult_1_Z[29]), .D(n574), 
        .Y(n576) );
  ao22d1_hd U667 ( .A(w_mult_2_Z[28]), .B(n853), .C(w_mult_1_Z[28]), .D(n574), 
        .Y(n578) );
  ao22d1_hd U670 ( .A(w_mult_2_Z[27]), .B(n853), .C(w_mult_1_Z[27]), .D(n852), 
        .Y(n580) );
  ao22d1_hd U673 ( .A(w_mult_2_Z[26]), .B(n853), .C(w_mult_1_Z[26]), .D(n574), 
        .Y(n582) );
  ao22d1_hd U676 ( .A(w_mult_2_Z[25]), .B(n853), .C(w_mult_1_Z[25]), .D(n574), 
        .Y(n584) );
  ao22d1_hd U679 ( .A(w_mult_2_Z[24]), .B(n853), .C(w_mult_1_Z[24]), .D(n574), 
        .Y(n586) );
  ao22d1_hd U682 ( .A(w_mult_2_Z[23]), .B(n853), .C(w_mult_1_Z[23]), .D(n574), 
        .Y(n588) );
  ao22d1_hd U685 ( .A(w_mult_2_Z[22]), .B(n853), .C(w_mult_1_Z[22]), .D(n574), 
        .Y(n590) );
  ao22d1_hd U688 ( .A(w_mult_2_Z[21]), .B(n853), .C(w_mult_1_Z[21]), .D(n574), 
        .Y(n592) );
  ao22d1_hd U691 ( .A(w_mult_2_Z[20]), .B(n853), .C(w_mult_1_Z[20]), .D(n852), 
        .Y(n594) );
  ao22d1_hd U694 ( .A(w_mult_2_Z[19]), .B(n573), .C(w_mult_1_Z[19]), .D(n574), 
        .Y(n596) );
  ao22d1_hd U697 ( .A(w_mult_2_Z[18]), .B(n573), .C(w_mult_1_Z[18]), .D(n574), 
        .Y(n598) );
  ao22d1_hd U700 ( .A(w_mult_2_Z[17]), .B(n853), .C(w_mult_1_Z[17]), .D(n574), 
        .Y(n600) );
  ao22d1_hd U703 ( .A(w_mult_2_Z[16]), .B(n853), .C(w_mult_1_Z[16]), .D(n574), 
        .Y(n602) );
  ao22d1_hd U706 ( .A(w_mult_2_Z[15]), .B(n853), .C(w_mult_1_Z[15]), .D(n574), 
        .Y(n604) );
  ao22d1_hd U709 ( .A(w_mult_2_Z[14]), .B(n853), .C(w_mult_1_Z[14]), .D(n574), 
        .Y(n606) );
  ao22d1_hd U712 ( .A(w_mult_2_Z[13]), .B(n853), .C(w_mult_1_Z[13]), .D(n574), 
        .Y(n608) );
  ao22d1_hd U715 ( .A(w_mult_2_Z[12]), .B(n853), .C(w_mult_1_Z[12]), .D(n574), 
        .Y(n610) );
  ao22d1_hd U718 ( .A(w_mult_2_Z[11]), .B(n853), .C(w_mult_1_Z[11]), .D(n574), 
        .Y(n612) );
  ao22d1_hd U721 ( .A(w_mult_2_Z[10]), .B(n853), .C(w_mult_1_Z[10]), .D(n574), 
        .Y(n614) );
  ao22d1_hd U724 ( .A(w_mult_2_Z[9]), .B(n853), .C(w_mult_1_Z[9]), .D(n852), 
        .Y(n616) );
  ao22d1_hd U727 ( .A(w_mult_2_Z[8]), .B(n853), .C(w_mult_1_Z[8]), .D(n852), 
        .Y(n618) );
  ao22d1_hd U730 ( .A(w_mult_2_Z[7]), .B(n853), .C(w_mult_1_Z[7]), .D(n852), 
        .Y(n620) );
  ao22d1_hd U733 ( .A(w_mult_2_Z[6]), .B(n853), .C(w_mult_1_Z[6]), .D(n852), 
        .Y(n622) );
  ao22d1_hd U736 ( .A(w_mult_2_Z[5]), .B(n853), .C(w_mult_1_Z[5]), .D(n852), 
        .Y(n624) );
  ao22d1_hd U739 ( .A(w_mult_2_Z[4]), .B(n573), .C(w_mult_1_Z[4]), .D(n852), 
        .Y(n626) );
  ao22d1_hd U742 ( .A(w_mult_2_Z[3]), .B(n853), .C(w_mult_1_Z[3]), .D(n852), 
        .Y(n628) );
  ao22d1_hd U745 ( .A(w_mult_2_Z[2]), .B(n853), .C(w_mult_1_Z[2]), .D(n852), 
        .Y(n630) );
  ao22d1_hd U748 ( .A(w_mult_2_Z[1]), .B(n573), .C(w_mult_1_Z[1]), .D(n852), 
        .Y(n632) );
  ao22d1_hd U751 ( .A(w_mult_2_Z[0]), .B(n853), .C(w_mult_1_Z[0]), .D(n852), 
        .Y(n634) );
  scg4d1_hd U765 ( .A(n557), .B(r_add_2_B[31]), .C(n834), .D(r_x_data[127]), 
        .E(n855), .F(w_mult_2_Z[31]), .G(w_mult_3_Z[31]), .H(n854), .Y(n794)
         );
  ao22d1_hd U802 ( .A(n853), .B(w_mult_2_Z[31]), .C(w_mult_1_Z[31]), .D(n852), 
        .Y(n651) );
  ivd1_hd U833 ( .A(i_RSTN), .Y(N23) );
  fd2qd1_hd r_counter_reg_1_ ( .D(n791), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_counter_1_) );
  fd1eqd1_hd r_mult_3_AB_STB_reg ( .D(N1343), .E(N1403), .CK(i_CLK), .Q(
        r_mult_3_AB_STB) );
  fd2qd1_hd r_mult_3_Z_ACK_reg ( .D(n497), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_Z_ACK) );
  fd2qd1_hd r_mult_1_AB_STB_reg ( .D(n491), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_AB_STB) );
  fd2qd1_hd r_mult_2_AB_STB_reg ( .D(n490), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_AB_STB) );
  fd2qd1_hd r_mult_2_A_reg_2_ ( .D(n169), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[2]) );
  fd2qd1_hd r_mult_2_A_reg_11_ ( .D(n160), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[11]) );
  fd2qd1_hd r_mult_2_A_reg_16_ ( .D(n155), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[16]) );
  fd2qd1_hd r_mult_2_A_reg_23_ ( .D(n148), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[23]) );
  fd2qd1_hd r_mult_2_A_reg_30_ ( .D(n141), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[30]) );
  fd2qd1_hd r_mult_3_A_reg_30_ ( .D(n78), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[30]) );
  fd2qd1_hd r_mult_2_A_reg_1_ ( .D(n170), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[1]) );
  fd2qd1_hd r_mult_2_A_reg_4_ ( .D(n167), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[4]) );
  fd2qd1_hd r_mult_2_A_reg_7_ ( .D(n164), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[7]) );
  fd2qd1_hd r_mult_2_A_reg_9_ ( .D(n162), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[9]) );
  fd2qd1_hd r_mult_2_A_reg_13_ ( .D(n158), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[13]) );
  fd2qd1_hd r_mult_2_A_reg_14_ ( .D(n157), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[14]) );
  fd2qd1_hd r_mult_2_A_reg_19_ ( .D(n152), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[19]) );
  fd2qd1_hd r_mult_2_A_reg_20_ ( .D(n151), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[20]) );
  fd2qd1_hd r_mult_2_A_reg_21_ ( .D(n150), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[21]) );
  fd2qd1_hd r_mult_2_A_reg_31_ ( .D(n140), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[31]) );
  fd2qd1_hd r_mult_3_A_reg_2_ ( .D(n106), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[2]) );
  fd2qd1_hd r_mult_3_A_reg_10_ ( .D(n98), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[10]) );
  fd2qd1_hd r_mult_3_A_reg_11_ ( .D(n97), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[11]) );
  fd2qd1_hd r_mult_3_A_reg_15_ ( .D(n93), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[15]) );
  fd2qd1_hd r_mult_3_A_reg_18_ ( .D(n90), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[18]) );
  fd2qd1_hd r_mult_3_A_reg_21_ ( .D(n87), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[21]) );
  fd2qd1_hd r_mult_3_A_reg_22_ ( .D(n86), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[22]) );
  fd2qd1_hd r_mult_3_A_reg_23_ ( .D(n85), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[23]) );
  fd2qd1_hd r_mult_3_A_reg_24_ ( .D(n84), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[24]) );
  fd2qd1_hd r_mult_3_A_reg_31_ ( .D(n77), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[31]) );
  fd2qd1_hd r_mult_3_B_reg_31_ ( .D(n501), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[31]) );
  fd2qd1_hd r_mult_3_B_reg_0_ ( .D(n139), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[0]) );
  fd2qd1_hd r_mult_3_B_reg_1_ ( .D(n138), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[1]) );
  fd2qd1_hd r_mult_3_B_reg_2_ ( .D(n137), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[2]) );
  fd2qd1_hd r_mult_3_B_reg_3_ ( .D(n136), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[3]) );
  fd2qd1_hd r_mult_3_B_reg_4_ ( .D(n135), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[4]) );
  fd2qd1_hd r_mult_3_B_reg_5_ ( .D(n134), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[5]) );
  fd2qd1_hd r_mult_3_B_reg_6_ ( .D(n133), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[6]) );
  fd2qd1_hd r_mult_3_B_reg_7_ ( .D(n132), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[7]) );
  fd2qd1_hd r_mult_3_B_reg_8_ ( .D(n131), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[8]) );
  fd2qd1_hd r_mult_3_B_reg_9_ ( .D(n130), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[9]) );
  fd2qd1_hd r_mult_3_B_reg_10_ ( .D(n129), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[10]) );
  fd2qd1_hd r_mult_3_B_reg_11_ ( .D(n128), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[11]) );
  fd2qd1_hd r_mult_3_B_reg_12_ ( .D(n127), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[12]) );
  fd2qd1_hd r_mult_3_B_reg_13_ ( .D(n126), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[13]) );
  fd2qd1_hd r_mult_3_B_reg_14_ ( .D(n125), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[14]) );
  fd2qd1_hd r_mult_3_B_reg_15_ ( .D(n124), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[15]) );
  fd2qd1_hd r_mult_3_B_reg_16_ ( .D(n123), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[16]) );
  fd2qd1_hd r_mult_3_B_reg_17_ ( .D(n122), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[17]) );
  fd2qd1_hd r_mult_3_B_reg_18_ ( .D(n121), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[18]) );
  fd2qd1_hd r_mult_3_B_reg_19_ ( .D(n120), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[19]) );
  fd2qd1_hd r_mult_3_B_reg_20_ ( .D(n119), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[20]) );
  fd2qd1_hd r_mult_3_B_reg_21_ ( .D(n118), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[21]) );
  fd2qd1_hd r_mult_3_B_reg_22_ ( .D(n117), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[22]) );
  fd2qd1_hd r_mult_3_B_reg_23_ ( .D(n116), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[23]) );
  fd2qd1_hd r_mult_3_B_reg_24_ ( .D(n115), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[24]) );
  fd2qd1_hd r_mult_3_B_reg_25_ ( .D(n114), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[25]) );
  fd2qd1_hd r_mult_3_B_reg_26_ ( .D(n113), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[26]) );
  fd2qd1_hd r_mult_3_B_reg_27_ ( .D(n112), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[27]) );
  fd2qd1_hd r_mult_3_B_reg_28_ ( .D(n111), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[28]) );
  fd2qd1_hd r_mult_3_B_reg_29_ ( .D(n110), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[29]) );
  fd2qd1_hd r_mult_3_B_reg_30_ ( .D(n109), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_0_ ( .D(n76), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[0]) );
  fd2qd1_hd r_mult_1_B_reg_1_ ( .D(n75), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[1]) );
  fd2qd1_hd r_mult_1_B_reg_2_ ( .D(n74), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[2]) );
  fd2qd1_hd r_mult_1_B_reg_3_ ( .D(n73), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[3]) );
  fd2qd1_hd r_mult_1_B_reg_4_ ( .D(n72), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[4]) );
  fd2qd1_hd r_mult_1_B_reg_5_ ( .D(n71), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[5]) );
  fd2qd1_hd r_mult_1_B_reg_6_ ( .D(n70), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[6]) );
  fd2qd1_hd r_mult_1_B_reg_7_ ( .D(n69), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[7]) );
  fd2qd1_hd r_mult_1_B_reg_8_ ( .D(n68), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[8]) );
  fd2qd1_hd r_mult_1_B_reg_9_ ( .D(n67), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[9]) );
  fd2qd1_hd r_mult_1_B_reg_10_ ( .D(n66), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[10]) );
  fd2qd1_hd r_mult_1_B_reg_11_ ( .D(n65), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[11]) );
  fd2qd1_hd r_mult_1_B_reg_12_ ( .D(n64), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[12]) );
  fd2qd1_hd r_mult_1_B_reg_13_ ( .D(n63), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[13]) );
  fd2qd1_hd r_mult_1_B_reg_14_ ( .D(n62), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[14]) );
  fd2qd1_hd r_mult_1_B_reg_15_ ( .D(n61), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[15]) );
  fd2qd1_hd r_mult_1_B_reg_16_ ( .D(n60), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[16]) );
  fd2qd1_hd r_mult_1_B_reg_17_ ( .D(n59), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[17]) );
  fd2qd1_hd r_mult_1_B_reg_18_ ( .D(n58), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[18]) );
  fd2qd1_hd r_mult_1_B_reg_19_ ( .D(n57), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[19]) );
  fd2qd1_hd r_mult_1_B_reg_20_ ( .D(n56), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[20]) );
  fd2qd1_hd r_mult_1_B_reg_21_ ( .D(n55), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[21]) );
  fd2qd1_hd r_mult_1_B_reg_22_ ( .D(n54), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[22]) );
  fd2qd1_hd r_mult_1_B_reg_30_ ( .D(n46), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_31_ ( .D(n45), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[31]) );
  fd2qd1_hd r_mult_2_B_reg_31_ ( .D(n499), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[31]) );
  fd2qd1_hd r_mult_1_Z_ACK_reg ( .D(n493), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_Z_ACK) );
  fd2qd1_hd r_mult_2_Z_ACK_reg ( .D(n492), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_Z_ACK) );
  fd2qd1_hd r_mult_2_B_reg_0_ ( .D(n202), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[0]) );
  fd2qd1_hd r_mult_2_B_reg_1_ ( .D(n201), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[1]) );
  fd2qd1_hd r_mult_2_B_reg_2_ ( .D(n200), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[2]) );
  fd2qd1_hd r_mult_2_B_reg_3_ ( .D(n199), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[3]) );
  fd2qd1_hd r_mult_2_B_reg_4_ ( .D(n198), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[4]) );
  fd2qd1_hd r_mult_2_B_reg_5_ ( .D(n197), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[5]) );
  fd2qd1_hd r_mult_2_B_reg_6_ ( .D(n196), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[6]) );
  fd2qd1_hd r_mult_2_B_reg_7_ ( .D(n195), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[7]) );
  fd2qd1_hd r_mult_2_B_reg_8_ ( .D(n194), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[8]) );
  fd2qd1_hd r_mult_2_B_reg_9_ ( .D(n193), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[9]) );
  fd2qd1_hd r_mult_2_B_reg_10_ ( .D(n192), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[10]) );
  fd2qd1_hd r_mult_2_B_reg_11_ ( .D(n191), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[11]) );
  fd2qd1_hd r_mult_2_B_reg_12_ ( .D(n190), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[12]) );
  fd2qd1_hd r_mult_2_B_reg_13_ ( .D(n189), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[13]) );
  fd2qd1_hd r_mult_2_B_reg_14_ ( .D(n188), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[14]) );
  fd2qd1_hd r_mult_2_B_reg_15_ ( .D(n187), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[15]) );
  fd2qd1_hd r_mult_2_B_reg_16_ ( .D(n186), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[16]) );
  fd2qd1_hd r_mult_2_B_reg_17_ ( .D(n185), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[17]) );
  fd2qd1_hd r_mult_2_B_reg_18_ ( .D(n184), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[18]) );
  fd2qd1_hd r_mult_2_B_reg_19_ ( .D(n183), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[19]) );
  fd2qd1_hd r_mult_2_B_reg_20_ ( .D(n182), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[20]) );
  fd2qd1_hd r_mult_2_B_reg_21_ ( .D(n181), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[21]) );
  fd2qd1_hd r_mult_2_B_reg_22_ ( .D(n180), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[22]) );
  fd2qd1_hd r_mult_2_B_reg_23_ ( .D(n179), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[23]) );
  fd2qd1_hd r_mult_2_B_reg_24_ ( .D(n178), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[24]) );
  fd2qd1_hd r_mult_2_B_reg_25_ ( .D(n177), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[25]) );
  fd2qd1_hd r_mult_2_B_reg_26_ ( .D(n176), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[26]) );
  fd2qd1_hd r_mult_2_B_reg_27_ ( .D(n175), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[27]) );
  fd2qd1_hd r_mult_2_B_reg_28_ ( .D(n174), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[28]) );
  fd2qd1_hd r_mult_2_B_reg_29_ ( .D(n173), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[29]) );
  fd2qd1_hd r_mult_2_B_reg_30_ ( .D(n172), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[30]) );
  fd2qd1_hd r_mult_2_A_reg_12_ ( .D(n159), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[12]) );
  fd2qd1_hd r_mult_2_A_reg_18_ ( .D(n153), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[18]) );
  fd2qd1_hd r_mult_1_B_reg_23_ ( .D(n53), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[23]) );
  fd2qd1_hd r_mult_1_B_reg_24_ ( .D(n52), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[24]) );
  fd2qd1_hd r_mult_1_B_reg_25_ ( .D(n51), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[25]) );
  fd2qd1_hd r_mult_1_B_reg_26_ ( .D(n50), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[26]) );
  fd2qd1_hd r_mult_1_B_reg_27_ ( .D(n49), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[27]) );
  fd2qd1_hd r_mult_1_B_reg_28_ ( .D(n48), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[28]) );
  fd2qd1_hd r_mult_1_B_reg_29_ ( .D(n47), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[29]) );
  fd2qd1_hd r_mult_2_A_reg_0_ ( .D(n171), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[0]) );
  fd2qd1_hd r_mult_2_A_reg_5_ ( .D(n166), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[5]) );
  fd2qd1_hd r_mult_2_A_reg_15_ ( .D(n156), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[15]) );
  fd2qd1_hd r_mult_2_A_reg_17_ ( .D(n154), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[17]) );
  fd2qd1_hd r_mult_2_A_reg_24_ ( .D(n147), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[24]) );
  fd2qd1_hd r_mult_3_A_reg_0_ ( .D(n108), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[0]) );
  fd2qd1_hd r_mult_3_A_reg_1_ ( .D(n107), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[1]) );
  fd2qd1_hd r_mult_3_A_reg_6_ ( .D(n102), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[6]) );
  fd2qd1_hd r_mult_3_A_reg_8_ ( .D(n100), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[8]) );
  fd2qd1_hd r_mult_3_A_reg_9_ ( .D(n99), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[9]) );
  fd2qd1_hd r_mult_3_A_reg_13_ ( .D(n95), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[13]) );
  fd2qd1_hd r_mult_3_A_reg_14_ ( .D(n94), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[14]) );
  fd2qd1_hd r_mult_3_A_reg_16_ ( .D(n92), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[16]) );
  fd2qd1_hd r_mult_3_A_reg_19_ ( .D(n89), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[19]) );
  fd2qd1_hd r_mult_3_A_reg_20_ ( .D(n88), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[20]) );
  fd2qd1_hd r_mult_2_A_reg_3_ ( .D(n168), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[3]) );
  fd2qd1_hd r_mult_2_A_reg_6_ ( .D(n165), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[6]) );
  fd2qd1_hd r_mult_2_A_reg_8_ ( .D(n163), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[8]) );
  fd2qd1_hd r_mult_2_A_reg_10_ ( .D(n161), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[10]) );
  fd2qd1_hd r_mult_2_A_reg_22_ ( .D(n149), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[22]) );
  fd2qd1_hd r_mult_2_A_reg_25_ ( .D(n146), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[25]) );
  fd2qd1_hd r_mult_2_A_reg_26_ ( .D(n145), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[26]) );
  fd2qd1_hd r_mult_2_A_reg_27_ ( .D(n144), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[27]) );
  fd2qd1_hd r_mult_2_A_reg_28_ ( .D(n143), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[28]) );
  fd2qd1_hd r_mult_2_A_reg_29_ ( .D(n142), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_0_ ( .D(n502), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[0]) );
  fd2qd1_hd r_mult_1_A_reg_2_ ( .D(n43), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[2]) );
  fd2qd1_hd r_mult_1_A_reg_3_ ( .D(n42), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[3]) );
  fd2qd1_hd r_mult_1_A_reg_4_ ( .D(n41), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[4]) );
  fd2qd1_hd r_mult_1_A_reg_5_ ( .D(n40), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[5]) );
  fd2qd1_hd r_mult_1_A_reg_7_ ( .D(n38), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[7]) );
  fd2qd1_hd r_mult_1_A_reg_10_ ( .D(n35), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[10]) );
  fd2qd1_hd r_mult_1_A_reg_11_ ( .D(n34), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[11]) );
  fd2qd1_hd r_mult_1_A_reg_13_ ( .D(n32), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[13]) );
  fd2qd1_hd r_mult_1_A_reg_14_ ( .D(n31), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[14]) );
  fd2qd1_hd r_mult_1_A_reg_15_ ( .D(n30), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[15]) );
  fd2qd1_hd r_mult_1_A_reg_17_ ( .D(n28), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[17]) );
  fd2qd1_hd r_mult_1_A_reg_18_ ( .D(n27), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[18]) );
  fd2qd1_hd r_mult_1_A_reg_19_ ( .D(n26), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[19]) );
  fd2qd1_hd r_mult_1_A_reg_21_ ( .D(n24), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[21]) );
  fd2qd1_hd r_mult_1_A_reg_22_ ( .D(n23), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[22]) );
  fd2qd1_hd r_mult_1_A_reg_23_ ( .D(n22), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[23]) );
  fd2qd1_hd r_mult_1_A_reg_24_ ( .D(n21), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[24]) );
  fd2qd1_hd r_mult_1_A_reg_25_ ( .D(n20), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[25]) );
  fd2qd1_hd r_mult_1_A_reg_26_ ( .D(n19), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[26]) );
  fd2qd1_hd r_mult_1_A_reg_27_ ( .D(n18), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[27]) );
  fd2qd1_hd r_mult_1_A_reg_28_ ( .D(n17), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[28]) );
  fd2qd1_hd r_mult_1_A_reg_29_ ( .D(n16), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_1_ ( .D(n44), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_6_ ( .D(n39), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[6]) );
  fd2qd1_hd r_mult_1_A_reg_8_ ( .D(n37), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[8]) );
  fd2qd1_hd r_mult_1_A_reg_9_ ( .D(n36), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[9]) );
  fd2qd1_hd r_mult_1_A_reg_12_ ( .D(n33), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[12]) );
  fd2qd1_hd r_mult_1_A_reg_16_ ( .D(n29), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[16]) );
  fd2qd1_hd r_mult_1_A_reg_20_ ( .D(n25), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[20]) );
  fd2qd1_hd r_mult_1_A_reg_30_ ( .D(n15), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[30]) );
  fd2qd1_hd r_mult_1_A_reg_31_ ( .D(n14), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[31]) );
  fd2qd1_hd r_add_2_B_reg_31_ ( .D(n794), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[31]) );
  fd2qd1_hd r_add_1_B_reg_19_ ( .D(n672), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[19]) );
  fd2qd1_hd r_add_2_B_reg_0_ ( .D(n755), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[0]) );
  fd2qd1_hd r_add_2_A_reg_0_ ( .D(n723), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[0]) );
  fd2qd1_hd r_add_2_B_reg_1_ ( .D(n754), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[1]) );
  fd2qd1_hd r_add_2_A_reg_1_ ( .D(n722), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[1]) );
  fd2qd1_hd r_add_2_B_reg_2_ ( .D(n753), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[2]) );
  fd2qd1_hd r_add_2_A_reg_2_ ( .D(n721), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[2]) );
  fd2qd1_hd r_add_2_B_reg_3_ ( .D(n752), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[3]) );
  fd2qd1_hd r_add_2_A_reg_3_ ( .D(n720), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[3]) );
  fd2qd1_hd r_add_2_B_reg_4_ ( .D(n751), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[4]) );
  fd2qd1_hd r_add_2_A_reg_4_ ( .D(n719), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[4]) );
  fd2qd1_hd r_add_2_B_reg_5_ ( .D(n750), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[5]) );
  fd2qd1_hd r_add_2_A_reg_5_ ( .D(n718), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[5]) );
  fd2qd1_hd r_add_2_B_reg_6_ ( .D(n749), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[6]) );
  fd2qd1_hd r_add_2_A_reg_6_ ( .D(n717), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[6]) );
  fd2qd1_hd r_add_2_B_reg_7_ ( .D(n748), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[7]) );
  fd2qd1_hd r_add_2_A_reg_7_ ( .D(n716), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[7]) );
  fd2qd1_hd r_add_2_B_reg_8_ ( .D(n747), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[8]) );
  fd2qd1_hd r_add_2_A_reg_8_ ( .D(n715), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[8]) );
  fd2qd1_hd r_add_2_B_reg_9_ ( .D(n746), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[9]) );
  fd2qd1_hd r_add_2_A_reg_9_ ( .D(n714), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[9]) );
  fd2qd1_hd r_add_2_B_reg_10_ ( .D(n745), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[10]) );
  fd2qd1_hd r_add_2_A_reg_10_ ( .D(n713), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[10]) );
  fd2qd1_hd r_add_2_B_reg_11_ ( .D(n744), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[11]) );
  fd2qd1_hd r_add_2_A_reg_11_ ( .D(n712), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[11]) );
  fd2qd1_hd r_add_2_B_reg_12_ ( .D(n743), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[12]) );
  fd2qd1_hd r_add_2_A_reg_12_ ( .D(n711), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[12]) );
  fd2qd1_hd r_add_2_B_reg_13_ ( .D(n742), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[13]) );
  fd2qd1_hd r_add_2_A_reg_13_ ( .D(n710), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[13]) );
  fd2qd1_hd r_add_2_B_reg_14_ ( .D(n741), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[14]) );
  fd2qd1_hd r_add_2_A_reg_14_ ( .D(n709), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[14]) );
  fd2qd1_hd r_add_2_B_reg_15_ ( .D(n740), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[15]) );
  fd2qd1_hd r_add_2_A_reg_15_ ( .D(n708), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[15]) );
  fd2qd1_hd r_add_2_B_reg_16_ ( .D(n739), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[16]) );
  fd2qd1_hd r_add_2_A_reg_16_ ( .D(n707), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[16]) );
  fd2qd1_hd r_add_2_B_reg_17_ ( .D(n738), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[17]) );
  fd2qd1_hd r_add_2_A_reg_17_ ( .D(n706), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[17]) );
  fd2qd1_hd r_add_2_B_reg_18_ ( .D(n737), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[18]) );
  fd2qd1_hd r_add_2_A_reg_18_ ( .D(n705), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[18]) );
  fd2qd1_hd r_add_2_B_reg_19_ ( .D(n736), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[19]) );
  fd2qd1_hd r_add_2_A_reg_19_ ( .D(n704), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[19]) );
  fd2qd1_hd r_add_2_B_reg_20_ ( .D(n735), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[20]) );
  fd2qd1_hd r_add_2_A_reg_20_ ( .D(n703), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[20]) );
  fd2qd1_hd r_add_2_B_reg_21_ ( .D(n734), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[21]) );
  fd2qd1_hd r_add_2_A_reg_21_ ( .D(n702), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[21]) );
  fd2qd1_hd r_add_2_B_reg_22_ ( .D(n733), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[22]) );
  fd2qd1_hd r_add_2_A_reg_22_ ( .D(n701), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[22]) );
  fd2qd1_hd r_add_2_B_reg_23_ ( .D(n732), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[23]) );
  fd2qd1_hd r_add_2_A_reg_23_ ( .D(n700), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[23]) );
  fd2qd1_hd r_add_2_B_reg_24_ ( .D(n731), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[24]) );
  fd2qd1_hd r_add_2_A_reg_24_ ( .D(n699), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[24]) );
  fd2qd1_hd r_add_2_B_reg_25_ ( .D(n730), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[25]) );
  fd2qd1_hd r_add_2_A_reg_25_ ( .D(n698), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[25]) );
  fd2qd1_hd r_add_2_B_reg_26_ ( .D(n729), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[26]) );
  fd2qd1_hd r_add_2_A_reg_26_ ( .D(n697), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[26]) );
  fd2qd1_hd r_add_2_B_reg_27_ ( .D(n728), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[27]) );
  fd2qd1_hd r_add_2_A_reg_27_ ( .D(n696), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[27]) );
  fd2qd1_hd r_add_2_B_reg_28_ ( .D(n727), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[28]) );
  fd2qd1_hd r_add_2_A_reg_28_ ( .D(n695), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[28]) );
  fd2qd1_hd r_add_2_B_reg_29_ ( .D(n726), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[29]) );
  fd2qd1_hd r_add_2_A_reg_29_ ( .D(n694), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[29]) );
  fd2qd1_hd r_add_2_B_reg_30_ ( .D(n725), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[30]) );
  fd2qd1_hd r_add_2_A_reg_30_ ( .D(n693), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[30]) );
  fd2qd1_hd r_add_2_A_reg_31_ ( .D(n692), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[31]) );
  fd2qd1_hd r_add_1_B_reg_31_ ( .D(n660), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[31]) );
  fd2qd1_hd r_add_1_B_reg_0_ ( .D(n691), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[0]) );
  fd2qd1_hd r_add_1_B_reg_1_ ( .D(n690), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[1]) );
  fd2qd1_hd r_add_1_B_reg_2_ ( .D(n689), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[2]) );
  fd2qd1_hd r_add_1_B_reg_3_ ( .D(n688), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[3]) );
  fd2qd1_hd r_add_1_B_reg_4_ ( .D(n687), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[4]) );
  fd2qd1_hd r_add_1_B_reg_5_ ( .D(n686), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[5]) );
  fd2qd1_hd r_add_1_B_reg_6_ ( .D(n685), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[6]) );
  fd2qd1_hd r_add_1_B_reg_7_ ( .D(n684), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[7]) );
  fd2qd1_hd r_add_1_B_reg_8_ ( .D(n683), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[8]) );
  fd2qd1_hd r_add_1_B_reg_9_ ( .D(n682), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[9]) );
  fd2qd1_hd r_add_1_B_reg_10_ ( .D(n681), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[10]) );
  fd2qd1_hd r_add_1_B_reg_11_ ( .D(n680), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[11]) );
  fd2qd1_hd r_add_1_B_reg_12_ ( .D(n679), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[12]) );
  fd2qd1_hd r_add_1_B_reg_13_ ( .D(n678), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[13]) );
  fd2qd1_hd r_add_1_B_reg_14_ ( .D(n677), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[14]) );
  fd2qd1_hd r_add_1_B_reg_15_ ( .D(n676), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[15]) );
  fd2qd1_hd r_add_1_B_reg_16_ ( .D(n675), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[16]) );
  fd2qd1_hd r_add_1_B_reg_17_ ( .D(n674), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[17]) );
  fd2qd1_hd r_add_1_B_reg_18_ ( .D(n673), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[18]) );
  fd2qd1_hd r_add_1_B_reg_20_ ( .D(n671), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[20]) );
  fd2qd1_hd r_add_1_B_reg_21_ ( .D(n670), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[21]) );
  fd2qd1_hd r_add_1_B_reg_22_ ( .D(n669), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[22]) );
  fd2qd1_hd r_add_1_B_reg_23_ ( .D(n668), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[23]) );
  fd2qd1_hd r_add_1_B_reg_24_ ( .D(n667), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[24]) );
  fd2qd1_hd r_add_1_B_reg_25_ ( .D(n666), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[25]) );
  fd2qd1_hd r_add_1_B_reg_26_ ( .D(n665), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[26]) );
  fd2qd1_hd r_add_1_B_reg_27_ ( .D(n664), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[27]) );
  fd2qd1_hd r_add_1_B_reg_28_ ( .D(n663), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[28]) );
  fd2qd1_hd r_add_1_B_reg_29_ ( .D(n662), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[29]) );
  fd2qd1_hd r_add_1_B_reg_30_ ( .D(n661), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[30]) );
  fd2qd1_hd r_x_data_reg_147_ ( .D(n342), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[147]) );
  fd2qd1_hd r_x_data_reg_128_ ( .D(n361), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[128]) );
  fd2qd1_hd r_x_data_reg_129_ ( .D(n360), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[129]) );
  fd2qd1_hd r_x_data_reg_130_ ( .D(n359), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[130]) );
  fd2qd1_hd r_x_data_reg_131_ ( .D(n358), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[131]) );
  fd2qd1_hd r_x_data_reg_132_ ( .D(n357), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[132]) );
  fd2qd1_hd r_x_data_reg_133_ ( .D(n356), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[133]) );
  fd2qd1_hd r_x_data_reg_134_ ( .D(n355), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[134]) );
  fd2qd1_hd r_x_data_reg_135_ ( .D(n354), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[135]) );
  fd2qd1_hd r_x_data_reg_136_ ( .D(n353), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[136]) );
  fd2qd1_hd r_x_data_reg_137_ ( .D(n352), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[137]) );
  fd2qd1_hd r_x_data_reg_138_ ( .D(n351), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[138]) );
  fd2qd1_hd r_x_data_reg_139_ ( .D(n350), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[139]) );
  fd2qd1_hd r_x_data_reg_140_ ( .D(n349), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[140]) );
  fd2qd1_hd r_x_data_reg_141_ ( .D(n348), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[141]) );
  fd2qd1_hd r_x_data_reg_142_ ( .D(n347), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[142]) );
  fd2qd1_hd r_x_data_reg_143_ ( .D(n346), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[143]) );
  fd2qd1_hd r_x_data_reg_144_ ( .D(n345), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[144]) );
  fd2qd1_hd r_x_data_reg_145_ ( .D(n344), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[145]) );
  fd2qd1_hd r_x_data_reg_146_ ( .D(n343), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[146]) );
  fd2qd1_hd r_x_data_reg_148_ ( .D(n341), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[148]) );
  fd2qd1_hd r_x_data_reg_149_ ( .D(n340), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[149]) );
  fd2qd1_hd r_x_data_reg_150_ ( .D(n339), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[150]) );
  fd2qd1_hd r_x_data_reg_151_ ( .D(n338), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[151]) );
  fd2qd1_hd r_x_data_reg_152_ ( .D(n337), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[152]) );
  fd2qd1_hd r_x_data_reg_153_ ( .D(n336), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[153]) );
  fd2qd1_hd r_x_data_reg_154_ ( .D(n335), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[154]) );
  fd2qd1_hd r_x_data_reg_155_ ( .D(n334), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[155]) );
  fd2qd1_hd r_x_data_reg_156_ ( .D(n333), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[156]) );
  fd2qd1_hd r_x_data_reg_157_ ( .D(n332), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[157]) );
  fd2qd1_hd r_x_data_reg_158_ ( .D(n331), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[158]) );
  fd2qd1_hd r_x_data_reg_159_ ( .D(n330), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[159]) );
  fd2qd1_hd r_y_data_reg_96_ ( .D(n234), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[96]) );
  fd2qd1_hd r_y_data_reg_97_ ( .D(n233), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[97]) );
  fd2qd1_hd r_y_data_reg_98_ ( .D(n232), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[98]) );
  fd2qd1_hd r_y_data_reg_99_ ( .D(n231), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[99]) );
  fd2qd1_hd r_y_data_reg_100_ ( .D(n230), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[100]) );
  fd2qd1_hd r_y_data_reg_101_ ( .D(n229), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[101]) );
  fd2qd1_hd r_y_data_reg_102_ ( .D(n228), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[102]) );
  fd2qd1_hd r_y_data_reg_103_ ( .D(n227), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[103]) );
  fd2qd1_hd r_y_data_reg_104_ ( .D(n226), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[104]) );
  fd2qd1_hd r_y_data_reg_105_ ( .D(n225), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[105]) );
  fd2qd1_hd r_y_data_reg_106_ ( .D(n224), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[106]) );
  fd2qd1_hd r_y_data_reg_107_ ( .D(n223), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[107]) );
  fd2qd1_hd r_y_data_reg_108_ ( .D(n222), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[108]) );
  fd2qd1_hd r_y_data_reg_109_ ( .D(n221), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[109]) );
  fd2qd1_hd r_y_data_reg_110_ ( .D(n220), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[110]) );
  fd2qd1_hd r_y_data_reg_111_ ( .D(n219), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[111]) );
  fd2qd1_hd r_y_data_reg_112_ ( .D(n218), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[112]) );
  fd2qd1_hd r_y_data_reg_113_ ( .D(n217), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[113]) );
  fd2qd1_hd r_y_data_reg_114_ ( .D(n216), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[114]) );
  fd2qd1_hd r_y_data_reg_115_ ( .D(n215), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[115]) );
  fd2qd1_hd r_y_data_reg_116_ ( .D(n214), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[116]) );
  fd2qd1_hd r_y_data_reg_117_ ( .D(n213), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[117]) );
  fd2qd1_hd r_y_data_reg_118_ ( .D(n212), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[118]) );
  fd2qd1_hd r_y_data_reg_119_ ( .D(n211), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[119]) );
  fd2qd1_hd r_y_data_reg_120_ ( .D(n210), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[120]) );
  fd2qd1_hd r_y_data_reg_121_ ( .D(n209), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[121]) );
  fd2qd1_hd r_y_data_reg_122_ ( .D(n208), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[122]) );
  fd2qd1_hd r_y_data_reg_123_ ( .D(n207), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[123]) );
  fd2qd1_hd r_y_data_reg_124_ ( .D(n206), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[124]) );
  fd2qd1_hd r_y_data_reg_125_ ( .D(n205), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[125]) );
  fd2qd1_hd r_y_data_reg_126_ ( .D(n204), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[126]) );
  fd2qd1_hd r_y_data_reg_127_ ( .D(n203), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[127]) );
  fd2qd1_hd r_add_1_A_reg_0_ ( .D(n787), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[0]) );
  fd2qd1_hd r_add_1_A_reg_1_ ( .D(n786), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[1]) );
  fd2qd1_hd r_add_1_A_reg_2_ ( .D(n785), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[2]) );
  fd2qd1_hd r_add_1_A_reg_3_ ( .D(n784), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[3]) );
  fd2qd1_hd r_add_1_A_reg_4_ ( .D(n783), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[4]) );
  fd2qd1_hd r_add_1_A_reg_5_ ( .D(n782), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[5]) );
  fd2qd1_hd r_add_1_A_reg_6_ ( .D(n781), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[6]) );
  fd2qd1_hd r_add_1_A_reg_7_ ( .D(n780), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[7]) );
  fd2qd1_hd r_add_1_A_reg_8_ ( .D(n779), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[8]) );
  fd2qd1_hd r_add_1_A_reg_9_ ( .D(n778), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[9]) );
  fd2qd1_hd r_add_1_A_reg_10_ ( .D(n777), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[10]) );
  fd2qd1_hd r_add_1_A_reg_11_ ( .D(n776), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[11]) );
  fd2qd1_hd r_add_1_A_reg_12_ ( .D(n775), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[12]) );
  fd2qd1_hd r_add_1_A_reg_13_ ( .D(n774), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[13]) );
  fd2qd1_hd r_add_1_A_reg_14_ ( .D(n773), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[14]) );
  fd2qd1_hd r_add_1_A_reg_15_ ( .D(n772), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[15]) );
  fd2qd1_hd r_add_1_A_reg_16_ ( .D(n771), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[16]) );
  fd2qd1_hd r_add_1_A_reg_17_ ( .D(n770), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[17]) );
  fd2qd1_hd r_add_1_A_reg_18_ ( .D(n769), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[18]) );
  fd2qd1_hd r_add_1_A_reg_19_ ( .D(n768), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[19]) );
  fd2qd1_hd r_add_1_A_reg_20_ ( .D(n767), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[20]) );
  fd2qd1_hd r_add_1_A_reg_21_ ( .D(n766), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[21]) );
  fd2qd1_hd r_add_1_A_reg_22_ ( .D(n765), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[22]) );
  fd2qd1_hd r_add_1_A_reg_23_ ( .D(n764), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[23]) );
  fd2qd1_hd r_add_1_A_reg_24_ ( .D(n763), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[24]) );
  fd2qd1_hd r_add_1_A_reg_25_ ( .D(n762), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[25]) );
  fd2qd1_hd r_add_1_A_reg_26_ ( .D(n761), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[26]) );
  fd2qd1_hd r_add_1_A_reg_27_ ( .D(n760), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[27]) );
  fd2qd1_hd r_add_1_A_reg_28_ ( .D(n759), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[28]) );
  fd2qd1_hd r_add_1_A_reg_29_ ( .D(n758), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[29]) );
  fd2qd1_hd r_add_1_A_reg_30_ ( .D(n757), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[30]) );
  fd2qd1_hd r_add_1_A_reg_31_ ( .D(n826), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[31]) );
  fd2qd1_hd r_mult_3_A_reg_3_ ( .D(n105), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[3]) );
  fd2qd1_hd r_mult_3_A_reg_4_ ( .D(n104), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[4]) );
  fd2qd1_hd r_mult_3_A_reg_5_ ( .D(n103), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[5]) );
  fd2qd1_hd r_mult_3_A_reg_7_ ( .D(n101), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[7]) );
  fd2qd1_hd r_mult_3_A_reg_12_ ( .D(n96), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[12]) );
  fd2qd1_hd r_mult_3_A_reg_17_ ( .D(n91), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[17]) );
  fd2qd1_hd r_mult_3_A_reg_25_ ( .D(n83), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[25]) );
  fd2qd1_hd r_mult_3_A_reg_26_ ( .D(n82), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[26]) );
  fd2qd1_hd r_mult_3_A_reg_27_ ( .D(n81), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[27]) );
  fd2qd1_hd r_mult_3_A_reg_28_ ( .D(n80), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[28]) );
  fd2qd1_hd r_mult_3_A_reg_29_ ( .D(n79), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[29]) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(n827), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[31]) );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(n795), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[0]) );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(n796), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[1]) );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(n797), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[2]) );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(n798), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[3]) );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(n799), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[4]) );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(n800), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[5]) );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(n801), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[6]) );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(n802), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[7]) );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(n803), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[8]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(n804), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[9]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(n805), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(n806), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(n807), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(n808), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(n809), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(n810), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(n811), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(n812), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(n813), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(n814), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(n815), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(n816), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(n817), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(n818), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(n819), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(n820), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(n821), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(n822), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(n823), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(n824), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(n825), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd r_x_data_reg_64_ ( .D(n425), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[64]) );
  fd2qd1_hd r_x_data_reg_65_ ( .D(n424), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[65]) );
  fd2qd1_hd r_x_data_reg_66_ ( .D(n423), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[66]) );
  fd2qd1_hd r_x_data_reg_67_ ( .D(n422), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[67]) );
  fd2qd1_hd r_x_data_reg_68_ ( .D(n421), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[68]) );
  fd2qd1_hd r_x_data_reg_69_ ( .D(n420), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[69]) );
  fd2qd1_hd r_x_data_reg_70_ ( .D(n419), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[70]) );
  fd2qd1_hd r_x_data_reg_71_ ( .D(n418), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[71]) );
  fd2qd1_hd r_x_data_reg_72_ ( .D(n417), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[72]) );
  fd2qd1_hd r_x_data_reg_73_ ( .D(n416), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[73]) );
  fd2qd1_hd r_x_data_reg_74_ ( .D(n415), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[74]) );
  fd2qd1_hd r_x_data_reg_75_ ( .D(n414), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[75]) );
  fd2qd1_hd r_x_data_reg_76_ ( .D(n413), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[76]) );
  fd2qd1_hd r_x_data_reg_77_ ( .D(n412), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[77]) );
  fd2qd1_hd r_x_data_reg_78_ ( .D(n411), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[78]) );
  fd2qd1_hd r_x_data_reg_79_ ( .D(n410), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[79]) );
  fd2qd1_hd r_x_data_reg_80_ ( .D(n409), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[80]) );
  fd2qd1_hd r_x_data_reg_81_ ( .D(n408), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[81]) );
  fd2qd1_hd r_x_data_reg_82_ ( .D(n407), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[82]) );
  fd2qd1_hd r_x_data_reg_83_ ( .D(n406), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[83]) );
  fd2qd1_hd r_x_data_reg_84_ ( .D(n405), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[84]) );
  fd2qd1_hd r_x_data_reg_85_ ( .D(n404), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[85]) );
  fd2qd1_hd r_x_data_reg_86_ ( .D(n403), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[86]) );
  fd2qd1_hd r_x_data_reg_94_ ( .D(n395), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[94]) );
  fd2qd1_hd r_x_data_reg_95_ ( .D(n394), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[95]) );
  fd2qd1_hd r_y_data_reg_64_ ( .D(n266), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[64]) );
  fd2qd1_hd r_y_data_reg_65_ ( .D(n265), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[65]) );
  fd2qd1_hd r_y_data_reg_66_ ( .D(n264), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[66]) );
  fd2qd1_hd r_y_data_reg_67_ ( .D(n263), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[67]) );
  fd2qd1_hd r_y_data_reg_68_ ( .D(n262), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[68]) );
  fd2qd1_hd r_y_data_reg_69_ ( .D(n261), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[69]) );
  fd2qd1_hd r_y_data_reg_70_ ( .D(n260), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[70]) );
  fd2qd1_hd r_y_data_reg_71_ ( .D(n259), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[71]) );
  fd2qd1_hd r_y_data_reg_72_ ( .D(n258), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[72]) );
  fd2qd1_hd r_y_data_reg_73_ ( .D(n257), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[73]) );
  fd2qd1_hd r_y_data_reg_74_ ( .D(n256), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[74]) );
  fd2qd1_hd r_y_data_reg_75_ ( .D(n255), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[75]) );
  fd2qd1_hd r_y_data_reg_76_ ( .D(n254), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[76]) );
  fd2qd1_hd r_y_data_reg_77_ ( .D(n253), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[77]) );
  fd2qd1_hd r_y_data_reg_78_ ( .D(n252), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[78]) );
  fd2qd1_hd r_y_data_reg_79_ ( .D(n251), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[79]) );
  fd2qd1_hd r_y_data_reg_80_ ( .D(n250), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[80]) );
  fd2qd1_hd r_y_data_reg_81_ ( .D(n249), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[81]) );
  fd2qd1_hd r_y_data_reg_82_ ( .D(n248), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[82]) );
  fd2qd1_hd r_y_data_reg_83_ ( .D(n247), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[83]) );
  fd2qd1_hd r_y_data_reg_84_ ( .D(n246), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[84]) );
  fd2qd1_hd r_y_data_reg_85_ ( .D(n245), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[85]) );
  fd2qd1_hd r_y_data_reg_86_ ( .D(n244), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[86]) );
  fd2qd1_hd r_y_data_reg_87_ ( .D(n243), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[87]) );
  fd2qd1_hd r_y_data_reg_88_ ( .D(n242), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[88]) );
  fd2qd1_hd r_y_data_reg_89_ ( .D(n241), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[89]) );
  fd2qd1_hd r_y_data_reg_90_ ( .D(n240), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[90]) );
  fd2qd1_hd r_y_data_reg_91_ ( .D(n239), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[91]) );
  fd2qd1_hd r_y_data_reg_92_ ( .D(n238), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[92]) );
  fd2qd1_hd r_y_data_reg_93_ ( .D(n237), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[93]) );
  fd2qd1_hd r_y_data_reg_94_ ( .D(n236), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[94]) );
  fd2qd1_hd r_y_data_reg_95_ ( .D(n235), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[95]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(n500), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_x_data_reg_32_ ( .D(n457), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[32]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(n456), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(n455), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[34]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(n454), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(n453), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(n452), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[37]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(n451), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(n450), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(n449), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(n448), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(n447), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(n446), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(n445), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(n444), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(n443), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(n442), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(n441), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(n440), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(n439), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(n438), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[51]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(n437), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(n436), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(n435), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(n434), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(n433), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(n432), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(n431), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[58]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(n430), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(n429), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(n428), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(n427), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_96_ ( .D(n393), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[96]) );
  fd2qd1_hd r_x_data_reg_97_ ( .D(n392), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[97]) );
  fd2qd1_hd r_x_data_reg_98_ ( .D(n391), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[98]) );
  fd2qd1_hd r_x_data_reg_99_ ( .D(n390), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[99]) );
  fd2qd1_hd r_x_data_reg_100_ ( .D(n389), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[100]) );
  fd2qd1_hd r_x_data_reg_101_ ( .D(n388), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[101]) );
  fd2qd1_hd r_x_data_reg_102_ ( .D(n387), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[102]) );
  fd2qd1_hd r_x_data_reg_103_ ( .D(n386), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[103]) );
  fd2qd1_hd r_x_data_reg_104_ ( .D(n385), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[104]) );
  fd2qd1_hd r_x_data_reg_105_ ( .D(n384), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[105]) );
  fd2qd1_hd r_x_data_reg_106_ ( .D(n383), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[106]) );
  fd2qd1_hd r_x_data_reg_107_ ( .D(n382), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[107]) );
  fd2qd1_hd r_x_data_reg_108_ ( .D(n381), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[108]) );
  fd2qd1_hd r_x_data_reg_109_ ( .D(n380), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[109]) );
  fd2qd1_hd r_x_data_reg_110_ ( .D(n379), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[110]) );
  fd2qd1_hd r_x_data_reg_111_ ( .D(n378), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[111]) );
  fd2qd1_hd r_x_data_reg_112_ ( .D(n377), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[112]) );
  fd2qd1_hd r_x_data_reg_113_ ( .D(n376), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[113]) );
  fd2qd1_hd r_x_data_reg_114_ ( .D(n375), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[114]) );
  fd2qd1_hd r_x_data_reg_115_ ( .D(n374), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[115]) );
  fd2qd1_hd r_x_data_reg_116_ ( .D(n373), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[116]) );
  fd2qd1_hd r_x_data_reg_117_ ( .D(n372), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[117]) );
  fd2qd1_hd r_x_data_reg_118_ ( .D(n371), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[118]) );
  fd2qd1_hd r_x_data_reg_119_ ( .D(n370), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[119]) );
  fd2qd1_hd r_x_data_reg_120_ ( .D(n369), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[120]) );
  fd2qd1_hd r_x_data_reg_121_ ( .D(n368), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[121]) );
  fd2qd1_hd r_x_data_reg_122_ ( .D(n367), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[122]) );
  fd2qd1_hd r_x_data_reg_123_ ( .D(n366), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[123]) );
  fd2qd1_hd r_x_data_reg_124_ ( .D(n365), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[124]) );
  fd2qd1_hd r_x_data_reg_125_ ( .D(n364), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[125]) );
  fd2qd1_hd r_x_data_reg_126_ ( .D(n363), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[126]) );
  fd2qd1_hd r_y_data_reg_0_ ( .D(n329), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[0]) );
  fd2qd1_hd r_y_data_reg_1_ ( .D(n328), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[1]) );
  fd2qd1_hd r_y_data_reg_2_ ( .D(n327), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[2]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(n326), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[3]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(n325), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(n324), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(n323), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(n322), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(n321), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(n320), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(n319), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(n318), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(n317), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(n316), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(n315), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(n314), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(n313), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(n312), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(n311), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(n310), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(n309), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(n308), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(n307), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(n306), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(n305), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(n304), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(n303), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(n302), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(n301), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(n300), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(n299), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_32_ ( .D(n298), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[32]) );
  fd2qd1_hd r_y_data_reg_33_ ( .D(n297), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[33]) );
  fd2qd1_hd r_y_data_reg_34_ ( .D(n296), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[34]) );
  fd2qd1_hd r_y_data_reg_35_ ( .D(n295), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[35]) );
  fd2qd1_hd r_y_data_reg_36_ ( .D(n294), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[36]) );
  fd2qd1_hd r_y_data_reg_37_ ( .D(n293), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[37]) );
  fd2qd1_hd r_y_data_reg_38_ ( .D(n292), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[38]) );
  fd2qd1_hd r_y_data_reg_39_ ( .D(n291), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[39]) );
  fd2qd1_hd r_y_data_reg_40_ ( .D(n290), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[40]) );
  fd2qd1_hd r_y_data_reg_41_ ( .D(n289), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[41]) );
  fd2qd1_hd r_y_data_reg_42_ ( .D(n288), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[42]) );
  fd2qd1_hd r_y_data_reg_43_ ( .D(n287), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[43]) );
  fd2qd1_hd r_y_data_reg_44_ ( .D(n286), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[44]) );
  fd2qd1_hd r_y_data_reg_45_ ( .D(n285), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[45]) );
  fd2qd1_hd r_y_data_reg_46_ ( .D(n284), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[46]) );
  fd2qd1_hd r_y_data_reg_47_ ( .D(n283), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[47]) );
  fd2qd1_hd r_y_data_reg_48_ ( .D(n282), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[48]) );
  fd2qd1_hd r_y_data_reg_49_ ( .D(n281), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[49]) );
  fd2qd1_hd r_y_data_reg_50_ ( .D(n280), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[50]) );
  fd2qd1_hd r_y_data_reg_51_ ( .D(n279), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[51]) );
  fd2qd1_hd r_y_data_reg_52_ ( .D(n278), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[52]) );
  fd2qd1_hd r_y_data_reg_53_ ( .D(n277), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[53]) );
  fd2qd1_hd r_y_data_reg_54_ ( .D(n276), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[54]) );
  fd2qd1_hd r_y_data_reg_55_ ( .D(n275), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[55]) );
  fd2qd1_hd r_y_data_reg_56_ ( .D(n274), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[56]) );
  fd2qd1_hd r_y_data_reg_57_ ( .D(n273), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[57]) );
  fd2qd1_hd r_y_data_reg_58_ ( .D(n272), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[58]) );
  fd2qd1_hd r_y_data_reg_59_ ( .D(n271), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[59]) );
  fd2qd1_hd r_y_data_reg_60_ ( .D(n270), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[60]) );
  fd2qd1_hd r_y_data_reg_61_ ( .D(n269), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[61]) );
  fd2qd1_hd r_y_data_reg_62_ ( .D(n268), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[62]) );
  fd2qd1_hd r_y_data_reg_63_ ( .D(n267), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[63]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(n426), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[63]) );
  fd2qd1_hd r_x_data_reg_127_ ( .D(n362), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[127]) );
  fd2qd1_hd r_x_data_reg_87_ ( .D(n402), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[87]) );
  fd2qd1_hd r_x_data_reg_88_ ( .D(n401), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[88]) );
  fd2qd1_hd r_x_data_reg_89_ ( .D(n400), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[89]) );
  fd2qd1_hd r_x_data_reg_90_ ( .D(n399), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[90]) );
  fd2qd1_hd r_x_data_reg_91_ ( .D(n398), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[91]) );
  fd2qd1_hd r_x_data_reg_92_ ( .D(n397), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[92]) );
  fd2qd1_hd r_x_data_reg_93_ ( .D(n396), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[93]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(n489), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(n488), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(n487), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(n486), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(n485), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(n484), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[5]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(n483), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(n482), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(n481), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(n480), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(n479), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(n478), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(n477), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(n476), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(n475), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(n474), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(n473), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(n472), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(n471), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(n470), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(n469), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(n468), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(n467), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(n466), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(n465), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(n464), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(n463), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(n462), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(n461), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(n460), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(n459), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(n458), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[31]) );
  fd2qd1_hd r_add_1_Z_ACK_reg ( .D(n793), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_Z_ACK) );
  fd2qd1_hd r_add_2_Z_ACK_reg ( .D(n756), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_Z_ACK) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n724), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_add_1_AB_STB_reg ( .D(n789), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_AB_STB) );
  fd2qd1_hd r_add_2_AB_STB_reg ( .D(n788), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_AB_STB) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n833), .E(N1402), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(N1383), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_pstate_0_) );
  scg4d1_hd U641 ( .A(n557), .B(r_add_2_B[17]), .C(w_mult_2_Z[17]), .D(n855), 
        .E(r_x_data[113]), .F(n834), .G(w_mult_3_Z[17]), .H(n854), .Y(n738) );
  scg4d1_hd U644 ( .A(n557), .B(r_add_2_B[14]), .C(w_mult_2_Z[14]), .D(n855), 
        .E(r_x_data[110]), .F(n832), .G(w_mult_3_Z[14]), .H(n854), .Y(n741) );
  scg4d1_hd U635 ( .A(n557), .B(r_add_2_B[23]), .C(w_mult_2_Z[23]), .D(n855), 
        .E(r_x_data[119]), .F(n832), .G(w_mult_3_Z[23]), .H(n854), .Y(n732) );
  scg4d1_hd U647 ( .A(n557), .B(r_add_2_B[11]), .C(w_mult_2_Z[11]), .D(n855), 
        .E(r_x_data[107]), .F(n830), .G(w_mult_3_Z[11]), .H(n854), .Y(n744) );
  scg4d1_hd U648 ( .A(n557), .B(r_add_2_B[10]), .C(w_mult_2_Z[10]), .D(n855), 
        .E(r_x_data[106]), .F(n830), .G(w_mult_3_Z[10]), .H(n854), .Y(n745) );
  scg4d1_hd U658 ( .A(n557), .B(r_add_2_B[0]), .C(w_mult_2_Z[0]), .D(n855), 
        .E(r_x_data[96]), .F(n830), .G(w_mult_3_Z[0]), .H(n854), .Y(n755) );
  scg4d1_hd U654 ( .A(n557), .B(r_add_2_B[4]), .C(w_mult_2_Z[4]), .D(n855), 
        .E(r_x_data[100]), .F(n832), .G(w_mult_3_Z[4]), .H(n854), .Y(n751) );
  scg4d1_hd U657 ( .A(n557), .B(r_add_2_B[1]), .C(w_mult_2_Z[1]), .D(n855), 
        .E(r_x_data[97]), .F(n830), .G(w_mult_3_Z[1]), .H(n854), .Y(n754) );
  scg4d1_hd U656 ( .A(n557), .B(r_add_2_B[2]), .C(w_mult_2_Z[2]), .D(n855), 
        .E(r_x_data[98]), .F(n834), .G(w_mult_3_Z[2]), .H(n854), .Y(n753) );
  scg4d1_hd U633 ( .A(n557), .B(r_add_2_B[25]), .C(w_mult_2_Z[25]), .D(n855), 
        .E(r_x_data[121]), .F(n834), .G(w_mult_3_Z[25]), .H(n854), .Y(n730) );
  scg4d1_hd U632 ( .A(n557), .B(r_add_2_B[26]), .C(w_mult_2_Z[26]), .D(n855), 
        .E(r_x_data[122]), .F(n832), .G(w_mult_3_Z[26]), .H(n854), .Y(n729) );
  scg4d1_hd U655 ( .A(n557), .B(r_add_2_B[3]), .C(w_mult_2_Z[3]), .D(n855), 
        .E(r_x_data[99]), .F(n834), .G(w_mult_3_Z[3]), .H(n854), .Y(n752) );
  scg4d1_hd U640 ( .A(n557), .B(r_add_2_B[18]), .C(w_mult_2_Z[18]), .D(n855), 
        .E(r_x_data[114]), .F(n834), .G(w_mult_3_Z[18]), .H(n854), .Y(n737) );
  scg4d1_hd U642 ( .A(n557), .B(r_add_2_B[16]), .C(w_mult_2_Z[16]), .D(n855), 
        .E(r_x_data[112]), .F(n832), .G(w_mult_3_Z[16]), .H(n854), .Y(n739) );
  scg4d1_hd U636 ( .A(n557), .B(r_add_2_B[22]), .C(w_mult_2_Z[22]), .D(n855), 
        .E(r_x_data[118]), .F(n830), .G(w_mult_3_Z[22]), .H(n854), .Y(n733) );
  scg4d1_hd U629 ( .A(n557), .B(r_add_2_B[29]), .C(w_mult_2_Z[29]), .D(n855), 
        .E(r_x_data[125]), .F(n832), .G(w_mult_3_Z[29]), .H(n854), .Y(n726) );
  scg4d1_hd U650 ( .A(n557), .B(r_add_2_B[8]), .C(w_mult_2_Z[8]), .D(n855), 
        .E(r_x_data[104]), .F(n830), .G(w_mult_3_Z[8]), .H(n854), .Y(n747) );
  scg4d1_hd U649 ( .A(n557), .B(r_add_2_B[9]), .C(w_mult_2_Z[9]), .D(n855), 
        .E(r_x_data[105]), .F(n832), .G(w_mult_3_Z[9]), .H(n854), .Y(n746) );
  scg4d1_hd U651 ( .A(n557), .B(r_add_2_B[7]), .C(w_mult_2_Z[7]), .D(n855), 
        .E(r_x_data[103]), .F(n832), .G(w_mult_3_Z[7]), .H(n854), .Y(n748) );
  scg4d1_hd U645 ( .A(n557), .B(r_add_2_B[13]), .C(w_mult_2_Z[13]), .D(n855), 
        .E(r_x_data[109]), .F(n834), .G(w_mult_3_Z[13]), .H(n854), .Y(n742) );
  scg4d1_hd U631 ( .A(n557), .B(r_add_2_B[27]), .C(w_mult_2_Z[27]), .D(n855), 
        .E(r_x_data[123]), .F(n832), .G(w_mult_3_Z[27]), .H(n854), .Y(n728) );
  scg4d1_hd U652 ( .A(n557), .B(r_add_2_B[6]), .C(w_mult_2_Z[6]), .D(n855), 
        .E(r_x_data[102]), .F(n830), .G(w_mult_3_Z[6]), .H(n854), .Y(n749) );
  scg4d1_hd U630 ( .A(n557), .B(r_add_2_B[28]), .C(w_mult_2_Z[28]), .D(n855), 
        .E(r_x_data[124]), .F(n830), .G(w_mult_3_Z[28]), .H(n854), .Y(n727) );
  scg4d1_hd U653 ( .A(n557), .B(r_add_2_B[5]), .C(w_mult_2_Z[5]), .D(n855), 
        .E(r_x_data[101]), .F(n834), .G(w_mult_3_Z[5]), .H(n854), .Y(n750) );
  scg4d1_hd U634 ( .A(n557), .B(r_add_2_B[24]), .C(w_mult_2_Z[24]), .D(n855), 
        .E(r_x_data[120]), .F(n834), .G(w_mult_3_Z[24]), .H(n854), .Y(n731) );
  scg4d1_hd U646 ( .A(n557), .B(r_add_2_B[12]), .C(w_mult_2_Z[12]), .D(n855), 
        .E(r_x_data[108]), .F(n834), .G(w_mult_3_Z[12]), .H(n854), .Y(n743) );
  scg4d1_hd U628 ( .A(n557), .B(r_add_2_B[30]), .C(w_mult_2_Z[30]), .D(n855), 
        .E(r_x_data[126]), .F(n832), .G(w_mult_3_Z[30]), .H(n854), .Y(n725) );
  fd3d1_hd r_pstate_reg_1_ ( .D(n498), .CK(i_CLK), .SN(i_RSTN), .Q(n542), .QN(
        n908) );
  fd3d1_hd r_counter_reg_0_ ( .D(n496), .CK(i_CLK), .SN(i_RSTN), .Q(n548), 
        .QN(n1040) );
  fd3d1_hd r_counter_reg_2_ ( .D(n494), .CK(i_CLK), .SN(i_RSTN), .Q(n495), 
        .QN(n1077) );
  clknd2d1_hd U844 ( .A(n1077), .B(w_add_1_Z_STB), .Y(n917) );
  clknd2d1_hd U845 ( .A(n829), .B(n962), .Y(n1076) );
  clknd2d1_hd U846 ( .A(N1396), .B(n829), .Y(n1032) );
  clknd2d1_hd U847 ( .A(n865), .B(n868), .Y(N1396) );
  clknd2d1_hd U848 ( .A(n916), .B(n1040), .Y(n1078) );
  clknd2d1_hd U849 ( .A(r_counter_1_), .B(N739), .Y(n904) );
  clknd2d1_hd U850 ( .A(n962), .B(n495), .Y(n899) );
  clknd2d1_hd U851 ( .A(n1079), .B(n901), .Y(N1401) );
  clknd2d1_hd U852 ( .A(w_add_2_Z_STB), .B(w_add_1_Z_STB), .Y(n1035) );
  clknd2d1_hd U853 ( .A(r_counter_1_), .B(n920), .Y(n1037) );
  clknd2d1_hd U854 ( .A(n1030), .B(N1401), .Y(n964) );
  clknd2d1_hd U855 ( .A(n829), .B(n1029), .Y(n1028) );
  clknd2d2_hd U856 ( .A(o_X_DATA_READY), .B(i_X_DATA_VALID), .Y(n828) );
  clknd2d1_hd U857 ( .A(n647), .B(n1029), .Y(n1033) );
  nr2ad1_hd U858 ( .A(n1079), .B(n1078), .Y(n4) );
  clknd2d1_hd U859 ( .A(n866), .B(n868), .Y(n867) );
  clknd2d4_hd U860 ( .A(n647), .B(n906), .Y(n861) );
  clknd2d1_hd U861 ( .A(n829), .B(n906), .Y(n866) );
  clknd2d1_hd U862 ( .A(r_counter_1_), .B(n1040), .Y(n960) );
  clknd2d1_hd U863 ( .A(n843), .B(i_X_DATA[31]), .Y(n1044) );
  clknd2d1_hd U864 ( .A(n849), .B(i_X_DATA[30]), .Y(n1045) );
  clknd2d1_hd U865 ( .A(n844), .B(i_X_DATA[29]), .Y(n1046) );
  clknd2d1_hd U866 ( .A(n848), .B(i_X_DATA[28]), .Y(n1047) );
  clknd2d1_hd U867 ( .A(n842), .B(i_X_DATA[27]), .Y(n1048) );
  clknd2d1_hd U868 ( .A(n846), .B(i_X_DATA[26]), .Y(n1049) );
  clknd2d1_hd U869 ( .A(n845), .B(i_X_DATA[25]), .Y(n1050) );
  clknd2d1_hd U870 ( .A(n847), .B(i_X_DATA[24]), .Y(n1051) );
  clknd2d1_hd U871 ( .A(n842), .B(i_X_DATA[23]), .Y(n1052) );
  clknd2d1_hd U872 ( .A(n848), .B(i_X_DATA[22]), .Y(n1053) );
  clknd2d1_hd U873 ( .A(n843), .B(i_X_DATA[21]), .Y(n1054) );
  clknd2d1_hd U874 ( .A(n848), .B(i_X_DATA[20]), .Y(n1055) );
  clknd2d1_hd U875 ( .A(n849), .B(i_X_DATA[19]), .Y(n1056) );
  clknd2d1_hd U876 ( .A(n844), .B(i_X_DATA[18]), .Y(n1057) );
  clknd2d1_hd U877 ( .A(n844), .B(i_X_DATA[17]), .Y(n1058) );
  clknd2d1_hd U878 ( .A(n845), .B(i_X_DATA[16]), .Y(n1059) );
  clknd2d1_hd U879 ( .A(n842), .B(i_X_DATA[15]), .Y(n1060) );
  clknd2d1_hd U880 ( .A(n846), .B(i_X_DATA[14]), .Y(n1061) );
  clknd2d1_hd U881 ( .A(n847), .B(i_X_DATA[13]), .Y(n1062) );
  clknd2d1_hd U882 ( .A(n845), .B(i_X_DATA[12]), .Y(n1063) );
  clknd2d1_hd U883 ( .A(n843), .B(i_X_DATA[11]), .Y(n1064) );
  clknd2d1_hd U884 ( .A(n847), .B(i_X_DATA[10]), .Y(n1065) );
  clknd2d1_hd U885 ( .A(n846), .B(i_X_DATA[9]), .Y(n1066) );
  clknd2d1_hd U886 ( .A(n847), .B(i_X_DATA[8]), .Y(n1067) );
  clknd2d1_hd U887 ( .A(n846), .B(i_X_DATA[7]), .Y(n1068) );
  clknd2d1_hd U888 ( .A(n847), .B(i_X_DATA[6]), .Y(n1069) );
  clknd2d1_hd U889 ( .A(n846), .B(i_X_DATA[5]), .Y(n1070) );
  clknd2d1_hd U890 ( .A(n873), .B(n895), .Y(n16) );
  clknd2d1_hd U891 ( .A(n873), .B(n893), .Y(n17) );
  clknd2d1_hd U892 ( .A(n873), .B(n892), .Y(n18) );
  clknd2d1_hd U893 ( .A(n873), .B(n891), .Y(n19) );
  clknd2d1_hd U894 ( .A(n873), .B(n890), .Y(n20) );
  clknd2d1_hd U895 ( .A(n873), .B(n889), .Y(n21) );
  clknd2d1_hd U896 ( .A(n888), .B(n857), .Y(n22) );
  clknd2d1_hd U897 ( .A(n873), .B(n887), .Y(n23) );
  clknd2d1_hd U898 ( .A(n873), .B(n886), .Y(n24) );
  clknd2d1_hd U899 ( .A(n885), .B(n857), .Y(n26) );
  clknd2d1_hd U900 ( .A(n884), .B(n872), .Y(n27) );
  clknd2d1_hd U901 ( .A(n883), .B(n872), .Y(n28) );
  clknd2d1_hd U902 ( .A(n882), .B(n872), .Y(n30) );
  clknd2d1_hd U903 ( .A(n881), .B(n857), .Y(n31) );
  clknd2d1_hd U904 ( .A(n880), .B(n857), .Y(n32) );
  clknd2d1_hd U905 ( .A(n879), .B(n872), .Y(n34) );
  clknd2d1_hd U906 ( .A(n878), .B(n872), .Y(n35) );
  clknd2d1_hd U907 ( .A(n873), .B(n877), .Y(n38) );
  clknd2d1_hd U908 ( .A(n876), .B(n857), .Y(n40) );
  clknd2d1_hd U909 ( .A(n875), .B(n872), .Y(n41) );
  clknd2d1_hd U910 ( .A(n873), .B(n874), .Y(n42) );
  clknd2d1_hd U911 ( .A(n871), .B(n872), .Y(n43) );
  clknd2d1_hd U912 ( .A(n863), .B(n857), .Y(n502) );
  clknd2d1_hd U913 ( .A(n1043), .B(n960), .Y(n961) );
  ivd2_hd U914 ( .A(n1027), .Y(n839) );
  clknd2d4_hd U915 ( .A(n829), .B(n954), .Y(n955) );
  ivd4_hd U916 ( .A(n857), .Y(n830) );
  scg10d1_hd U917 ( .A(n833), .B(o_Y_DATA[5]), .C(r_y_data[5]), .D(n843), .Y(
        n324) );
  scg10d1_hd U918 ( .A(n833), .B(o_Y_DATA[0]), .C(r_y_data[0]), .D(n846), .Y(
        n329) );
  scg10d1_hd U919 ( .A(n833), .B(r_x_data[114]), .C(r_x_data[146]), .D(n847), 
        .Y(n343) );
  scg10d1_hd U920 ( .A(n833), .B(r_x_data[116]), .C(r_x_data[148]), .D(n849), 
        .Y(n341) );
  scg10d1_hd U921 ( .A(n833), .B(r_x_data[118]), .C(r_x_data[150]), .D(n845), 
        .Y(n339) );
  scg10d1_hd U922 ( .A(n833), .B(r_x_data[119]), .C(r_x_data[151]), .D(n844), 
        .Y(n338) );
  scg10d1_hd U923 ( .A(n833), .B(r_x_data[120]), .C(r_x_data[152]), .D(n842), 
        .Y(n337) );
  scg10d1_hd U924 ( .A(n833), .B(r_x_data[126]), .C(r_x_data[158]), .D(n848), 
        .Y(n331) );
  scg10d1_hd U925 ( .A(n833), .B(r_x_data[121]), .C(r_x_data[153]), .D(n843), 
        .Y(n336) );
  scg10d1_hd U926 ( .A(n833), .B(r_x_data[122]), .C(r_x_data[154]), .D(n846), 
        .Y(n335) );
  scg10d1_hd U927 ( .A(n833), .B(r_x_data[124]), .C(r_x_data[156]), .D(n847), 
        .Y(n333) );
  scg10d1_hd U928 ( .A(n833), .B(r_x_data[123]), .C(r_x_data[155]), .D(n849), 
        .Y(n334) );
  scg10d1_hd U929 ( .A(n833), .B(o_Y_DATA[2]), .C(r_y_data[2]), .D(n845), .Y(
        n327) );
  nid8_hd U930 ( .A(n828), .Y(n833) );
  nid2_hd U931 ( .A(n573), .Y(n853) );
  ad2bd2_hd U932 ( .B(n568), .AN(n1040), .Y(n558) );
  or2d4_hd U933 ( .A(n899), .B(n918), .Y(n857) );
  nid4_hd U934 ( .A(n861), .Y(n831) );
  scg10d1_hd U935 ( .A(n833), .B(r_x_data[103]), .C(r_x_data[135]), .D(n847), 
        .Y(n354) );
  scg10d1_hd U936 ( .A(n833), .B(r_x_data[113]), .C(r_x_data[145]), .D(n849), 
        .Y(n344) );
  scg10d1_hd U937 ( .A(n833), .B(r_x_data[102]), .C(r_x_data[134]), .D(n847), 
        .Y(n355) );
  scg10d1_hd U938 ( .A(n833), .B(r_x_data[100]), .C(r_x_data[132]), .D(n846), 
        .Y(n357) );
  scg10d1_hd U939 ( .A(n833), .B(r_x_data[99]), .C(r_x_data[131]), .D(n843), 
        .Y(n358) );
  scg10d1_hd U940 ( .A(n833), .B(r_x_data[106]), .C(r_x_data[138]), .D(n846), 
        .Y(n351) );
  scg10d1_hd U941 ( .A(n833), .B(r_x_data[98]), .C(r_x_data[130]), .D(n849), 
        .Y(n359) );
  scg10d1_hd U942 ( .A(n833), .B(r_x_data[108]), .C(r_x_data[140]), .D(n843), 
        .Y(n349) );
  scg10d1_hd U943 ( .A(n833), .B(r_x_data[115]), .C(r_x_data[147]), .D(n849), 
        .Y(n342) );
  scg10d1_hd U944 ( .A(n833), .B(r_x_data[109]), .C(r_x_data[141]), .D(n849), 
        .Y(n348) );
  scg10d1_hd U945 ( .A(n833), .B(r_x_data[117]), .C(r_x_data[149]), .D(n849), 
        .Y(n340) );
  scg10d1_hd U946 ( .A(n833), .B(r_x_data[110]), .C(r_x_data[142]), .D(n843), 
        .Y(n347) );
  scg10d1_hd U947 ( .A(n833), .B(r_x_data[94]), .C(r_x_data[126]), .D(n848), 
        .Y(n363) );
  scg10d1_hd U948 ( .A(n833), .B(r_x_data[93]), .C(r_x_data[125]), .D(n842), 
        .Y(n364) );
  scg10d1_hd U949 ( .A(n833), .B(r_x_data[92]), .C(r_x_data[124]), .D(n844), 
        .Y(n365) );
  scg10d1_hd U950 ( .A(n833), .B(r_x_data[95]), .C(r_x_data[127]), .D(n845), 
        .Y(n362) );
  scg10d1_hd U951 ( .A(n833), .B(r_y_data[95]), .C(r_y_data[127]), .D(n848), 
        .Y(n203) );
  scg10d1_hd U952 ( .A(n833), .B(o_Y_DATA[20]), .C(r_y_data[20]), .D(n849), 
        .Y(n309) );
  scg10d1_hd U953 ( .A(n833), .B(o_Y_DATA[18]), .C(r_y_data[18]), .D(n849), 
        .Y(n311) );
  scg10d1_hd U954 ( .A(n833), .B(o_Y_DATA[13]), .C(r_y_data[13]), .D(n849), 
        .Y(n316) );
  scg10d1_hd U955 ( .A(n833), .B(o_Y_DATA[12]), .C(r_y_data[12]), .D(n849), 
        .Y(n317) );
  scg10d1_hd U956 ( .A(n833), .B(o_Y_DATA[9]), .C(r_y_data[9]), .D(n849), .Y(
        n320) );
  ad2d1_hd U957 ( .A(N739), .B(w_mult_3_Z_STB), .Y(n506) );
  ad4d1_hd U958 ( .A(w_add_1_Z_STB), .B(w_add_2_Z_STB), .C(w_mult_1_Z_STB), 
        .D(w_mult_2_Z_STB), .Y(N739) );
  ad2bd2_hd U959 ( .B(n920), .AN(n1028), .Y(n574) );
  ivd4_hd U960 ( .A(n857), .Y(n832) );
  ao21d2_hd U961 ( .A(n1037), .B(n1078), .C(n1032), .Y(n559) );
  nd2d4_hd U962 ( .A(N1396), .B(n647), .Y(n557) );
  nid3_hd U963 ( .A(n864), .Y(n907) );
  scg10d1_hd U964 ( .A(n851), .B(r_y_data[68]), .C(r_y_data[100]), .D(n846), 
        .Y(n230) );
  scg10d1_hd U965 ( .A(n850), .B(r_x_data[79]), .C(r_x_data[111]), .D(n843), 
        .Y(n378) );
  scg10d1_hd U966 ( .A(n851), .B(r_y_data[67]), .C(r_y_data[99]), .D(n846), 
        .Y(n231) );
  scg10d1_hd U967 ( .A(n850), .B(r_x_data[74]), .C(r_x_data[106]), .D(n842), 
        .Y(n383) );
  scg10d1_hd U968 ( .A(n851), .B(r_x_data[65]), .C(r_x_data[97]), .D(n842), 
        .Y(n392) );
  scg10d1_hd U969 ( .A(n851), .B(r_y_data[69]), .C(r_y_data[101]), .D(n846), 
        .Y(n229) );
  scg10d1_hd U970 ( .A(n851), .B(r_x_data[52]), .C(r_x_data[84]), .D(n843), 
        .Y(n405) );
  scg10d1_hd U971 ( .A(n851), .B(r_y_data[76]), .C(r_y_data[108]), .D(n846), 
        .Y(n222) );
  scg10d1_hd U972 ( .A(n850), .B(r_x_data[64]), .C(r_x_data[96]), .D(n842), 
        .Y(n393) );
  scg10d1_hd U973 ( .A(n851), .B(r_y_data[70]), .C(r_y_data[102]), .D(n846), 
        .Y(n228) );
  scg10d1_hd U974 ( .A(n851), .B(r_x_data[51]), .C(r_x_data[83]), .D(n843), 
        .Y(n406) );
  scg10d1_hd U975 ( .A(n850), .B(r_x_data[78]), .C(r_x_data[110]), .D(n842), 
        .Y(n379) );
  scg10d1_hd U976 ( .A(n850), .B(r_x_data[73]), .C(r_x_data[105]), .D(n843), 
        .Y(n384) );
  scg10d1_hd U977 ( .A(n850), .B(r_x_data[61]), .C(r_x_data[93]), .D(n842), 
        .Y(n396) );
  scg10d1_hd U978 ( .A(n851), .B(r_x_data[50]), .C(r_x_data[82]), .D(n843), 
        .Y(n407) );
  scg10d1_hd U979 ( .A(n851), .B(r_y_data[66]), .C(r_y_data[98]), .D(n846), 
        .Y(n232) );
  scg10d1_hd U980 ( .A(n850), .B(r_x_data[72]), .C(r_x_data[104]), .D(n842), 
        .Y(n385) );
  scg10d1_hd U981 ( .A(n850), .B(r_x_data[55]), .C(r_x_data[87]), .D(n842), 
        .Y(n402) );
  scg10d1_hd U982 ( .A(n851), .B(r_x_data[49]), .C(r_x_data[81]), .D(n843), 
        .Y(n408) );
  scg10d1_hd U983 ( .A(n850), .B(r_x_data[66]), .C(r_x_data[98]), .D(n842), 
        .Y(n391) );
  scg10d1_hd U984 ( .A(n851), .B(r_x_data[60]), .C(r_x_data[92]), .D(n842), 
        .Y(n397) );
  scg10d1_hd U985 ( .A(n850), .B(r_x_data[71]), .C(r_x_data[103]), .D(n843), 
        .Y(n386) );
  scg10d1_hd U986 ( .A(n851), .B(r_y_data[71]), .C(r_y_data[103]), .D(n847), 
        .Y(n227) );
  scg10d1_hd U987 ( .A(n851), .B(r_y_data[72]), .C(r_y_data[104]), .D(n846), 
        .Y(n226) );
  scg10d1_hd U988 ( .A(n850), .B(r_x_data[59]), .C(r_x_data[91]), .D(n842), 
        .Y(n398) );
  scg10d1_hd U989 ( .A(n851), .B(r_x_data[56]), .C(r_x_data[88]), .D(n842), 
        .Y(n401) );
  scg10d1_hd U990 ( .A(n850), .B(r_x_data[67]), .C(r_x_data[99]), .D(n842), 
        .Y(n390) );
  scg10d1_hd U991 ( .A(n850), .B(r_x_data[70]), .C(r_x_data[102]), .D(n842), 
        .Y(n387) );
  scg10d1_hd U992 ( .A(n850), .B(r_x_data[77]), .C(r_x_data[109]), .D(n843), 
        .Y(n380) );
  scg10d1_hd U993 ( .A(n851), .B(r_y_data[73]), .C(r_y_data[105]), .D(n847), 
        .Y(n225) );
  scg10d1_hd U994 ( .A(n851), .B(r_x_data[68]), .C(r_x_data[100]), .D(n842), 
        .Y(n389) );
  scg10d1_hd U995 ( .A(n851), .B(r_y_data[65]), .C(r_y_data[97]), .D(n846), 
        .Y(n233) );
  scg10d1_hd U996 ( .A(n850), .B(r_x_data[57]), .C(r_x_data[89]), .D(n842), 
        .Y(n400) );
  scg10d1_hd U997 ( .A(n851), .B(r_y_data[75]), .C(r_y_data[107]), .D(n847), 
        .Y(n223) );
  scg10d1_hd U998 ( .A(n851), .B(r_y_data[74]), .C(r_y_data[106]), .D(n846), 
        .Y(n224) );
  scg10d1_hd U999 ( .A(n850), .B(r_x_data[76]), .C(r_x_data[108]), .D(n842), 
        .Y(n381) );
  scg10d1_hd U1000 ( .A(n850), .B(r_x_data[125]), .C(r_x_data[157]), .D(n849), 
        .Y(n332) );
  scg10d1_hd U1001 ( .A(n851), .B(r_y_data[64]), .C(r_y_data[96]), .D(n846), 
        .Y(n234) );
  scg10d1_hd U1002 ( .A(n850), .B(r_x_data[58]), .C(r_x_data[90]), .D(n842), 
        .Y(n399) );
  scg10d1_hd U1003 ( .A(n850), .B(r_x_data[69]), .C(r_x_data[101]), .D(n842), 
        .Y(n388) );
  scg10d1_hd U1004 ( .A(n850), .B(r_x_data[75]), .C(r_x_data[107]), .D(n843), 
        .Y(n382) );
  scg10d1_hd U1005 ( .A(n851), .B(r_y_data[56]), .C(r_y_data[88]), .D(n846), 
        .Y(n242) );
  scg10d1_hd U1006 ( .A(n851), .B(r_y_data[57]), .C(r_y_data[89]), .D(n846), 
        .Y(n241) );
  scg10d1_hd U1007 ( .A(n851), .B(r_y_data[58]), .C(r_y_data[90]), .D(n846), 
        .Y(n240) );
  scg10d1_hd U1008 ( .A(n851), .B(r_y_data[59]), .C(r_y_data[91]), .D(n846), 
        .Y(n239) );
  scg10d1_hd U1009 ( .A(n851), .B(r_y_data[60]), .C(r_y_data[92]), .D(n846), 
        .Y(n238) );
  scg10d1_hd U1010 ( .A(n851), .B(r_y_data[61]), .C(r_y_data[93]), .D(n846), 
        .Y(n237) );
  scg10d1_hd U1011 ( .A(n851), .B(r_y_data[62]), .C(r_y_data[94]), .D(n846), 
        .Y(n236) );
  scg10d1_hd U1012 ( .A(n851), .B(r_y_data[63]), .C(r_y_data[95]), .D(n846), 
        .Y(n235) );
  scg10d1_hd U1013 ( .A(n850), .B(r_x_data[91]), .C(r_x_data[123]), .D(n847), 
        .Y(n366) );
  scg10d1_hd U1014 ( .A(n850), .B(r_x_data[90]), .C(r_x_data[122]), .D(n846), 
        .Y(n367) );
  scg10d1_hd U1015 ( .A(n850), .B(r_x_data[89]), .C(r_x_data[121]), .D(n843), 
        .Y(n368) );
  scg10d1_hd U1016 ( .A(n850), .B(r_x_data[88]), .C(r_x_data[120]), .D(n849), 
        .Y(n369) );
  scg10d1_hd U1017 ( .A(n851), .B(r_x_data[87]), .C(r_x_data[119]), .D(n849), 
        .Y(n370) );
  scg10d1_hd U1018 ( .A(n850), .B(r_x_data[86]), .C(r_x_data[118]), .D(n842), 
        .Y(n371) );
  scg10d1_hd U1019 ( .A(n850), .B(r_x_data[85]), .C(r_x_data[117]), .D(n843), 
        .Y(n372) );
  scg10d1_hd U1020 ( .A(n850), .B(r_x_data[84]), .C(r_x_data[116]), .D(n842), 
        .Y(n373) );
  scg10d1_hd U1021 ( .A(n850), .B(r_x_data[80]), .C(r_x_data[112]), .D(n842), 
        .Y(n377) );
  scg10d1_hd U1022 ( .A(n850), .B(r_x_data[54]), .C(r_x_data[86]), .D(n843), 
        .Y(n403) );
  scg10d1_hd U1023 ( .A(n851), .B(r_y_data[77]), .C(r_y_data[109]), .D(n847), 
        .Y(n221) );
  scg10d1_hd U1024 ( .A(n850), .B(r_x_data[53]), .C(r_x_data[85]), .D(n843), 
        .Y(n404) );
  scg10d1_hd U1025 ( .A(n850), .B(r_x_data[83]), .C(r_x_data[115]), .D(n843), 
        .Y(n374) );
  scg10d1_hd U1026 ( .A(n850), .B(r_x_data[81]), .C(r_x_data[113]), .D(n843), 
        .Y(n376) );
  scg10d1_hd U1027 ( .A(n850), .B(r_x_data[82]), .C(r_x_data[114]), .D(n842), 
        .Y(n375) );
  scg10d1_hd U1028 ( .A(n850), .B(r_x_data[62]), .C(r_x_data[94]), .D(n842), 
        .Y(n395) );
  scg10d1_hd U1029 ( .A(n850), .B(r_x_data[63]), .C(r_x_data[95]), .D(n842), 
        .Y(n394) );
  scg10d1_hd U1030 ( .A(n850), .B(r_x_data[107]), .C(r_x_data[139]), .D(n842), 
        .Y(n350) );
  scg10d1_hd U1031 ( .A(n850), .B(o_Y_DATA[31]), .C(r_y_data[31]), .D(n845), 
        .Y(n500) );
  scg10d1_hd U1032 ( .A(n833), .B(r_y_data[32]), .C(r_y_data[64]), .D(n849), 
        .Y(n266) );
  scg10d1_hd U1033 ( .A(n833), .B(r_y_data[34]), .C(r_y_data[66]), .D(n847), 
        .Y(n264) );
  scg10d1_hd U1034 ( .A(n850), .B(r_x_data[105]), .C(r_x_data[137]), .D(n844), 
        .Y(n352) );
  scg10d1_hd U1035 ( .A(n833), .B(r_y_data[35]), .C(r_y_data[67]), .D(n848), 
        .Y(n263) );
  scg10d1_hd U1036 ( .A(n833), .B(r_y_data[55]), .C(r_y_data[87]), .D(n846), 
        .Y(n243) );
  scg10d1_hd U1037 ( .A(n833), .B(r_y_data[54]), .C(r_y_data[86]), .D(n847), 
        .Y(n244) );
  scg10d1_hd U1038 ( .A(n850), .B(r_x_data[0]), .C(r_x_data[32]), .D(n845), 
        .Y(n457) );
  scg10d1_hd U1039 ( .A(n833), .B(r_y_data[36]), .C(r_y_data[68]), .D(n846), 
        .Y(n262) );
  scg10d1_hd U1040 ( .A(n850), .B(r_x_data[1]), .C(r_x_data[33]), .D(n845), 
        .Y(n456) );
  scg10d1_hd U1041 ( .A(n833), .B(r_y_data[37]), .C(r_y_data[69]), .D(n848), 
        .Y(n261) );
  scg10d1_hd U1042 ( .A(n850), .B(r_x_data[104]), .C(r_x_data[136]), .D(n845), 
        .Y(n353) );
  scg10d1_hd U1043 ( .A(n833), .B(r_y_data[33]), .C(r_y_data[65]), .D(n848), 
        .Y(n265) );
  scg10d1_hd U1044 ( .A(n833), .B(r_y_data[38]), .C(r_y_data[70]), .D(n843), 
        .Y(n260) );
  scg10d1_hd U1045 ( .A(n833), .B(r_y_data[39]), .C(r_y_data[71]), .D(n847), 
        .Y(n259) );
  scg10d1_hd U1046 ( .A(n833), .B(r_y_data[40]), .C(r_y_data[72]), .D(n847), 
        .Y(n258) );
  scg10d1_hd U1047 ( .A(n833), .B(r_y_data[53]), .C(r_y_data[85]), .D(n847), 
        .Y(n245) );
  scg10d1_hd U1048 ( .A(n833), .B(r_y_data[52]), .C(r_y_data[84]), .D(n847), 
        .Y(n246) );
  scg10d1_hd U1049 ( .A(n833), .B(r_y_data[51]), .C(r_y_data[83]), .D(n847), 
        .Y(n247) );
  scg10d1_hd U1050 ( .A(n833), .B(r_y_data[41]), .C(r_y_data[73]), .D(n847), 
        .Y(n257) );
  scg10d1_hd U1051 ( .A(n850), .B(r_x_data[101]), .C(r_x_data[133]), .D(n849), 
        .Y(n356) );
  scg10d1_hd U1052 ( .A(n833), .B(r_y_data[42]), .C(r_y_data[74]), .D(n847), 
        .Y(n256) );
  scg10d1_hd U1053 ( .A(n833), .B(r_y_data[50]), .C(r_y_data[82]), .D(n847), 
        .Y(n248) );
  scg10d1_hd U1054 ( .A(n833), .B(r_y_data[43]), .C(r_y_data[75]), .D(n847), 
        .Y(n255) );
  scg10d1_hd U1055 ( .A(n833), .B(r_y_data[44]), .C(r_y_data[76]), .D(n847), 
        .Y(n254) );
  scg10d1_hd U1056 ( .A(n833), .B(r_y_data[49]), .C(r_y_data[81]), .D(n847), 
        .Y(n249) );
  scg10d1_hd U1057 ( .A(n850), .B(r_x_data[97]), .C(r_x_data[129]), .D(n849), 
        .Y(n360) );
  scg10d1_hd U1058 ( .A(n833), .B(r_y_data[45]), .C(r_y_data[77]), .D(n847), 
        .Y(n253) );
  scg10d1_hd U1059 ( .A(n850), .B(r_x_data[96]), .C(r_x_data[128]), .D(n849), 
        .Y(n361) );
  scg10d1_hd U1060 ( .A(n833), .B(r_y_data[48]), .C(r_y_data[80]), .D(n847), 
        .Y(n250) );
  scg10d1_hd U1061 ( .A(n833), .B(r_y_data[47]), .C(r_y_data[79]), .D(n847), 
        .Y(n251) );
  scg10d1_hd U1062 ( .A(n833), .B(r_y_data[46]), .C(r_y_data[78]), .D(n847), 
        .Y(n252) );
  scg10d1_hd U1063 ( .A(n850), .B(r_x_data[127]), .C(r_x_data[159]), .D(n847), 
        .Y(n330) );
  scg10d1_hd U1064 ( .A(n850), .B(r_y_data[78]), .C(r_y_data[110]), .D(n846), 
        .Y(n220) );
  scg10d1_hd U1065 ( .A(n850), .B(r_y_data[79]), .C(r_y_data[111]), .D(n847), 
        .Y(n219) );
  scg10d1_hd U1066 ( .A(n850), .B(r_y_data[80]), .C(r_y_data[112]), .D(n846), 
        .Y(n218) );
  scg10d1_hd U1067 ( .A(n850), .B(r_y_data[81]), .C(r_y_data[113]), .D(n847), 
        .Y(n217) );
  scg10d1_hd U1068 ( .A(n850), .B(r_y_data[82]), .C(r_y_data[114]), .D(n846), 
        .Y(n216) );
  scg10d1_hd U1069 ( .A(n850), .B(r_y_data[83]), .C(r_y_data[115]), .D(n847), 
        .Y(n215) );
  scg10d1_hd U1070 ( .A(n850), .B(r_y_data[84]), .C(r_y_data[116]), .D(n846), 
        .Y(n214) );
  scg10d1_hd U1071 ( .A(n850), .B(r_y_data[85]), .C(r_y_data[117]), .D(n847), 
        .Y(n213) );
  scg10d1_hd U1072 ( .A(n850), .B(r_y_data[86]), .C(r_y_data[118]), .D(n846), 
        .Y(n212) );
  scg10d1_hd U1073 ( .A(n850), .B(r_y_data[87]), .C(r_y_data[119]), .D(n845), 
        .Y(n211) );
  scg10d1_hd U1074 ( .A(n850), .B(r_y_data[88]), .C(r_y_data[120]), .D(n845), 
        .Y(n210) );
  scg10d1_hd U1075 ( .A(n850), .B(r_y_data[89]), .C(r_y_data[121]), .D(n845), 
        .Y(n209) );
  scg10d1_hd U1076 ( .A(n850), .B(r_y_data[90]), .C(r_y_data[122]), .D(n845), 
        .Y(n208) );
  scg10d1_hd U1077 ( .A(n850), .B(r_y_data[91]), .C(r_y_data[123]), .D(n845), 
        .Y(n207) );
  scg10d1_hd U1078 ( .A(n850), .B(r_y_data[92]), .C(r_y_data[124]), .D(n845), 
        .Y(n206) );
  scg10d1_hd U1079 ( .A(n850), .B(r_y_data[93]), .C(r_y_data[125]), .D(n845), 
        .Y(n205) );
  scg10d1_hd U1080 ( .A(n833), .B(r_y_data[94]), .C(r_y_data[126]), .D(n848), 
        .Y(n204) );
  scg10d1_hd U1081 ( .A(n850), .B(r_x_data[32]), .C(r_x_data[64]), .D(n844), 
        .Y(n425) );
  scg10d1_hd U1082 ( .A(n850), .B(r_x_data[33]), .C(r_x_data[65]), .D(n844), 
        .Y(n424) );
  scg10d1_hd U1083 ( .A(n850), .B(r_x_data[34]), .C(r_x_data[66]), .D(n844), 
        .Y(n423) );
  scg10d1_hd U1084 ( .A(n850), .B(r_x_data[36]), .C(r_x_data[68]), .D(n844), 
        .Y(n421) );
  scg10d1_hd U1085 ( .A(n850), .B(r_x_data[37]), .C(r_x_data[69]), .D(n844), 
        .Y(n420) );
  scg10d1_hd U1086 ( .A(n850), .B(r_x_data[38]), .C(r_x_data[70]), .D(n844), 
        .Y(n419) );
  scg10d1_hd U1087 ( .A(n850), .B(r_x_data[39]), .C(r_x_data[71]), .D(n844), 
        .Y(n418) );
  scg10d1_hd U1088 ( .A(n850), .B(r_x_data[40]), .C(r_x_data[72]), .D(n843), 
        .Y(n417) );
  scg10d1_hd U1089 ( .A(n850), .B(r_x_data[41]), .C(r_x_data[73]), .D(n843), 
        .Y(n416) );
  scg10d1_hd U1090 ( .A(n850), .B(r_x_data[42]), .C(r_x_data[74]), .D(n843), 
        .Y(n415) );
  scg10d1_hd U1091 ( .A(n850), .B(r_x_data[43]), .C(r_x_data[75]), .D(n843), 
        .Y(n414) );
  scg10d1_hd U1092 ( .A(n850), .B(r_x_data[44]), .C(r_x_data[76]), .D(n843), 
        .Y(n413) );
  scg10d1_hd U1093 ( .A(n850), .B(r_x_data[45]), .C(r_x_data[77]), .D(n843), 
        .Y(n412) );
  scg10d1_hd U1094 ( .A(n850), .B(r_x_data[46]), .C(r_x_data[78]), .D(n843), 
        .Y(n411) );
  scg10d1_hd U1095 ( .A(n850), .B(r_x_data[112]), .C(r_x_data[144]), .D(n846), 
        .Y(n345) );
  scg10d1_hd U1096 ( .A(n850), .B(r_x_data[47]), .C(r_x_data[79]), .D(n843), 
        .Y(n410) );
  scg10d1_hd U1097 ( .A(n850), .B(r_x_data[48]), .C(r_x_data[80]), .D(n843), 
        .Y(n409) );
  scg10d1_hd U1098 ( .A(n850), .B(r_x_data[111]), .C(r_x_data[143]), .D(n849), 
        .Y(n346) );
  scg10d1_hd U1099 ( .A(n833), .B(r_y_data[12]), .C(r_y_data[44]), .D(n842), 
        .Y(n286) );
  scg10d1_hd U1100 ( .A(n850), .B(r_x_data[30]), .C(r_x_data[62]), .D(n844), 
        .Y(n427) );
  scg10d1_hd U1101 ( .A(n833), .B(r_y_data[11]), .C(r_y_data[43]), .D(n844), 
        .Y(n287) );
  scg10d1_hd U1102 ( .A(n850), .B(r_x_data[29]), .C(r_x_data[61]), .D(n844), 
        .Y(n428) );
  scg10d1_hd U1103 ( .A(n833), .B(r_y_data[13]), .C(r_y_data[45]), .D(n845), 
        .Y(n285) );
  scg10d1_hd U1104 ( .A(n850), .B(r_x_data[28]), .C(r_x_data[60]), .D(n844), 
        .Y(n429) );
  scg10d1_hd U1105 ( .A(n833), .B(r_y_data[10]), .C(r_y_data[42]), .D(n849), 
        .Y(n288) );
  scg10d1_hd U1106 ( .A(n850), .B(r_x_data[27]), .C(r_x_data[59]), .D(n844), 
        .Y(n430) );
  scg10d1_hd U1107 ( .A(n850), .B(o_Y_DATA[1]), .C(r_y_data[1]), .D(n843), .Y(
        n328) );
  scg10d1_hd U1108 ( .A(n850), .B(r_x_data[26]), .C(r_x_data[58]), .D(n844), 
        .Y(n431) );
  scg10d1_hd U1109 ( .A(n833), .B(r_y_data[9]), .C(r_y_data[41]), .D(n847), 
        .Y(n289) );
  scg10d1_hd U1110 ( .A(n833), .B(r_y_data[14]), .C(r_y_data[46]), .D(n846), 
        .Y(n284) );
  scg10d1_hd U1111 ( .A(n850), .B(r_x_data[25]), .C(r_x_data[57]), .D(n844), 
        .Y(n432) );
  scg10d1_hd U1112 ( .A(n833), .B(r_y_data[8]), .C(r_y_data[40]), .D(n843), 
        .Y(n290) );
  scg10d1_hd U1113 ( .A(n833), .B(r_y_data[15]), .C(r_y_data[47]), .D(n848), 
        .Y(n283) );
  scg10d1_hd U1114 ( .A(n850), .B(r_x_data[24]), .C(r_x_data[56]), .D(n844), 
        .Y(n433) );
  scg10d1_hd U1115 ( .A(n850), .B(o_Y_DATA[3]), .C(r_y_data[3]), .D(n848), .Y(
        n326) );
  scg10d1_hd U1116 ( .A(n850), .B(r_x_data[23]), .C(r_x_data[55]), .D(n845), 
        .Y(n434) );
  scg10d1_hd U1117 ( .A(n833), .B(r_y_data[7]), .C(r_y_data[39]), .D(n848), 
        .Y(n291) );
  scg10d1_hd U1118 ( .A(n833), .B(r_y_data[16]), .C(r_y_data[48]), .D(n842), 
        .Y(n282) );
  scg10d1_hd U1119 ( .A(n833), .B(r_y_data[17]), .C(r_y_data[49]), .D(n844), 
        .Y(n281) );
  scg10d1_hd U1120 ( .A(n833), .B(r_y_data[6]), .C(r_y_data[38]), .D(n848), 
        .Y(n292) );
  scg10d1_hd U1121 ( .A(n850), .B(r_x_data[22]), .C(r_x_data[54]), .D(n844), 
        .Y(n435) );
  scg10d1_hd U1122 ( .A(n850), .B(o_Y_DATA[4]), .C(r_y_data[4]), .D(n842), .Y(
        n325) );
  scg10d1_hd U1123 ( .A(n833), .B(r_y_data[18]), .C(r_y_data[50]), .D(n845), 
        .Y(n280) );
  scg10d1_hd U1124 ( .A(n833), .B(r_y_data[5]), .C(r_y_data[37]), .D(n848), 
        .Y(n293) );
  scg10d1_hd U1125 ( .A(n850), .B(r_x_data[21]), .C(r_x_data[53]), .D(n845), 
        .Y(n436) );
  scg10d1_hd U1126 ( .A(n833), .B(r_y_data[4]), .C(r_y_data[36]), .D(n848), 
        .Y(n294) );
  scg10d1_hd U1127 ( .A(n833), .B(r_y_data[19]), .C(r_y_data[51]), .D(n849), 
        .Y(n279) );
  scg10d1_hd U1128 ( .A(n850), .B(r_x_data[20]), .C(r_x_data[52]), .D(n844), 
        .Y(n437) );
  scg10d1_hd U1129 ( .A(n850), .B(o_Y_DATA[6]), .C(r_y_data[6]), .D(n844), .Y(
        n323) );
  scg10d1_hd U1130 ( .A(n833), .B(r_y_data[3]), .C(r_y_data[35]), .D(n848), 
        .Y(n295) );
  scg10d1_hd U1131 ( .A(n833), .B(r_y_data[20]), .C(r_y_data[52]), .D(n847), 
        .Y(n278) );
  scg10d1_hd U1132 ( .A(n833), .B(r_y_data[2]), .C(r_y_data[34]), .D(n848), 
        .Y(n296) );
  scg10d1_hd U1133 ( .A(n850), .B(r_x_data[19]), .C(r_x_data[51]), .D(n845), 
        .Y(n438) );
  scg10d1_hd U1134 ( .A(n850), .B(o_Y_DATA[7]), .C(r_y_data[7]), .D(n849), .Y(
        n322) );
  scg10d1_hd U1135 ( .A(n833), .B(r_y_data[21]), .C(r_y_data[53]), .D(n846), 
        .Y(n277) );
  scg10d1_hd U1136 ( .A(n833), .B(r_y_data[1]), .C(r_y_data[33]), .D(n848), 
        .Y(n297) );
  scg10d1_hd U1137 ( .A(n850), .B(r_x_data[18]), .C(r_x_data[50]), .D(n844), 
        .Y(n439) );
  scg10d1_hd U1138 ( .A(n850), .B(o_Y_DATA[8]), .C(r_y_data[8]), .D(n849), .Y(
        n321) );
  scg10d1_hd U1139 ( .A(n833), .B(r_y_data[0]), .C(r_y_data[32]), .D(n848), 
        .Y(n298) );
  scg10d1_hd U1140 ( .A(n850), .B(r_x_data[17]), .C(r_x_data[49]), .D(n845), 
        .Y(n440) );
  scg10d1_hd U1141 ( .A(n833), .B(r_y_data[22]), .C(r_y_data[54]), .D(n843), 
        .Y(n276) );
  scg10d1_hd U1142 ( .A(n850), .B(r_x_data[16]), .C(r_x_data[48]), .D(n844), 
        .Y(n441) );
  scg10d1_hd U1143 ( .A(n833), .B(o_Y_DATA[30]), .C(r_y_data[30]), .D(n848), 
        .Y(n299) );
  scg10d1_hd U1144 ( .A(n850), .B(r_x_data[15]), .C(r_x_data[47]), .D(n845), 
        .Y(n442) );
  scg10d1_hd U1145 ( .A(n850), .B(r_x_data[14]), .C(r_x_data[46]), .D(n844), 
        .Y(n443) );
  scg10d1_hd U1146 ( .A(n833), .B(r_y_data[23]), .C(r_y_data[55]), .D(n848), 
        .Y(n275) );
  scg10d1_hd U1147 ( .A(n833), .B(o_Y_DATA[29]), .C(r_y_data[29]), .D(n848), 
        .Y(n300) );
  scg10d1_hd U1148 ( .A(n850), .B(r_x_data[13]), .C(r_x_data[45]), .D(n845), 
        .Y(n444) );
  scg10d1_hd U1149 ( .A(n850), .B(o_Y_DATA[10]), .C(r_y_data[10]), .D(n849), 
        .Y(n319) );
  scg10d1_hd U1150 ( .A(n833), .B(o_Y_DATA[28]), .C(r_y_data[28]), .D(n848), 
        .Y(n301) );
  scg10d1_hd U1151 ( .A(n850), .B(r_x_data[12]), .C(r_x_data[44]), .D(n844), 
        .Y(n445) );
  scg10d1_hd U1152 ( .A(n833), .B(o_Y_DATA[27]), .C(r_y_data[27]), .D(n848), 
        .Y(n302) );
  scg10d1_hd U1153 ( .A(n833), .B(r_y_data[24]), .C(r_y_data[56]), .D(n848), 
        .Y(n274) );
  scg10d1_hd U1154 ( .A(n833), .B(r_y_data[31]), .C(r_y_data[63]), .D(n848), 
        .Y(n267) );
  scg10d1_hd U1155 ( .A(n850), .B(o_Y_DATA[11]), .C(r_y_data[11]), .D(n849), 
        .Y(n318) );
  scg10d1_hd U1156 ( .A(n850), .B(o_Y_DATA[16]), .C(r_y_data[16]), .D(n849), 
        .Y(n313) );
  scg10d1_hd U1157 ( .A(n833), .B(r_y_data[25]), .C(r_y_data[57]), .D(n848), 
        .Y(n273) );
  scg10d1_hd U1158 ( .A(n850), .B(r_x_data[35]), .C(r_x_data[67]), .D(n844), 
        .Y(n422) );
  scg10d1_hd U1159 ( .A(n850), .B(r_x_data[11]), .C(r_x_data[43]), .D(n845), 
        .Y(n446) );
  scg10d1_hd U1160 ( .A(n833), .B(r_y_data[30]), .C(r_y_data[62]), .D(n842), 
        .Y(n268) );
  scg10d1_hd U1161 ( .A(n828), .B(o_Y_DATA[19]), .C(r_y_data[19]), .D(n849), 
        .Y(n310) );
  scg10d1_hd U1162 ( .A(n850), .B(o_Y_DATA[21]), .C(r_y_data[21]), .D(n849), 
        .Y(n308) );
  scg10d1_hd U1163 ( .A(n833), .B(r_y_data[29]), .C(r_y_data[61]), .D(n848), 
        .Y(n269) );
  scg10d1_hd U1164 ( .A(n850), .B(r_x_data[2]), .C(r_x_data[34]), .D(n845), 
        .Y(n455) );
  scg10d1_hd U1165 ( .A(n850), .B(r_x_data[10]), .C(r_x_data[42]), .D(n844), 
        .Y(n447) );
  scg10d1_hd U1166 ( .A(n850), .B(o_Y_DATA[17]), .C(r_y_data[17]), .D(n849), 
        .Y(n312) );
  scg10d1_hd U1167 ( .A(n833), .B(o_Y_DATA[26]), .C(r_y_data[26]), .D(n848), 
        .Y(n303) );
  scg10d1_hd U1168 ( .A(n850), .B(r_x_data[6]), .C(r_x_data[38]), .D(n845), 
        .Y(n451) );
  scg10d1_hd U1169 ( .A(n833), .B(o_Y_DATA[24]), .C(r_y_data[24]), .D(n848), 
        .Y(n305) );
  scg10d1_hd U1170 ( .A(n833), .B(r_y_data[26]), .C(r_y_data[58]), .D(n844), 
        .Y(n272) );
  scg10d1_hd U1171 ( .A(n850), .B(r_x_data[7]), .C(r_x_data[39]), .D(n845), 
        .Y(n450) );
  scg10d1_hd U1172 ( .A(n833), .B(r_y_data[28]), .C(r_y_data[60]), .D(n845), 
        .Y(n270) );
  scg10d1_hd U1173 ( .A(n850), .B(r_x_data[8]), .C(r_x_data[40]), .D(n844), 
        .Y(n449) );
  scg10d1_hd U1174 ( .A(n833), .B(o_Y_DATA[23]), .C(r_y_data[23]), .D(n848), 
        .Y(n306) );
  scg10d1_hd U1175 ( .A(n850), .B(r_x_data[4]), .C(r_x_data[36]), .D(n845), 
        .Y(n453) );
  scg10d1_hd U1176 ( .A(n850), .B(r_x_data[3]), .C(r_x_data[35]), .D(n845), 
        .Y(n454) );
  scg10d1_hd U1177 ( .A(n850), .B(r_x_data[5]), .C(r_x_data[37]), .D(n845), 
        .Y(n452) );
  scg10d1_hd U1178 ( .A(n828), .B(o_Y_DATA[14]), .C(r_y_data[14]), .D(n849), 
        .Y(n315) );
  scg10d1_hd U1179 ( .A(n833), .B(o_Y_DATA[22]), .C(r_y_data[22]), .D(n849), 
        .Y(n307) );
  scg10d1_hd U1180 ( .A(n850), .B(r_x_data[31]), .C(r_x_data[63]), .D(n844), 
        .Y(n426) );
  scg10d1_hd U1181 ( .A(n833), .B(o_Y_DATA[25]), .C(r_y_data[25]), .D(n848), 
        .Y(n304) );
  scg10d1_hd U1182 ( .A(n850), .B(o_Y_DATA[15]), .C(r_y_data[15]), .D(n849), 
        .Y(n314) );
  scg10d1_hd U1183 ( .A(n850), .B(r_x_data[9]), .C(r_x_data[41]), .D(n845), 
        .Y(n448) );
  scg10d1_hd U1184 ( .A(n833), .B(r_y_data[27]), .C(r_y_data[59]), .D(n848), 
        .Y(n271) );
  or4d1_hd U1185 ( .A(n1079), .B(n1077), .C(n1040), .D(n904), .Y(n868) );
  nid6_hd U1186 ( .A(n828), .Y(n850) );
  clknd2d1_hd U1187 ( .A(n849), .B(i_X_DATA[2]), .Y(n1073) );
  clknd2d1_hd U1188 ( .A(n844), .B(i_X_DATA[0]), .Y(n1075) );
  clknd2d1_hd U1189 ( .A(n845), .B(i_X_DATA[1]), .Y(n1074) );
  clknd2d1_hd U1190 ( .A(n842), .B(i_X_DATA[3]), .Y(n1072) );
  clknd2d1_hd U1191 ( .A(n848), .B(i_X_DATA[4]), .Y(n1071) );
  nr2ad1_hd U1192 ( .A(n830), .B(n862), .Y(n873) );
  ivd1_hd U1193 ( .A(n906), .Y(n865) );
  nid2_hd U1194 ( .A(n1034), .Y(n841) );
  ivd1_hd U1195 ( .A(n839), .Y(n836) );
  ivd1_hd U1196 ( .A(n1079), .Y(n829) );
  nid2_hd U1197 ( .A(n850), .Y(n851) );
  nid2_hd U1198 ( .A(n954), .Y(n835) );
  nid2_hd U1199 ( .A(n568), .Y(n854) );
  nid2_hd U1200 ( .A(n567), .Y(n855) );
  nid2_hd U1201 ( .A(n559), .Y(n856) );
  ivd1_hd U1202 ( .A(n839), .Y(n837) );
  ivd1_hd U1203 ( .A(n839), .Y(n838) );
  ivd1_hd U1204 ( .A(n5), .Y(n918) );
  nr2d1_hd U1205 ( .A(n902), .B(n900), .Y(n5) );
  ivd1_hd U1206 ( .A(n659), .Y(n900) );
  nr2bd1_hd U1207 ( .AN(w_mult_3_AB_ACK), .B(n903), .Y(n659) );
  nid2_hd U1208 ( .A(n574), .Y(n852) );
  nd2bd1_hd U1209 ( .AN(N1396), .B(n915), .Y(n1029) );
  ivd1_hd U1210 ( .A(n870), .Y(n902) );
  nr2bd1_hd U1211 ( .AN(r_pstate_0_), .B(n908), .Y(n870) );
  nd2d1_hd U1212 ( .A(n908), .B(n909), .Y(n1079) );
  ivd1_hd U1213 ( .A(N1401), .Y(n963) );
  oa22d1_hd U1214 ( .A(n1078), .B(n918), .C(n917), .D(n1076), .Y(n954) );
  nd2d1_hd U1215 ( .A(n906), .B(n7), .Y(n872) );
  nr2d1_hd U1216 ( .A(n956), .B(n1032), .Y(n568) );
  ao21d1_hd U1217 ( .A(n1037), .B(n1078), .C(n1028), .Y(n1034) );
  nid4_hd U1218 ( .A(n1033), .Y(n840) );
  oa21d1_hd U1219 ( .A(n900), .B(n899), .C(n870), .Y(n647) );
  nr2d1_hd U1220 ( .A(r_counter_1_), .B(n1040), .Y(n962) );
  nr2d1_hd U1221 ( .A(n1028), .B(n1078), .Y(n573) );
  nd2bd1_hd U1222 ( .AN(n1028), .B(n1042), .Y(n1027) );
  nr2d1_hd U1223 ( .A(n1077), .B(n960), .Y(n1042) );
  scg22d2_hd U1224 ( .A(n506), .B(n905), .C(n1079), .D(n902), .Y(n906) );
  ivd1_hd U1225 ( .A(r_pstate_0_), .Y(n909) );
  scg6d1_hd U1226 ( .A(r_add_1_Z_ACK), .B(n957), .C(n958), .Y(n793) );
  ivd1_hd U1227 ( .A(n1030), .Y(n957) );
  ivd2_hd U1228 ( .A(n833), .Y(n844) );
  ivd2_hd U1229 ( .A(n833), .Y(n845) );
  ivd2_hd U1230 ( .A(n833), .Y(n849) );
  ivd2_hd U1231 ( .A(n833), .Y(n848) );
  ivd2_hd U1232 ( .A(n833), .Y(n847) );
  ivd2_hd U1233 ( .A(n833), .Y(n846) );
  ivd2_hd U1234 ( .A(n833), .Y(n843) );
  ivd2_hd U1235 ( .A(n833), .Y(n842) );
  nd2d1_hd U1236 ( .A(n896), .B(n906), .Y(n894) );
  nd2d1_hd U1237 ( .A(n898), .B(n896), .Y(n860) );
  nr2d1_hd U1238 ( .A(n959), .B(n958), .Y(n1041) );
  clknd2d4_hd U1239 ( .A(n898), .B(n647), .Y(n858) );
  ivd1_hd U1240 ( .A(n897), .Y(n898) );
  ad2bd2_hd U1241 ( .B(n4), .AN(n865), .Y(n864) );
  ivd4_hd U1242 ( .A(n872), .Y(n862) );
  nr2d1_hd U1243 ( .A(n1077), .B(n1076), .Y(n7) );
  ivd4_hd U1244 ( .A(n857), .Y(n834) );
  ivd1_hd U1245 ( .A(w_add_1_Z[10]), .Y(n986) );
  ivd1_hd U1246 ( .A(w_add_1_Z[11]), .Y(n988) );
  ivd1_hd U1247 ( .A(w_add_1_Z[12]), .Y(n990) );
  ivd1_hd U1248 ( .A(n916), .Y(n956) );
  ivd1_hd U1249 ( .A(w_add_1_Z[15]), .Y(n996) );
  ivd1_hd U1250 ( .A(w_add_1_Z[14]), .Y(n994) );
  ivd1_hd U1251 ( .A(w_add_1_Z[17]), .Y(n1000) );
  ivd1_hd U1252 ( .A(w_add_1_Z[16]), .Y(n998) );
  ivd1_hd U1253 ( .A(w_add_1_Z[13]), .Y(n992) );
  ivd1_hd U1254 ( .A(w_add_1_Z[18]), .Y(n1002) );
  ivd1_hd U1255 ( .A(w_add_1_Z[19]), .Y(n1004) );
  ivd1_hd U1256 ( .A(w_add_1_Z[24]), .Y(n1014) );
  ivd1_hd U1257 ( .A(w_add_1_Z[25]), .Y(n1016) );
  ivd1_hd U1258 ( .A(w_add_1_Z[23]), .Y(n1012) );
  ivd1_hd U1259 ( .A(w_add_1_Z[21]), .Y(n1008) );
  ivd1_hd U1260 ( .A(w_add_1_Z[22]), .Y(n1010) );
  ivd1_hd U1261 ( .A(w_add_1_Z[28]), .Y(n1022) );
  ivd1_hd U1262 ( .A(w_add_1_Z[29]), .Y(n1024) );
  ivd1_hd U1263 ( .A(w_add_1_Z[26]), .Y(n1018) );
  ivd1_hd U1264 ( .A(w_add_1_Z[27]), .Y(n1020) );
  ivd1_hd U1265 ( .A(w_add_1_Z[20]), .Y(n1006) );
  ivd1_hd U1266 ( .A(w_add_1_Z[9]), .Y(n984) );
  ivd1_hd U1267 ( .A(w_add_1_Z[30]), .Y(n1026) );
  ivd1_hd U1268 ( .A(w_add_1_Z[8]), .Y(n982) );
  ivd1_hd U1269 ( .A(w_add_1_Z[6]), .Y(n978) );
  ivd1_hd U1270 ( .A(w_add_1_Z[7]), .Y(n980) );
  ivd1_hd U1271 ( .A(w_add_1_Z[5]), .Y(n976) );
  ivd1_hd U1272 ( .A(w_add_1_Z[0]), .Y(n966) );
  ivd1_hd U1273 ( .A(w_add_1_Z[2]), .Y(n970) );
  ivd1_hd U1274 ( .A(w_add_1_Z[3]), .Y(n972) );
  ivd1_hd U1275 ( .A(w_add_1_Z[31]), .Y(n922) );
  ivd1_hd U1276 ( .A(w_add_1_Z[1]), .Y(n968) );
  nd4d1_hd U1277 ( .A(w_add_1_AB_ACK), .B(w_add_2_AB_ACK), .C(w_mult_1_AB_ACK), 
        .D(w_mult_2_AB_ACK), .Y(n903) );
  nr2d1_hd U1278 ( .A(n1077), .B(n1040), .Y(n920) );
  nr2d1_hd U1279 ( .A(r_counter_1_), .B(n1077), .Y(n916) );
  ivd1_hd U1280 ( .A(w_add_1_Z[4]), .Y(n974) );
  nr2d1_hd U1281 ( .A(n908), .B(n909), .Y(n1030) );
  nd2d1_hd U1282 ( .A(n1079), .B(n857), .Y(n896) );
  nr2d4_hd U1283 ( .A(n1079), .B(n897), .Y(n859) );
  nr2d1_hd U1284 ( .A(r_pstate_0_), .B(n908), .Y(n959) );
  nr2d1_hd U1285 ( .A(n1037), .B(n1032), .Y(n567) );
  nr2d1_hd U1286 ( .A(n1077), .B(r_counter_1_), .Y(n905) );
  scg2d1_hd U1287 ( .A(w_mult_1_Z[30]), .B(n907), .C(r_mult_1_A[30]), .D(n831), 
        .Y(n15) );
  scg2d1_hd U1288 ( .A(w_mult_1_Z[12]), .B(n864), .C(r_mult_1_A[12]), .D(n831), 
        .Y(n33) );
  scg2d1_hd U1289 ( .A(w_mult_1_Z[31]), .B(n864), .C(r_mult_1_A[31]), .D(n831), 
        .Y(n14) );
  scg14d1_hd U1290 ( .A(r_mult_3_A[29]), .B(n858), .C(n860), .Y(n79) );
  scg14d1_hd U1291 ( .A(r_mult_3_A[28]), .B(n858), .C(n860), .Y(n80) );
  scg14d1_hd U1292 ( .A(r_mult_3_A[27]), .B(n858), .C(n860), .Y(n81) );
  scg14d1_hd U1293 ( .A(r_mult_3_A[26]), .B(n858), .C(n860), .Y(n82) );
  scg14d1_hd U1294 ( .A(r_mult_3_A[25]), .B(n858), .C(n860), .Y(n83) );
  scg14d1_hd U1295 ( .A(r_mult_3_A[17]), .B(n858), .C(n860), .Y(n91) );
  scg14d1_hd U1296 ( .A(r_mult_3_A[12]), .B(n858), .C(n860), .Y(n96) );
  scg14d1_hd U1297 ( .A(r_mult_3_A[7]), .B(n858), .C(n860), .Y(n101) );
  scg14d1_hd U1298 ( .A(r_mult_3_A[5]), .B(n858), .C(n860), .Y(n103) );
  scg14d1_hd U1299 ( .A(r_mult_3_A[4]), .B(n858), .C(n860), .Y(n104) );
  scg14d1_hd U1300 ( .A(r_mult_3_A[3]), .B(n858), .C(n860), .Y(n105) );
  scg2d1_hd U1301 ( .A(w_mult_1_Z[9]), .B(n907), .C(r_mult_1_A[9]), .D(n861), 
        .Y(n36) );
  scg2d1_hd U1302 ( .A(w_mult_1_Z[20]), .B(n907), .C(r_mult_1_A[20]), .D(n861), 
        .Y(n25) );
  scg2d1_hd U1303 ( .A(w_mult_1_Z[16]), .B(n864), .C(r_mult_1_A[16]), .D(n861), 
        .Y(n29) );
  scg2d1_hd U1304 ( .A(w_mult_1_Z[8]), .B(n907), .C(r_mult_1_A[8]), .D(n861), 
        .Y(n37) );
  scg2d1_hd U1305 ( .A(w_mult_1_Z[6]), .B(n864), .C(r_mult_1_A[6]), .D(n861), 
        .Y(n39) );
  scg2d1_hd U1306 ( .A(w_mult_1_Z[1]), .B(n864), .C(r_mult_1_A[1]), .D(n861), 
        .Y(n44) );
  scg6d1_hd U1307 ( .A(r_mult_3_A[9]), .B(n858), .C(n859), .Y(n99) );
  scg14d1_hd U1308 ( .A(r_mult_3_A[10]), .B(n858), .C(n857), .Y(n98) );
  scg14d1_hd U1309 ( .A(r_mult_3_A[11]), .B(n858), .C(n857), .Y(n97) );
  scg6d1_hd U1310 ( .A(r_mult_3_A[13]), .B(n858), .C(n859), .Y(n95) );
  scg6d1_hd U1311 ( .A(r_mult_3_A[14]), .B(n858), .C(n859), .Y(n94) );
  scg14d1_hd U1312 ( .A(r_mult_3_A[15]), .B(n858), .C(n857), .Y(n93) );
  scg6d1_hd U1313 ( .A(r_mult_3_A[16]), .B(n858), .C(n859), .Y(n92) );
  scg14d1_hd U1314 ( .A(r_mult_3_A[18]), .B(n858), .C(n857), .Y(n90) );
  scg6d1_hd U1315 ( .A(r_mult_3_A[19]), .B(n858), .C(n859), .Y(n89) );
  scg6d1_hd U1316 ( .A(r_mult_3_A[20]), .B(n858), .C(n859), .Y(n88) );
  scg14d1_hd U1317 ( .A(r_mult_3_A[21]), .B(n858), .C(n857), .Y(n87) );
  scg14d1_hd U1318 ( .A(r_mult_3_A[22]), .B(n858), .C(n860), .Y(n86) );
  scg14d1_hd U1319 ( .A(r_mult_3_A[23]), .B(n858), .C(n857), .Y(n85) );
  scg14d1_hd U1320 ( .A(r_mult_3_A[24]), .B(n858), .C(n857), .Y(n84) );
  ad2d1_hd U1321 ( .A(r_mult_3_A[30]), .B(n858), .Y(n78) );
  scg14d1_hd U1322 ( .A(r_mult_3_A[31]), .B(n858), .C(n857), .Y(n77) );
  scg5d1_hd U1323 ( .A(n831), .B(r_mult_1_B[0]), .C(n862), .D(w_add_1_Z[0]), 
        .E(n834), .F(r_x_data[64]), .Y(n76) );
  scg5d1_hd U1324 ( .A(n831), .B(r_mult_1_B[1]), .C(n862), .D(w_add_1_Z[1]), 
        .E(n834), .F(r_x_data[65]), .Y(n75) );
  scg5d1_hd U1325 ( .A(n831), .B(r_mult_1_B[2]), .C(n862), .D(w_add_1_Z[2]), 
        .E(n834), .F(r_x_data[66]), .Y(n74) );
  scg5d1_hd U1326 ( .A(n861), .B(r_mult_1_B[3]), .C(n862), .D(w_add_1_Z[3]), 
        .E(n834), .F(r_x_data[67]), .Y(n73) );
  scg5d1_hd U1327 ( .A(n831), .B(r_mult_1_B[4]), .C(n862), .D(w_add_1_Z[4]), 
        .E(n834), .F(r_x_data[68]), .Y(n72) );
  scg5d1_hd U1328 ( .A(n831), .B(r_mult_1_B[5]), .C(n862), .D(w_add_1_Z[5]), 
        .E(n830), .F(r_x_data[69]), .Y(n71) );
  scg5d1_hd U1329 ( .A(n861), .B(r_mult_1_B[6]), .C(n862), .D(w_add_1_Z[6]), 
        .E(n830), .F(r_x_data[70]), .Y(n70) );
  scg5d1_hd U1330 ( .A(n831), .B(r_mult_1_B[7]), .C(n862), .D(w_add_1_Z[7]), 
        .E(n834), .F(r_x_data[71]), .Y(n69) );
  scg5d1_hd U1331 ( .A(n831), .B(r_mult_1_B[8]), .C(n862), .D(w_add_1_Z[8]), 
        .E(n830), .F(r_x_data[72]), .Y(n68) );
  scg5d1_hd U1332 ( .A(n831), .B(r_mult_1_B[9]), .C(n862), .D(w_add_1_Z[9]), 
        .E(n830), .F(r_x_data[73]), .Y(n67) );
  scg5d1_hd U1333 ( .A(n831), .B(r_mult_1_B[10]), .C(n862), .D(w_add_1_Z[10]), 
        .E(n834), .F(r_x_data[74]), .Y(n66) );
  scg5d1_hd U1334 ( .A(n831), .B(r_mult_1_B[11]), .C(n862), .D(w_add_1_Z[11]), 
        .E(n830), .F(r_x_data[75]), .Y(n65) );
  scg5d1_hd U1335 ( .A(n831), .B(r_mult_1_B[12]), .C(n862), .D(w_add_1_Z[12]), 
        .E(n832), .F(r_x_data[76]), .Y(n64) );
  scg5d1_hd U1336 ( .A(n831), .B(r_mult_1_B[13]), .C(n862), .D(w_add_1_Z[13]), 
        .E(n834), .F(r_x_data[77]), .Y(n63) );
  scg5d1_hd U1337 ( .A(n831), .B(r_mult_1_B[14]), .C(n862), .D(w_add_1_Z[14]), 
        .E(n830), .F(r_x_data[78]), .Y(n62) );
  scg5d1_hd U1338 ( .A(n831), .B(r_mult_1_B[15]), .C(n862), .D(w_add_1_Z[15]), 
        .E(n832), .F(r_x_data[79]), .Y(n61) );
  scg5d1_hd U1339 ( .A(n831), .B(r_mult_1_B[16]), .C(n862), .D(w_add_1_Z[16]), 
        .E(n830), .F(r_x_data[80]), .Y(n60) );
  scg5d1_hd U1340 ( .A(n831), .B(r_mult_1_B[17]), .C(n862), .D(w_add_1_Z[17]), 
        .E(n832), .F(r_x_data[81]), .Y(n59) );
  scg5d1_hd U1341 ( .A(n831), .B(r_mult_1_B[18]), .C(n862), .D(w_add_1_Z[18]), 
        .E(n834), .F(r_x_data[82]), .Y(n58) );
  scg5d1_hd U1342 ( .A(n831), .B(r_mult_1_B[19]), .C(n862), .D(w_add_1_Z[19]), 
        .E(n834), .F(r_x_data[83]), .Y(n57) );
  scg5d1_hd U1343 ( .A(n831), .B(r_mult_1_B[20]), .C(n862), .D(w_add_1_Z[20]), 
        .E(n830), .F(r_x_data[84]), .Y(n56) );
  scg5d1_hd U1344 ( .A(n831), .B(r_mult_1_B[21]), .C(n862), .D(w_add_1_Z[21]), 
        .E(n834), .F(r_x_data[85]), .Y(n55) );
  scg5d1_hd U1345 ( .A(n831), .B(r_mult_1_B[22]), .C(n862), .D(w_add_1_Z[22]), 
        .E(n832), .F(r_x_data[86]), .Y(n54) );
  scg4d1_hd U1346 ( .A(n831), .B(r_mult_1_B[23]), .C(n906), .D(n4), .E(n862), 
        .F(w_add_1_Z[23]), .G(n832), .H(r_x_data[87]), .Y(n53) );
  scg4d1_hd U1347 ( .A(n831), .B(r_mult_1_B[24]), .C(n906), .D(n4), .E(n862), 
        .F(w_add_1_Z[24]), .G(n832), .H(r_x_data[88]), .Y(n52) );
  scg4d1_hd U1348 ( .A(n831), .B(r_mult_1_B[25]), .C(n906), .D(n4), .E(n862), 
        .F(w_add_1_Z[25]), .G(n830), .H(r_x_data[89]), .Y(n51) );
  ao22d1_hd U1349 ( .A(w_mult_1_Z[0]), .B(n864), .C(r_mult_1_A[0]), .D(n831), 
        .Y(n863) );
  scg5d1_hd U1350 ( .A(n858), .B(r_mult_3_B[31]), .C(n834), .D(r_y_data[63]), 
        .E(n859), .F(r_y_data[95]), .Y(n501) );
  scg4d1_hd U1351 ( .A(n831), .B(r_mult_1_B[26]), .C(n906), .D(n4), .E(n862), 
        .F(w_add_1_Z[26]), .G(n832), .H(r_x_data[90]), .Y(n50) );
  scg4d1_hd U1352 ( .A(n831), .B(r_mult_2_B[31]), .C(n862), .D(w_add_2_Z[31]), 
        .E(r_y_data[31]), .F(n832), .G(r_y_data[127]), .H(n907), .Y(n499) );
  scg14d1_hd U1353 ( .A(n865), .B(r_mult_3_Z_ACK), .C(n866), .Y(n497) );
  scg6d1_hd U1354 ( .A(n865), .B(r_mult_1_Z_ACK), .C(n867), .Y(n493) );
  scg6d1_hd U1355 ( .A(n865), .B(r_mult_2_Z_ACK), .C(n867), .Y(n492) );
  scg14d1_hd U1356 ( .A(n963), .B(r_mult_1_AB_STB), .C(n869), .Y(n491) );
  scg14d1_hd U1357 ( .A(n963), .B(r_mult_2_AB_STB), .C(n869), .Y(n490) );
  scg18d1_hd U1358 ( .A(n1040), .B(r_counter_1_), .C(n1077), .D(N1401), .E(
        n870), .Y(n869) );
  scg4d1_hd U1359 ( .A(n831), .B(r_mult_1_B[27]), .C(n906), .D(n4), .E(n862), 
        .F(w_add_1_Z[27]), .G(n834), .H(r_x_data[91]), .Y(n49) );
  scg4d1_hd U1360 ( .A(n861), .B(r_mult_1_B[28]), .C(n906), .D(n4), .E(n862), 
        .F(w_add_1_Z[28]), .G(n834), .H(r_x_data[92]), .Y(n48) );
  scg4d1_hd U1361 ( .A(n831), .B(r_mult_1_B[29]), .C(n906), .D(n4), .E(n862), 
        .F(w_add_1_Z[29]), .G(n830), .H(r_x_data[93]), .Y(n47) );
  scg5d1_hd U1362 ( .A(n831), .B(r_mult_1_B[30]), .C(n862), .D(w_add_1_Z[30]), 
        .E(n834), .F(r_x_data[94]), .Y(n46) );
  scg5d1_hd U1363 ( .A(n831), .B(r_mult_1_B[31]), .C(n862), .D(w_add_1_Z[31]), 
        .E(n830), .F(r_x_data[95]), .Y(n45) );
  ao22d1_hd U1364 ( .A(w_mult_1_Z[2]), .B(n907), .C(r_mult_1_A[2]), .D(n831), 
        .Y(n871) );
  ao22d1_hd U1365 ( .A(w_mult_1_Z[3]), .B(n907), .C(r_mult_1_A[3]), .D(n861), 
        .Y(n874) );
  ao22d1_hd U1366 ( .A(w_mult_1_Z[4]), .B(n864), .C(r_mult_1_A[4]), .D(n831), 
        .Y(n875) );
  ao22d1_hd U1367 ( .A(w_mult_1_Z[5]), .B(n864), .C(r_mult_1_A[5]), .D(n861), 
        .Y(n876) );
  ao22d1_hd U1368 ( .A(w_mult_1_Z[7]), .B(n907), .C(r_mult_1_A[7]), .D(n831), 
        .Y(n877) );
  ao22d1_hd U1369 ( .A(w_mult_1_Z[10]), .B(n907), .C(r_mult_1_A[10]), .D(n831), 
        .Y(n878) );
  ao22d1_hd U1370 ( .A(w_mult_1_Z[11]), .B(n864), .C(r_mult_1_A[11]), .D(n831), 
        .Y(n879) );
  ao22d1_hd U1371 ( .A(w_mult_1_Z[13]), .B(n864), .C(r_mult_1_A[13]), .D(n831), 
        .Y(n880) );
  ao22d1_hd U1372 ( .A(w_mult_1_Z[14]), .B(n907), .C(r_mult_1_A[14]), .D(n861), 
        .Y(n881) );
  ao22d1_hd U1373 ( .A(w_mult_1_Z[15]), .B(n907), .C(r_mult_1_A[15]), .D(n831), 
        .Y(n882) );
  ao22d1_hd U1374 ( .A(w_mult_1_Z[17]), .B(n864), .C(r_mult_1_A[17]), .D(n861), 
        .Y(n883) );
  ao22d1_hd U1375 ( .A(w_mult_1_Z[18]), .B(n864), .C(r_mult_1_A[18]), .D(n861), 
        .Y(n884) );
  ao22d1_hd U1376 ( .A(w_mult_1_Z[19]), .B(n907), .C(r_mult_1_A[19]), .D(n861), 
        .Y(n885) );
  ao22d1_hd U1377 ( .A(w_mult_1_Z[21]), .B(n907), .C(r_mult_1_A[21]), .D(n831), 
        .Y(n886) );
  ao22d1_hd U1378 ( .A(w_mult_1_Z[22]), .B(n864), .C(r_mult_1_A[22]), .D(n861), 
        .Y(n887) );
  ao22d1_hd U1379 ( .A(w_mult_1_Z[23]), .B(n864), .C(r_mult_1_A[23]), .D(n861), 
        .Y(n888) );
  ao22d1_hd U1380 ( .A(w_mult_1_Z[24]), .B(n907), .C(r_mult_1_A[24]), .D(n861), 
        .Y(n889) );
  scg4d1_hd U1381 ( .A(n831), .B(r_mult_2_B[0]), .C(n862), .D(w_add_2_Z[0]), 
        .E(r_y_data[0]), .F(n830), .G(r_y_data[96]), .H(n907), .Y(n202) );
  scg4d1_hd U1382 ( .A(n831), .B(r_mult_2_B[1]), .C(n862), .D(w_add_2_Z[1]), 
        .E(r_y_data[1]), .F(n832), .G(r_y_data[97]), .H(n907), .Y(n201) );
  scg4d1_hd U1383 ( .A(n861), .B(r_mult_2_B[2]), .C(n862), .D(w_add_2_Z[2]), 
        .E(r_y_data[2]), .F(n832), .G(r_y_data[98]), .H(n907), .Y(n200) );
  ao22d1_hd U1384 ( .A(w_mult_1_Z[25]), .B(n907), .C(r_mult_1_A[25]), .D(n831), 
        .Y(n890) );
  scg4d1_hd U1385 ( .A(n831), .B(r_mult_2_B[3]), .C(n862), .D(w_add_2_Z[3]), 
        .E(r_y_data[3]), .F(n832), .G(r_y_data[99]), .H(n907), .Y(n199) );
  scg4d1_hd U1386 ( .A(n861), .B(r_mult_2_B[4]), .C(n862), .D(w_add_2_Z[4]), 
        .E(r_y_data[4]), .F(n832), .G(r_y_data[100]), .H(n907), .Y(n198) );
  scg4d1_hd U1387 ( .A(n861), .B(r_mult_2_B[5]), .C(n862), .D(w_add_2_Z[5]), 
        .E(r_y_data[5]), .F(n834), .G(r_y_data[101]), .H(n907), .Y(n197) );
  scg4d1_hd U1388 ( .A(n831), .B(r_mult_2_B[6]), .C(n862), .D(w_add_2_Z[6]), 
        .E(r_y_data[6]), .F(n834), .G(r_y_data[102]), .H(n907), .Y(n196) );
  scg4d1_hd U1389 ( .A(n831), .B(r_mult_2_B[7]), .C(n862), .D(w_add_2_Z[7]), 
        .E(r_y_data[7]), .F(n834), .G(r_y_data[103]), .H(n907), .Y(n195) );
  scg4d1_hd U1390 ( .A(n861), .B(r_mult_2_B[8]), .C(n862), .D(w_add_2_Z[8]), 
        .E(r_y_data[8]), .F(n834), .G(r_y_data[104]), .H(n907), .Y(n194) );
  scg4d1_hd U1391 ( .A(n831), .B(r_mult_2_B[9]), .C(n862), .D(w_add_2_Z[9]), 
        .E(r_y_data[9]), .F(n834), .G(r_y_data[105]), .H(n907), .Y(n193) );
  scg4d1_hd U1392 ( .A(n831), .B(r_mult_2_B[10]), .C(n862), .D(w_add_2_Z[10]), 
        .E(r_y_data[10]), .F(n830), .G(r_y_data[106]), .H(n907), .Y(n192) );
  scg4d1_hd U1393 ( .A(n861), .B(r_mult_2_B[11]), .C(n862), .D(w_add_2_Z[11]), 
        .E(r_y_data[11]), .F(n830), .G(r_y_data[107]), .H(n907), .Y(n191) );
  scg4d1_hd U1394 ( .A(n861), .B(r_mult_2_B[12]), .C(n862), .D(w_add_2_Z[12]), 
        .E(r_y_data[12]), .F(n832), .G(r_y_data[108]), .H(n907), .Y(n190) );
  ao22d1_hd U1395 ( .A(w_mult_1_Z[26]), .B(n864), .C(r_mult_1_A[26]), .D(n861), 
        .Y(n891) );
  scg4d1_hd U1396 ( .A(n861), .B(r_mult_2_B[13]), .C(n862), .D(w_add_2_Z[13]), 
        .E(r_y_data[13]), .F(n832), .G(r_y_data[109]), .H(n907), .Y(n189) );
  scg4d1_hd U1397 ( .A(n861), .B(r_mult_2_B[14]), .C(n862), .D(w_add_2_Z[14]), 
        .E(r_y_data[14]), .F(n834), .G(r_y_data[110]), .H(n907), .Y(n188) );
  scg4d1_hd U1398 ( .A(n861), .B(r_mult_2_B[15]), .C(n862), .D(w_add_2_Z[15]), 
        .E(r_y_data[15]), .F(n830), .G(r_y_data[111]), .H(n907), .Y(n187) );
  scg4d1_hd U1399 ( .A(n861), .B(r_mult_2_B[16]), .C(n862), .D(w_add_2_Z[16]), 
        .E(r_y_data[16]), .F(n832), .G(r_y_data[112]), .H(n907), .Y(n186) );
  scg4d1_hd U1400 ( .A(n861), .B(r_mult_2_B[17]), .C(n862), .D(w_add_2_Z[17]), 
        .E(r_y_data[17]), .F(n832), .G(r_y_data[113]), .H(n907), .Y(n185) );
  scg4d1_hd U1401 ( .A(n861), .B(r_mult_2_B[18]), .C(n862), .D(w_add_2_Z[18]), 
        .E(r_y_data[18]), .F(n834), .G(r_y_data[114]), .H(n907), .Y(n184) );
  scg4d1_hd U1402 ( .A(n861), .B(r_mult_2_B[19]), .C(n862), .D(w_add_2_Z[19]), 
        .E(r_y_data[19]), .F(n834), .G(r_y_data[115]), .H(n907), .Y(n183) );
  scg4d1_hd U1403 ( .A(n861), .B(r_mult_2_B[20]), .C(n862), .D(w_add_2_Z[20]), 
        .E(r_y_data[20]), .F(n830), .G(r_y_data[116]), .H(n907), .Y(n182) );
  scg4d1_hd U1404 ( .A(n861), .B(r_mult_2_B[21]), .C(n862), .D(w_add_2_Z[21]), 
        .E(r_y_data[21]), .F(n832), .G(r_y_data[117]), .H(n907), .Y(n181) );
  scg4d1_hd U1405 ( .A(n861), .B(r_mult_2_B[22]), .C(n862), .D(w_add_2_Z[22]), 
        .E(r_y_data[22]), .F(n832), .G(r_y_data[118]), .H(n907), .Y(n180) );
  ao22d1_hd U1406 ( .A(w_mult_1_Z[27]), .B(n864), .C(r_mult_1_A[27]), .D(n831), 
        .Y(n892) );
  scg4d1_hd U1407 ( .A(n861), .B(r_mult_2_B[23]), .C(n862), .D(w_add_2_Z[23]), 
        .E(r_y_data[23]), .F(n832), .G(r_y_data[119]), .H(n907), .Y(n179) );
  scg4d1_hd U1408 ( .A(n861), .B(r_mult_2_B[24]), .C(n862), .D(w_add_2_Z[24]), 
        .E(r_y_data[24]), .F(n834), .G(r_y_data[120]), .H(n907), .Y(n178) );
  scg4d1_hd U1409 ( .A(n861), .B(r_mult_2_B[25]), .C(n862), .D(w_add_2_Z[25]), 
        .E(r_y_data[25]), .F(n834), .G(r_y_data[121]), .H(n907), .Y(n177) );
  scg4d1_hd U1410 ( .A(n861), .B(r_mult_2_B[26]), .C(n862), .D(w_add_2_Z[26]), 
        .E(r_y_data[26]), .F(n830), .G(r_y_data[122]), .H(n864), .Y(n176) );
  scg4d1_hd U1411 ( .A(n831), .B(r_mult_2_B[27]), .C(n862), .D(w_add_2_Z[27]), 
        .E(r_y_data[27]), .F(n830), .G(r_y_data[123]), .H(n864), .Y(n175) );
  scg4d1_hd U1412 ( .A(n861), .B(r_mult_2_B[28]), .C(n862), .D(w_add_2_Z[28]), 
        .E(r_y_data[28]), .F(n832), .G(r_y_data[124]), .H(n907), .Y(n174) );
  scg4d1_hd U1413 ( .A(n831), .B(r_mult_2_B[29]), .C(n862), .D(w_add_2_Z[29]), 
        .E(r_y_data[29]), .F(n832), .G(r_y_data[125]), .H(n907), .Y(n173) );
  scg4d1_hd U1414 ( .A(n861), .B(r_mult_2_B[30]), .C(n862), .D(w_add_2_Z[30]), 
        .E(r_y_data[30]), .F(n832), .G(r_y_data[126]), .H(n864), .Y(n172) );
  scg6d1_hd U1415 ( .A(r_mult_2_A[0]), .B(n831), .C(n864), .Y(n171) );
  scg14d1_hd U1416 ( .A(r_mult_2_A[1]), .B(n831), .C(n857), .Y(n170) );
  ao22d1_hd U1417 ( .A(w_mult_1_Z[28]), .B(n907), .C(r_mult_1_A[28]), .D(n861), 
        .Y(n893) );
  ad2d1_hd U1418 ( .A(r_mult_2_A[2]), .B(n831), .Y(n169) );
  nd2bd1_hd U1419 ( .AN(r_mult_2_A[3]), .B(n894), .Y(n168) );
  scg14d1_hd U1420 ( .A(r_mult_2_A[4]), .B(n831), .C(n857), .Y(n167) );
  scg6d1_hd U1421 ( .A(r_mult_2_A[5]), .B(n831), .C(n862), .Y(n166) );
  nd2bd1_hd U1422 ( .AN(r_mult_2_A[6]), .B(n894), .Y(n165) );
  scg14d1_hd U1423 ( .A(r_mult_2_A[7]), .B(n831), .C(n866), .Y(n164) );
  nd2bd1_hd U1424 ( .AN(r_mult_2_A[8]), .B(n894), .Y(n163) );
  scg14d1_hd U1425 ( .A(r_mult_2_A[9]), .B(n831), .C(n873), .Y(n162) );
  nd2bd1_hd U1426 ( .AN(r_mult_2_A[10]), .B(n894), .Y(n161) );
  ad2d1_hd U1427 ( .A(r_mult_2_A[11]), .B(n831), .Y(n160) );
  ao22d1_hd U1428 ( .A(w_mult_1_Z[29]), .B(n907), .C(r_mult_1_A[29]), .D(n831), 
        .Y(n895) );
  scg17d1_hd U1429 ( .A(r_mult_2_A[12]), .B(n861), .C(n864), .D(n857), .Y(n159) );
  scg14d1_hd U1430 ( .A(r_mult_2_A[13]), .B(n831), .C(n857), .Y(n158) );
  scg14d1_hd U1431 ( .A(r_mult_2_A[14]), .B(n831), .C(n866), .Y(n157) );
  scg6d1_hd U1432 ( .A(r_mult_2_A[15]), .B(n861), .C(n907), .Y(n156) );
  ad2d1_hd U1433 ( .A(r_mult_2_A[16]), .B(n831), .Y(n155) );
  scg6d1_hd U1434 ( .A(r_mult_2_A[17]), .B(n831), .C(n907), .Y(n154) );
  scg17d1_hd U1435 ( .A(r_mult_2_A[18]), .B(n831), .C(n907), .D(n857), .Y(n153) );
  scg14d1_hd U1436 ( .A(r_mult_2_A[19]), .B(n831), .C(n866), .Y(n152) );
  scg14d1_hd U1437 ( .A(r_mult_2_A[20]), .B(n831), .C(n857), .Y(n151) );
  scg14d1_hd U1438 ( .A(r_mult_2_A[21]), .B(n831), .C(n873), .Y(n150) );
  nd2bd1_hd U1439 ( .AN(r_mult_2_A[22]), .B(n894), .Y(n149) );
  ad2d1_hd U1440 ( .A(r_mult_2_A[23]), .B(n831), .Y(n148) );
  scg6d1_hd U1441 ( .A(r_mult_2_A[24]), .B(n861), .C(n864), .Y(n147) );
  nd2bd1_hd U1442 ( .AN(r_mult_2_A[25]), .B(n894), .Y(n146) );
  nd2bd1_hd U1443 ( .AN(r_mult_2_A[26]), .B(n894), .Y(n145) );
  nd2bd1_hd U1444 ( .AN(r_mult_2_A[27]), .B(n894), .Y(n144) );
  nd2bd1_hd U1445 ( .AN(r_mult_2_A[28]), .B(n894), .Y(n143) );
  nd2bd1_hd U1446 ( .AN(r_mult_2_A[29]), .B(n894), .Y(n142) );
  ad2d1_hd U1447 ( .A(r_mult_2_A[30]), .B(n831), .Y(n141) );
  scg14d1_hd U1448 ( .A(r_mult_2_A[31]), .B(n831), .C(n866), .Y(n140) );
  scg5d1_hd U1449 ( .A(n858), .B(r_mult_3_B[0]), .C(n830), .D(r_y_data[32]), 
        .E(n859), .F(r_y_data[64]), .Y(n139) );
  scg5d1_hd U1450 ( .A(n858), .B(r_mult_3_B[1]), .C(n832), .D(r_y_data[33]), 
        .E(n859), .F(r_y_data[65]), .Y(n138) );
  scg5d1_hd U1451 ( .A(n858), .B(r_mult_3_B[2]), .C(n830), .D(r_y_data[34]), 
        .E(n859), .F(r_y_data[66]), .Y(n137) );
  scg5d1_hd U1452 ( .A(n858), .B(r_mult_3_B[3]), .C(n834), .D(r_y_data[35]), 
        .E(n859), .F(r_y_data[67]), .Y(n136) );
  scg5d1_hd U1453 ( .A(n858), .B(r_mult_3_B[4]), .C(n830), .D(r_y_data[36]), 
        .E(n859), .F(r_y_data[68]), .Y(n135) );
  scg5d1_hd U1454 ( .A(n858), .B(r_mult_3_B[5]), .C(n834), .D(r_y_data[37]), 
        .E(n859), .F(r_y_data[69]), .Y(n134) );
  scg5d1_hd U1455 ( .A(n858), .B(r_mult_3_B[6]), .C(n830), .D(r_y_data[38]), 
        .E(n859), .F(r_y_data[70]), .Y(n133) );
  scg5d1_hd U1456 ( .A(n858), .B(r_mult_3_B[7]), .C(n832), .D(r_y_data[39]), 
        .E(n859), .F(r_y_data[71]), .Y(n132) );
  scg5d1_hd U1457 ( .A(n858), .B(r_mult_3_B[8]), .C(n832), .D(r_y_data[40]), 
        .E(n859), .F(r_y_data[72]), .Y(n131) );
  scg5d1_hd U1458 ( .A(n858), .B(r_mult_3_B[9]), .C(n832), .D(r_y_data[41]), 
        .E(n859), .F(r_y_data[73]), .Y(n130) );
  scg5d1_hd U1459 ( .A(n858), .B(r_mult_3_B[10]), .C(n830), .D(r_y_data[42]), 
        .E(n859), .F(r_y_data[74]), .Y(n129) );
  scg5d1_hd U1460 ( .A(n858), .B(r_mult_3_B[11]), .C(n834), .D(r_y_data[43]), 
        .E(n859), .F(r_y_data[75]), .Y(n128) );
  scg5d1_hd U1461 ( .A(n858), .B(r_mult_3_B[12]), .C(n830), .D(r_y_data[44]), 
        .E(n859), .F(r_y_data[76]), .Y(n127) );
  scg5d1_hd U1462 ( .A(n858), .B(r_mult_3_B[13]), .C(n834), .D(r_y_data[45]), 
        .E(n859), .F(r_y_data[77]), .Y(n126) );
  scg5d1_hd U1463 ( .A(n858), .B(r_mult_3_B[14]), .C(n834), .D(r_y_data[46]), 
        .E(n859), .F(r_y_data[78]), .Y(n125) );
  scg5d1_hd U1464 ( .A(n858), .B(r_mult_3_B[15]), .C(n834), .D(r_y_data[47]), 
        .E(n859), .F(r_y_data[79]), .Y(n124) );
  scg5d1_hd U1465 ( .A(n858), .B(r_mult_3_B[16]), .C(n830), .D(r_y_data[48]), 
        .E(n859), .F(r_y_data[80]), .Y(n123) );
  scg5d1_hd U1466 ( .A(n858), .B(r_mult_3_B[17]), .C(n830), .D(r_y_data[49]), 
        .E(n859), .F(r_y_data[81]), .Y(n122) );
  scg5d1_hd U1467 ( .A(n858), .B(r_mult_3_B[18]), .C(n834), .D(r_y_data[50]), 
        .E(n859), .F(r_y_data[82]), .Y(n121) );
  scg5d1_hd U1468 ( .A(n858), .B(r_mult_3_B[19]), .C(n830), .D(r_y_data[51]), 
        .E(n859), .F(r_y_data[83]), .Y(n120) );
  scg5d1_hd U1469 ( .A(n858), .B(r_mult_3_B[20]), .C(n834), .D(r_y_data[52]), 
        .E(n859), .F(r_y_data[84]), .Y(n119) );
  scg5d1_hd U1470 ( .A(n858), .B(r_mult_3_B[21]), .C(n834), .D(r_y_data[53]), 
        .E(n859), .F(r_y_data[85]), .Y(n118) );
  scg5d1_hd U1471 ( .A(n858), .B(r_mult_3_B[22]), .C(n834), .D(r_y_data[54]), 
        .E(n859), .F(r_y_data[86]), .Y(n117) );
  scg5d1_hd U1472 ( .A(n858), .B(r_mult_3_B[23]), .C(n834), .D(r_y_data[55]), 
        .E(n859), .F(r_y_data[87]), .Y(n116) );
  scg5d1_hd U1473 ( .A(n858), .B(r_mult_3_B[24]), .C(n830), .D(r_y_data[56]), 
        .E(n859), .F(r_y_data[88]), .Y(n115) );
  scg5d1_hd U1474 ( .A(n858), .B(r_mult_3_B[25]), .C(n830), .D(r_y_data[57]), 
        .E(n859), .F(r_y_data[89]), .Y(n114) );
  scg5d1_hd U1475 ( .A(n858), .B(r_mult_3_B[26]), .C(n834), .D(r_y_data[58]), 
        .E(n859), .F(r_y_data[90]), .Y(n113) );
  scg5d1_hd U1476 ( .A(n858), .B(r_mult_3_B[27]), .C(n834), .D(r_y_data[59]), 
        .E(n859), .F(r_y_data[91]), .Y(n112) );
  scg5d1_hd U1477 ( .A(n858), .B(r_mult_3_B[28]), .C(n834), .D(r_y_data[60]), 
        .E(n859), .F(r_y_data[92]), .Y(n111) );
  scg5d1_hd U1478 ( .A(n858), .B(r_mult_3_B[29]), .C(n834), .D(r_y_data[61]), 
        .E(n859), .F(r_y_data[93]), .Y(n110) );
  scg5d1_hd U1479 ( .A(n858), .B(r_mult_3_B[30]), .C(n830), .D(r_y_data[62]), 
        .E(n859), .F(r_y_data[94]), .Y(n109) );
  scg6d1_hd U1480 ( .A(r_mult_3_A[0]), .B(n858), .C(n859), .Y(n108) );
  scg6d1_hd U1481 ( .A(r_mult_3_A[1]), .B(n858), .C(n859), .Y(n107) );
  scg14d1_hd U1482 ( .A(r_mult_3_A[2]), .B(n858), .C(n857), .Y(n106) );
  scg6d1_hd U1483 ( .A(r_mult_3_A[6]), .B(n858), .C(n859), .Y(n102) );
  scg6d1_hd U1484 ( .A(r_mult_3_A[8]), .B(n858), .C(n830), .Y(n100) );
  ao21d1_hd U1485 ( .A(n506), .B(n7), .C(n870), .Y(n897) );
  oa21d1_hd U1486 ( .A(n495), .B(n962), .C(n5), .Y(n901) );
  nr2d1_hd U1487 ( .A(n956), .B(n957), .Y(N1343) );
  ao211d1_hd U1488 ( .A(i_Y_ACK), .B(o_Y_DATA_VALID), .C(n542), .D(n909), .Y(
        n1038) );
  ivd1_hd U1489 ( .A(n917), .Y(n910) );
  ao22d1_hd U1490 ( .A(n916), .B(n506), .C(n962), .D(n910), .Y(n913) );
  ao21d1_hd U1491 ( .A(n1035), .B(n1040), .C(n1077), .Y(n911) );
  oa211d1_hd U1492 ( .A(N739), .B(n1040), .C(r_counter_1_), .D(n911), .Y(n912)
         );
  ao21d1_hd U1493 ( .A(n913), .B(n912), .C(n1079), .Y(n958) );
  ao211d1_hd U1494 ( .A(n959), .B(n843), .C(n1038), .D(n958), .Y(n914) );
  oa21d1_hd U1495 ( .A(n659), .B(n957), .C(n914), .Y(N1383) );
  nr2bd1_hd U1496 ( .AN(n959), .B(N23), .Y(N1402) );
  nr2d1_hd U1497 ( .A(N23), .B(n963), .Y(N1403) );
  nd4d1_hd U1498 ( .A(n829), .B(w_add_2_Z_STB), .C(w_add_1_Z_STB), .D(n1042), 
        .Y(n915) );
  scg4d1_hd U1499 ( .A(n840), .B(r_add_1_B[19]), .C(n841), .D(w_add_1_Z[19]), 
        .E(n834), .F(r_x_data[147]), .G(w_add_2_Z[19]), .H(n839), .Y(n672) );
  scg4d1_hd U1500 ( .A(n841), .B(w_add_1_Z[20]), .C(n840), .D(r_add_1_B[20]), 
        .E(n839), .F(w_add_2_Z[20]), .G(r_x_data[148]), .H(n834), .Y(n671) );
  scg4d1_hd U1501 ( .A(n841), .B(w_add_1_Z[21]), .C(n840), .D(r_add_1_B[21]), 
        .E(n839), .F(w_add_2_Z[21]), .G(r_x_data[149]), .H(n834), .Y(n670) );
  scg4d1_hd U1502 ( .A(n841), .B(w_add_1_Z[22]), .C(n840), .D(r_add_1_B[22]), 
        .E(n839), .F(w_add_2_Z[22]), .G(r_x_data[150]), .H(n834), .Y(n669) );
  scg4d1_hd U1503 ( .A(n841), .B(w_add_1_Z[23]), .C(n840), .D(r_add_1_B[23]), 
        .E(n839), .F(w_add_2_Z[23]), .G(r_x_data[151]), .H(n830), .Y(n668) );
  scg4d1_hd U1504 ( .A(n841), .B(w_add_1_Z[24]), .C(n840), .D(r_add_1_B[24]), 
        .E(n839), .F(w_add_2_Z[24]), .G(r_x_data[152]), .H(n834), .Y(n667) );
  scg4d1_hd U1505 ( .A(n841), .B(w_add_1_Z[25]), .C(n840), .D(r_add_1_B[25]), 
        .E(n839), .F(w_add_2_Z[25]), .G(r_x_data[153]), .H(n832), .Y(n666) );
  scg4d1_hd U1506 ( .A(n841), .B(w_add_1_Z[26]), .C(n840), .D(r_add_1_B[26]), 
        .E(n839), .F(w_add_2_Z[26]), .G(r_x_data[154]), .H(n834), .Y(n665) );
  scg4d1_hd U1507 ( .A(n841), .B(w_add_1_Z[27]), .C(n840), .D(r_add_1_B[27]), 
        .E(n839), .F(w_add_2_Z[27]), .G(r_x_data[155]), .H(n834), .Y(n664) );
  scg4d1_hd U1508 ( .A(n841), .B(w_add_1_Z[28]), .C(n840), .D(r_add_1_B[28]), 
        .E(n839), .F(w_add_2_Z[28]), .G(r_x_data[156]), .H(n830), .Y(n663) );
  scg4d1_hd U1509 ( .A(n1034), .B(w_add_1_Z[29]), .C(n840), .D(r_add_1_B[29]), 
        .E(n839), .F(w_add_2_Z[29]), .G(r_x_data[157]), .H(n832), .Y(n662) );
  scg4d1_hd U1510 ( .A(n1034), .B(w_add_1_Z[30]), .C(n840), .D(r_add_1_B[30]), 
        .E(n839), .F(w_add_2_Z[30]), .G(r_x_data[158]), .H(n832), .Y(n661) );
  scg4d1_hd U1511 ( .A(n1034), .B(w_add_1_Z[31]), .C(n840), .D(r_add_1_B[31]), 
        .E(n839), .F(w_add_2_Z[31]), .G(r_x_data[159]), .H(n832), .Y(n660) );
  ivd1_hd U1512 ( .A(o_Y_DATA[31]), .Y(n919) );
  oa22d1_hd U1513 ( .A(n922), .B(n955), .C(n835), .D(n919), .Y(n827) );
  ao22d1_hd U1514 ( .A(r_x_data[31]), .B(n830), .C(r_add_1_A[31]), .D(n840), 
        .Y(n921) );
  oa211d1_hd U1515 ( .A(n836), .B(n922), .C(n651), .D(n921), .Y(n826) );
  ivd1_hd U1516 ( .A(o_Y_DATA[30]), .Y(n923) );
  oa22d1_hd U1517 ( .A(n1026), .B(n955), .C(n835), .D(n923), .Y(n825) );
  ivd1_hd U1518 ( .A(o_Y_DATA[29]), .Y(n924) );
  oa22d1_hd U1519 ( .A(n1024), .B(n955), .C(n835), .D(n924), .Y(n824) );
  ivd1_hd U1520 ( .A(o_Y_DATA[28]), .Y(n925) );
  oa22d1_hd U1521 ( .A(n1022), .B(n955), .C(n835), .D(n925), .Y(n823) );
  ivd1_hd U1522 ( .A(o_Y_DATA[27]), .Y(n926) );
  oa22d1_hd U1523 ( .A(n1020), .B(n955), .C(n835), .D(n926), .Y(n822) );
  ivd1_hd U1524 ( .A(o_Y_DATA[26]), .Y(n927) );
  oa22d1_hd U1525 ( .A(n1018), .B(n955), .C(n835), .D(n927), .Y(n821) );
  ivd1_hd U1526 ( .A(o_Y_DATA[25]), .Y(n928) );
  oa22d1_hd U1527 ( .A(n1016), .B(n955), .C(n835), .D(n928), .Y(n820) );
  ivd1_hd U1528 ( .A(o_Y_DATA[24]), .Y(n929) );
  oa22d1_hd U1529 ( .A(n1014), .B(n955), .C(n835), .D(n929), .Y(n819) );
  ivd1_hd U1530 ( .A(o_Y_DATA[23]), .Y(n930) );
  oa22d1_hd U1531 ( .A(n1012), .B(n955), .C(n835), .D(n930), .Y(n818) );
  ivd1_hd U1532 ( .A(o_Y_DATA[22]), .Y(n931) );
  oa22d1_hd U1533 ( .A(n1010), .B(n955), .C(n835), .D(n931), .Y(n817) );
  ivd1_hd U1534 ( .A(o_Y_DATA[21]), .Y(n932) );
  oa22d1_hd U1535 ( .A(n1008), .B(n955), .C(n835), .D(n932), .Y(n816) );
  ivd1_hd U1536 ( .A(o_Y_DATA[20]), .Y(n933) );
  oa22d1_hd U1537 ( .A(n1006), .B(n955), .C(n835), .D(n933), .Y(n815) );
  ivd1_hd U1538 ( .A(o_Y_DATA[19]), .Y(n934) );
  oa22d1_hd U1539 ( .A(n1004), .B(n955), .C(n835), .D(n934), .Y(n814) );
  ivd1_hd U1540 ( .A(o_Y_DATA[18]), .Y(n935) );
  oa22d1_hd U1541 ( .A(n1002), .B(n955), .C(n835), .D(n935), .Y(n813) );
  ivd1_hd U1542 ( .A(o_Y_DATA[17]), .Y(n936) );
  oa22d1_hd U1543 ( .A(n1000), .B(n955), .C(n835), .D(n936), .Y(n812) );
  ivd1_hd U1544 ( .A(o_Y_DATA[16]), .Y(n937) );
  oa22d1_hd U1545 ( .A(n998), .B(n955), .C(n835), .D(n937), .Y(n811) );
  ivd1_hd U1546 ( .A(o_Y_DATA[15]), .Y(n938) );
  oa22d1_hd U1547 ( .A(n996), .B(n955), .C(n835), .D(n938), .Y(n810) );
  ivd1_hd U1548 ( .A(o_Y_DATA[14]), .Y(n939) );
  oa22d1_hd U1549 ( .A(n994), .B(n955), .C(n835), .D(n939), .Y(n809) );
  ivd1_hd U1550 ( .A(o_Y_DATA[13]), .Y(n940) );
  oa22d1_hd U1551 ( .A(n992), .B(n955), .C(n954), .D(n940), .Y(n808) );
  ivd1_hd U1552 ( .A(o_Y_DATA[12]), .Y(n941) );
  oa22d1_hd U1553 ( .A(n990), .B(n955), .C(n954), .D(n941), .Y(n807) );
  ivd1_hd U1554 ( .A(o_Y_DATA[11]), .Y(n942) );
  oa22d1_hd U1555 ( .A(n988), .B(n955), .C(n954), .D(n942), .Y(n806) );
  ivd1_hd U1556 ( .A(o_Y_DATA[10]), .Y(n943) );
  oa22d1_hd U1557 ( .A(n986), .B(n955), .C(n835), .D(n943), .Y(n805) );
  ivd1_hd U1558 ( .A(o_Y_DATA[9]), .Y(n944) );
  oa22d1_hd U1559 ( .A(n984), .B(n955), .C(n835), .D(n944), .Y(n804) );
  ivd1_hd U1560 ( .A(o_Y_DATA[8]), .Y(n945) );
  oa22d1_hd U1561 ( .A(n982), .B(n955), .C(n835), .D(n945), .Y(n803) );
  ivd1_hd U1562 ( .A(o_Y_DATA[7]), .Y(n946) );
  oa22d1_hd U1563 ( .A(n980), .B(n955), .C(n835), .D(n946), .Y(n802) );
  ivd1_hd U1564 ( .A(o_Y_DATA[6]), .Y(n947) );
  oa22d1_hd U1565 ( .A(n978), .B(n955), .C(n835), .D(n947), .Y(n801) );
  ivd1_hd U1566 ( .A(o_Y_DATA[5]), .Y(n948) );
  oa22d1_hd U1567 ( .A(n976), .B(n955), .C(n835), .D(n948), .Y(n800) );
  ivd1_hd U1568 ( .A(o_Y_DATA[4]), .Y(n949) );
  oa22d1_hd U1569 ( .A(n974), .B(n955), .C(n835), .D(n949), .Y(n799) );
  ivd1_hd U1570 ( .A(o_Y_DATA[3]), .Y(n950) );
  oa22d1_hd U1571 ( .A(n972), .B(n955), .C(n835), .D(n950), .Y(n798) );
  ivd1_hd U1572 ( .A(o_Y_DATA[2]), .Y(n951) );
  oa22d1_hd U1573 ( .A(n970), .B(n955), .C(n835), .D(n951), .Y(n797) );
  ivd1_hd U1574 ( .A(o_Y_DATA[1]), .Y(n952) );
  oa22d1_hd U1575 ( .A(n968), .B(n955), .C(n835), .D(n952), .Y(n796) );
  ivd1_hd U1576 ( .A(o_Y_DATA[0]), .Y(n953) );
  oa22d1_hd U1577 ( .A(n966), .B(n955), .C(n835), .D(n953), .Y(n795) );
  scg21d1_hd U1578 ( .A(n495), .B(r_counter_1_), .C(n1041), .D(n1079), .Y(
        n1043) );
  oa22ad1_hd U1579 ( .A(n962), .B(n961), .C(r_counter_1_), .D(n1041), .Y(n791)
         );
  scg14d1_hd U1580 ( .A(n963), .B(r_add_1_AB_STB), .C(n964), .Y(n789) );
  oa22ad1_hd U1581 ( .A(n1077), .B(n964), .C(n963), .D(r_add_2_AB_STB), .Y(
        n788) );
  ao22d1_hd U1582 ( .A(r_x_data[0]), .B(n830), .C(r_add_1_A[0]), .D(n840), .Y(
        n965) );
  oa211d1_hd U1583 ( .A(n836), .B(n966), .C(n634), .D(n965), .Y(n787) );
  ao22d1_hd U1584 ( .A(r_x_data[1]), .B(n830), .C(r_add_1_A[1]), .D(n840), .Y(
        n967) );
  oa211d1_hd U1585 ( .A(n836), .B(n968), .C(n632), .D(n967), .Y(n786) );
  ao22d1_hd U1586 ( .A(r_x_data[2]), .B(n834), .C(r_add_1_A[2]), .D(n840), .Y(
        n969) );
  oa211d1_hd U1587 ( .A(n836), .B(n970), .C(n630), .D(n969), .Y(n785) );
  ao22d1_hd U1588 ( .A(r_x_data[3]), .B(n834), .C(r_add_1_A[3]), .D(n840), .Y(
        n971) );
  oa211d1_hd U1589 ( .A(n836), .B(n972), .C(n628), .D(n971), .Y(n784) );
  ao22d1_hd U1590 ( .A(r_x_data[4]), .B(n834), .C(r_add_1_A[4]), .D(n840), .Y(
        n973) );
  oa211d1_hd U1591 ( .A(n836), .B(n974), .C(n626), .D(n973), .Y(n783) );
  ao22d1_hd U1592 ( .A(r_x_data[5]), .B(n834), .C(r_add_1_A[5]), .D(n840), .Y(
        n975) );
  oa211d1_hd U1593 ( .A(n836), .B(n976), .C(n624), .D(n975), .Y(n782) );
  ao22d1_hd U1594 ( .A(r_x_data[6]), .B(n834), .C(r_add_1_A[6]), .D(n840), .Y(
        n977) );
  oa211d1_hd U1595 ( .A(n836), .B(n978), .C(n622), .D(n977), .Y(n781) );
  ao22d1_hd U1596 ( .A(r_x_data[7]), .B(n834), .C(r_add_1_A[7]), .D(n840), .Y(
        n979) );
  oa211d1_hd U1597 ( .A(n836), .B(n980), .C(n620), .D(n979), .Y(n780) );
  ao22d1_hd U1598 ( .A(r_x_data[8]), .B(n834), .C(r_add_1_A[8]), .D(n840), .Y(
        n981) );
  oa211d1_hd U1599 ( .A(n836), .B(n982), .C(n618), .D(n981), .Y(n779) );
  ao22d1_hd U1600 ( .A(r_x_data[9]), .B(n832), .C(r_add_1_A[9]), .D(n840), .Y(
        n983) );
  oa211d1_hd U1601 ( .A(n836), .B(n984), .C(n616), .D(n983), .Y(n778) );
  ao22d1_hd U1602 ( .A(r_x_data[10]), .B(n832), .C(r_add_1_A[10]), .D(n840), 
        .Y(n985) );
  oa211d1_hd U1603 ( .A(n837), .B(n986), .C(n614), .D(n985), .Y(n777) );
  ao22d1_hd U1604 ( .A(r_x_data[11]), .B(n832), .C(r_add_1_A[11]), .D(n840), 
        .Y(n987) );
  oa211d1_hd U1605 ( .A(n837), .B(n988), .C(n612), .D(n987), .Y(n776) );
  ao22d1_hd U1606 ( .A(r_x_data[12]), .B(n832), .C(r_add_1_A[12]), .D(n840), 
        .Y(n989) );
  oa211d1_hd U1607 ( .A(n837), .B(n990), .C(n610), .D(n989), .Y(n775) );
  ao22d1_hd U1608 ( .A(r_x_data[13]), .B(n832), .C(r_add_1_A[13]), .D(n840), 
        .Y(n991) );
  oa211d1_hd U1609 ( .A(n837), .B(n992), .C(n608), .D(n991), .Y(n774) );
  ao22d1_hd U1610 ( .A(r_x_data[14]), .B(n832), .C(r_add_1_A[14]), .D(n840), 
        .Y(n993) );
  oa211d1_hd U1611 ( .A(n837), .B(n994), .C(n606), .D(n993), .Y(n773) );
  ao22d1_hd U1612 ( .A(r_x_data[15]), .B(n830), .C(r_add_1_A[15]), .D(n840), 
        .Y(n995) );
  oa211d1_hd U1613 ( .A(n837), .B(n996), .C(n604), .D(n995), .Y(n772) );
  ao22d1_hd U1614 ( .A(r_x_data[16]), .B(n830), .C(r_add_1_A[16]), .D(n840), 
        .Y(n997) );
  oa211d1_hd U1615 ( .A(n837), .B(n998), .C(n602), .D(n997), .Y(n771) );
  ao22d1_hd U1616 ( .A(r_x_data[17]), .B(n830), .C(r_add_1_A[17]), .D(n840), 
        .Y(n999) );
  oa211d1_hd U1617 ( .A(n837), .B(n1000), .C(n600), .D(n999), .Y(n770) );
  ao22d1_hd U1618 ( .A(r_x_data[18]), .B(n834), .C(r_add_1_A[18]), .D(n840), 
        .Y(n1001) );
  oa211d1_hd U1619 ( .A(n837), .B(n1002), .C(n598), .D(n1001), .Y(n769) );
  ao22d1_hd U1620 ( .A(r_x_data[19]), .B(n834), .C(r_add_1_A[19]), .D(n840), 
        .Y(n1003) );
  oa211d1_hd U1621 ( .A(n837), .B(n1004), .C(n596), .D(n1003), .Y(n768) );
  ao22d1_hd U1622 ( .A(r_x_data[20]), .B(n834), .C(r_add_1_A[20]), .D(n840), 
        .Y(n1005) );
  oa211d1_hd U1623 ( .A(n837), .B(n1006), .C(n594), .D(n1005), .Y(n767) );
  ao22d1_hd U1624 ( .A(r_x_data[21]), .B(n834), .C(r_add_1_A[21]), .D(n840), 
        .Y(n1007) );
  oa211d1_hd U1625 ( .A(n838), .B(n1008), .C(n592), .D(n1007), .Y(n766) );
  ao22d1_hd U1626 ( .A(r_x_data[22]), .B(n834), .C(r_add_1_A[22]), .D(n840), 
        .Y(n1009) );
  oa211d1_hd U1627 ( .A(n838), .B(n1010), .C(n590), .D(n1009), .Y(n765) );
  ao22d1_hd U1628 ( .A(r_x_data[23]), .B(n834), .C(r_add_1_A[23]), .D(n840), 
        .Y(n1011) );
  oa211d1_hd U1629 ( .A(n838), .B(n1012), .C(n588), .D(n1011), .Y(n764) );
  ao22d1_hd U1630 ( .A(r_x_data[24]), .B(n834), .C(r_add_1_A[24]), .D(n840), 
        .Y(n1013) );
  oa211d1_hd U1631 ( .A(n838), .B(n1014), .C(n586), .D(n1013), .Y(n763) );
  ao22d1_hd U1632 ( .A(r_x_data[25]), .B(n832), .C(r_add_1_A[25]), .D(n840), 
        .Y(n1015) );
  oa211d1_hd U1633 ( .A(n838), .B(n1016), .C(n584), .D(n1015), .Y(n762) );
  ao22d1_hd U1634 ( .A(r_x_data[26]), .B(n832), .C(r_add_1_A[26]), .D(n840), 
        .Y(n1017) );
  oa211d1_hd U1635 ( .A(n838), .B(n1018), .C(n582), .D(n1017), .Y(n761) );
  ao22d1_hd U1636 ( .A(r_x_data[27]), .B(n832), .C(r_add_1_A[27]), .D(n840), 
        .Y(n1019) );
  oa211d1_hd U1637 ( .A(n838), .B(n1020), .C(n580), .D(n1019), .Y(n760) );
  ao22d1_hd U1638 ( .A(r_x_data[28]), .B(n832), .C(r_add_1_A[28]), .D(n840), 
        .Y(n1021) );
  oa211d1_hd U1639 ( .A(n838), .B(n1022), .C(n578), .D(n1021), .Y(n759) );
  ao22d1_hd U1640 ( .A(r_x_data[29]), .B(n832), .C(r_add_1_A[29]), .D(n840), 
        .Y(n1023) );
  oa211d1_hd U1641 ( .A(n838), .B(n1024), .C(n576), .D(n1023), .Y(n758) );
  ao22d1_hd U1642 ( .A(r_x_data[30]), .B(n832), .C(r_add_1_A[30]), .D(n840), 
        .Y(n1025) );
  oa211d1_hd U1643 ( .A(n838), .B(n1026), .C(n572), .D(n1025), .Y(n757) );
  scg16d1_hd U1644 ( .A(r_add_2_Z_ACK), .B(n1029), .C(n1028), .Y(n756) );
  oa21d1_hd U1645 ( .A(n1030), .B(n829), .C(o_Y_DATA_VALID), .Y(n1031) );
  nd2bd1_hd U1646 ( .AN(n1038), .B(n1031), .Y(n724) );
  scg4d1_hd U1647 ( .A(n1034), .B(w_add_1_Z[0]), .C(n840), .D(r_add_1_B[0]), 
        .E(n839), .F(w_add_2_Z[0]), .G(r_x_data[128]), .H(n830), .Y(n691) );
  scg4d1_hd U1648 ( .A(n1034), .B(w_add_1_Z[1]), .C(n840), .D(r_add_1_B[1]), 
        .E(n839), .F(w_add_2_Z[1]), .G(r_x_data[129]), .H(n830), .Y(n690) );
  scg4d1_hd U1649 ( .A(n841), .B(w_add_1_Z[2]), .C(n840), .D(r_add_1_B[2]), 
        .E(n839), .F(w_add_2_Z[2]), .G(r_x_data[130]), .H(n834), .Y(n689) );
  scg4d1_hd U1650 ( .A(n841), .B(w_add_1_Z[3]), .C(n840), .D(r_add_1_B[3]), 
        .E(n839), .F(w_add_2_Z[3]), .G(r_x_data[131]), .H(n832), .Y(n688) );
  scg4d1_hd U1651 ( .A(n841), .B(w_add_1_Z[4]), .C(n840), .D(r_add_1_B[4]), 
        .E(n839), .F(w_add_2_Z[4]), .G(r_x_data[132]), .H(n834), .Y(n687) );
  scg4d1_hd U1652 ( .A(n841), .B(w_add_1_Z[5]), .C(n840), .D(r_add_1_B[5]), 
        .E(n839), .F(w_add_2_Z[5]), .G(r_x_data[133]), .H(n832), .Y(n686) );
  scg4d1_hd U1653 ( .A(n841), .B(w_add_1_Z[6]), .C(n840), .D(r_add_1_B[6]), 
        .E(n839), .F(w_add_2_Z[6]), .G(r_x_data[134]), .H(n832), .Y(n685) );
  scg4d1_hd U1654 ( .A(n841), .B(w_add_1_Z[7]), .C(n840), .D(r_add_1_B[7]), 
        .E(n839), .F(w_add_2_Z[7]), .G(r_x_data[135]), .H(n832), .Y(n684) );
  scg4d1_hd U1655 ( .A(n841), .B(w_add_1_Z[8]), .C(n840), .D(r_add_1_B[8]), 
        .E(n839), .F(w_add_2_Z[8]), .G(r_x_data[136]), .H(n832), .Y(n683) );
  scg4d1_hd U1656 ( .A(n841), .B(w_add_1_Z[9]), .C(n840), .D(r_add_1_B[9]), 
        .E(n839), .F(w_add_2_Z[9]), .G(r_x_data[137]), .H(n830), .Y(n682) );
  scg4d1_hd U1657 ( .A(n841), .B(w_add_1_Z[10]), .C(n840), .D(r_add_1_B[10]), 
        .E(n839), .F(w_add_2_Z[10]), .G(r_x_data[138]), .H(n832), .Y(n681) );
  scg4d1_hd U1658 ( .A(n841), .B(w_add_1_Z[11]), .C(n840), .D(r_add_1_B[11]), 
        .E(n839), .F(w_add_2_Z[11]), .G(r_x_data[139]), .H(n830), .Y(n680) );
  scg4d1_hd U1659 ( .A(n841), .B(w_add_1_Z[12]), .C(n840), .D(r_add_1_B[12]), 
        .E(n839), .F(w_add_2_Z[12]), .G(r_x_data[140]), .H(n834), .Y(n679) );
  scg4d1_hd U1660 ( .A(n841), .B(w_add_1_Z[13]), .C(n840), .D(r_add_1_B[13]), 
        .E(n839), .F(w_add_2_Z[13]), .G(r_x_data[141]), .H(n830), .Y(n678) );
  scg4d1_hd U1661 ( .A(n841), .B(w_add_1_Z[14]), .C(n840), .D(r_add_1_B[14]), 
        .E(n839), .F(w_add_2_Z[14]), .G(r_x_data[142]), .H(n834), .Y(n677) );
  scg4d1_hd U1662 ( .A(n841), .B(w_add_1_Z[15]), .C(n840), .D(r_add_1_B[15]), 
        .E(n839), .F(w_add_2_Z[15]), .G(r_x_data[143]), .H(n830), .Y(n676) );
  scg4d1_hd U1663 ( .A(n841), .B(w_add_1_Z[16]), .C(n840), .D(r_add_1_B[16]), 
        .E(n839), .F(w_add_2_Z[16]), .G(r_x_data[144]), .H(n832), .Y(n675) );
  scg4d1_hd U1664 ( .A(n841), .B(w_add_1_Z[17]), .C(n840), .D(r_add_1_B[17]), 
        .E(n839), .F(w_add_2_Z[17]), .G(r_x_data[145]), .H(n834), .Y(n674) );
  scg4d1_hd U1665 ( .A(n841), .B(w_add_1_Z[18]), .C(n840), .D(r_add_1_B[18]), 
        .E(n839), .F(w_add_2_Z[18]), .G(r_x_data[146]), .H(n832), .Y(n673) );
  scg21d1_hd U1666 ( .A(r_counter_1_), .B(n506), .C(n1077), .D(n1035), .Y(
        n1036) );
  oa21d1_hd U1667 ( .A(N739), .B(n1037), .C(n1036), .Y(n1039) );
  ao211d1_hd U1668 ( .A(n829), .B(n1039), .C(n1038), .D(n5), .Y(n498) );
  ao22d1_hd U1669 ( .A(n548), .B(n1043), .C(n1041), .D(n1040), .Y(n496) );
  ao22d1_hd U1670 ( .A(n1043), .B(n1042), .C(n1041), .D(n1077), .Y(n494) );
  scg14d1_hd U1671 ( .A(r_x_data[31]), .B(n850), .C(n1044), .Y(n458) );
  scg14d1_hd U1672 ( .A(r_x_data[30]), .B(n833), .C(n1045), .Y(n459) );
  scg14d1_hd U1673 ( .A(r_x_data[29]), .B(n850), .C(n1046), .Y(n460) );
  scg14d1_hd U1674 ( .A(r_x_data[28]), .B(n833), .C(n1047), .Y(n461) );
  scg14d1_hd U1675 ( .A(r_x_data[27]), .B(n850), .C(n1048), .Y(n462) );
  scg14d1_hd U1676 ( .A(r_x_data[26]), .B(n833), .C(n1049), .Y(n463) );
  scg14d1_hd U1677 ( .A(r_x_data[25]), .B(n850), .C(n1050), .Y(n464) );
  scg14d1_hd U1678 ( .A(r_x_data[24]), .B(n833), .C(n1051), .Y(n465) );
  scg14d1_hd U1679 ( .A(r_x_data[23]), .B(n833), .C(n1052), .Y(n466) );
  scg14d1_hd U1680 ( .A(r_x_data[22]), .B(n828), .C(n1053), .Y(n467) );
  scg14d1_hd U1681 ( .A(r_x_data[21]), .B(n828), .C(n1054), .Y(n468) );
  scg14d1_hd U1682 ( .A(r_x_data[20]), .B(n828), .C(n1055), .Y(n469) );
  scg14d1_hd U1683 ( .A(r_x_data[19]), .B(n828), .C(n1056), .Y(n470) );
  scg14d1_hd U1684 ( .A(r_x_data[18]), .B(n828), .C(n1057), .Y(n471) );
  scg14d1_hd U1685 ( .A(r_x_data[17]), .B(n833), .C(n1058), .Y(n472) );
  scg14d1_hd U1686 ( .A(r_x_data[16]), .B(n828), .C(n1059), .Y(n473) );
  scg14d1_hd U1687 ( .A(r_x_data[15]), .B(n828), .C(n1060), .Y(n474) );
  scg14d1_hd U1688 ( .A(r_x_data[14]), .B(n828), .C(n1061), .Y(n475) );
  scg14d1_hd U1689 ( .A(r_x_data[13]), .B(n828), .C(n1062), .Y(n476) );
  scg14d1_hd U1690 ( .A(r_x_data[12]), .B(n850), .C(n1063), .Y(n477) );
  scg14d1_hd U1691 ( .A(r_x_data[11]), .B(n833), .C(n1064), .Y(n478) );
  scg14d1_hd U1692 ( .A(r_x_data[10]), .B(n828), .C(n1065), .Y(n479) );
  scg14d1_hd U1693 ( .A(r_x_data[9]), .B(n833), .C(n1066), .Y(n480) );
  scg14d1_hd U1694 ( .A(r_x_data[8]), .B(n833), .C(n1067), .Y(n481) );
  scg14d1_hd U1695 ( .A(r_x_data[7]), .B(n833), .C(n1068), .Y(n482) );
  scg14d1_hd U1696 ( .A(r_x_data[6]), .B(n833), .C(n1069), .Y(n483) );
  scg14d1_hd U1697 ( .A(r_x_data[5]), .B(n833), .C(n1070), .Y(n484) );
  scg14d1_hd U1698 ( .A(r_x_data[4]), .B(n833), .C(n1071), .Y(n485) );
  scg14d1_hd U1699 ( .A(r_x_data[3]), .B(n833), .C(n1072), .Y(n486) );
  scg14d1_hd U1700 ( .A(r_x_data[2]), .B(n833), .C(n1073), .Y(n487) );
  scg14d1_hd U1701 ( .A(r_x_data[1]), .B(n833), .C(n1074), .Y(n488) );
  scg14d1_hd U1702 ( .A(r_x_data[0]), .B(n833), .C(n1075), .Y(n489) );
endmodule

