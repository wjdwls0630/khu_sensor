
module converter_f2i ( i_A, i_A_STB, o_A_ACK, o_Z, o_Z_STB, i_Z_ACK, i_CLK, 
        i_RST );
  input [31:0] i_A;
  output [31:0] o_Z;
  input i_A_STB, i_Z_ACK, i_CLK, i_RST;
  output o_A_ACK, o_Z_STB;
  wire   a_s, N65, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         RSOP_38_C1_CONTROL1, n1, n88, n113, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470;
  wire   [2:0] state;
  wire   [31:0] a;
  wire   [8:0] a_e;
  wire   [31:1] a_m;
  wire   [31:0] z;

  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n1), .CK(i_CLK), .Q(o_Z[0]) );
  fd1qd1_hd z_reg_30_ ( .D(n142), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_29_ ( .D(n143), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_28_ ( .D(n144), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_27_ ( .D(n145), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_26_ ( .D(n146), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_25_ ( .D(n147), .CK(i_CLK), .Q(z[25]) );
  fd1qd1_hd z_reg_24_ ( .D(n148), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n149), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_22_ ( .D(n150), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd z_reg_21_ ( .D(n151), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n152), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n153), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n154), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_17_ ( .D(n155), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n156), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_15_ ( .D(n157), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n158), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_13_ ( .D(n159), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n160), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_11_ ( .D(n161), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n162), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_9_ ( .D(n163), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n164), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_7_ ( .D(n165), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n166), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_5_ ( .D(n167), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_4_ ( .D(n168), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_3_ ( .D(n169), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_2_ ( .D(n170), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_0_ ( .D(n172), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_31_ ( .D(n141), .CK(i_CLK), .Q(z[31]) );
  fd1qd1_hd z_reg_1_ ( .D(n171), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n140), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd o_A_ACK_reg ( .D(n208), .CK(i_CLK), .Q(o_A_ACK) );
  fd1qd1_hd a_m_reg_31_ ( .D(n204), .CK(i_CLK), .Q(a_m[31]) );
  fd1qd1_hd a_m_reg_30_ ( .D(n173), .CK(i_CLK), .Q(a_m[30]) );
  fd1eqd1_hd a_e_reg_3_ ( .D(N177), .E(n88), .CK(i_CLK), .Q(a_e[3]) );
  fd1eqd1_hd a_e_reg_8_ ( .D(N182), .E(n88), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_0_ ( .D(n206), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd state_reg_2_ ( .D(n207), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_1_ ( .D(n205), .CK(i_CLK), .Q(state[1]) );
  fd1eqd1_hd a_e_reg_6_ ( .D(N180), .E(n88), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd a_m_reg_28_ ( .D(n175), .CK(i_CLK), .Q(a_m[28]) );
  fd1qd1_hd a_m_reg_26_ ( .D(n177), .CK(i_CLK), .Q(a_m[26]) );
  fd1eqd1_hd a_e_reg_0_ ( .D(N174), .E(n88), .CK(i_CLK), .Q(a_e[0]) );
  fd1eqd1_hd a_e_reg_4_ ( .D(N178), .E(n88), .CK(i_CLK), .Q(a_e[4]) );
  fd1eqd1_hd a_e_reg_2_ ( .D(N176), .E(n88), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd a_e_reg_1_ ( .D(N175), .E(n88), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_m_reg_29_ ( .D(n174), .CK(i_CLK), .Q(a_m[29]) );
  fd1qd1_hd a_m_reg_27_ ( .D(n176), .CK(i_CLK), .Q(a_m[27]) );
  fd1eqd1_hd a_e_reg_5_ ( .D(N179), .E(n88), .CK(i_CLK), .Q(a_e[5]) );
  fd1eqd1_hd a_e_reg_7_ ( .D(N181), .E(n88), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n179), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n181), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n183), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd a_m_reg_25_ ( .D(n178), .CK(i_CLK), .Q(a_m[25]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n180), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n182), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n185), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n187), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n184), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n186), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n189), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n191), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n193), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n188), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n190), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n192), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n197), .CK(i_CLK), .Q(a_m[6]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n195), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n196), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n194), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n199), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n201), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n202), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n198), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n200), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n203), .CK(i_CLK), .Q(N65) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n1), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n113), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n113), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n113), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n113), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n113), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n113), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n113), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n113), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n113), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n113), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n113), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n113), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n113), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n113), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n113), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n113), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n113), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n214), .CK(i_CLK), .Q(a_s) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n113), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n113), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n113), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n113), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n113), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n113), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n113), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n113), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n113), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n113), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n113), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n113), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n113), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n113), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n113), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n1), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n1), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n1), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n1), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n1), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n1), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n1), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n1), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n1), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n1), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n1), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n1), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n1), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n1), .CK(i_CLK), .Q(o_Z[1]) );
  clknd2d1_hd U223 ( .A(a[23]), .B(a[24]), .Y(n467) );
  clknd2d1_hd U224 ( .A(n453), .B(a_e[4]), .Y(n448) );
  clknd2d1_hd U225 ( .A(n444), .B(a_e[5]), .Y(n443) );
  clknd2d1_hd U226 ( .A(n449), .B(a[28]), .Y(n445) );
  clknd2d1_hd U227 ( .A(n427), .B(n237), .Y(n233) );
  clknd2d1_hd U228 ( .A(a_e[7]), .B(n438), .Y(n433) );
  clknd2d1_hd U229 ( .A(n220), .B(n448), .Y(n221) );
  clknd2d1_hd U230 ( .A(state[1]), .B(n225), .Y(n227) );
  clknd2d1_hd U231 ( .A(n461), .B(a[26]), .Y(n455) );
  clknd2d1_hd U232 ( .A(n427), .B(n215), .Y(n222) );
  clknd2d1_hd U233 ( .A(state[0]), .B(n219), .Y(n419) );
  clknd2d1_hd U234 ( .A(a_s), .B(n212), .Y(n424) );
  clknd2d1_hd U235 ( .A(n284), .B(n238), .Y(n285) );
  clknd2d1_hd U236 ( .A(n290), .B(n239), .Y(n294) );
  clknd2d1_hd U237 ( .A(n299), .B(n240), .Y(n303) );
  clknd2d1_hd U238 ( .A(n308), .B(n241), .Y(n312) );
  clknd2d1_hd U239 ( .A(n317), .B(n243), .Y(n321) );
  clknd2d1_hd U240 ( .A(n326), .B(n246), .Y(n330) );
  clknd2d1_hd U241 ( .A(n335), .B(n249), .Y(n339) );
  clknd2d1_hd U242 ( .A(n344), .B(n252), .Y(n348) );
  clknd2d1_hd U243 ( .A(n353), .B(n255), .Y(n357) );
  clknd2d1_hd U244 ( .A(n362), .B(n258), .Y(n366) );
  clknd2d1_hd U245 ( .A(n371), .B(n261), .Y(n375) );
  clknd2d1_hd U246 ( .A(n380), .B(n264), .Y(n384) );
  clknd2d1_hd U247 ( .A(n389), .B(n267), .Y(n393) );
  clknd2d1_hd U248 ( .A(n398), .B(n270), .Y(n402) );
  nid1_hd U249 ( .A(n414), .Y(n212) );
  clknd2d1_hd U250 ( .A(n407), .B(n273), .Y(n412) );
  clknd2d1_hd U251 ( .A(n418), .B(n422), .Y(n280) );
  clknd2d1_hd U252 ( .A(n432), .B(a[30]), .Y(n436) );
  clknd2d1_hd U253 ( .A(n447), .B(n446), .Y(N179) );
  clknd2d1_hd U254 ( .A(n464), .B(n463), .Y(N176) );
  clknd2d1_hd U255 ( .A(n452), .B(n451), .Y(N178) );
  clknd2d1_hd U256 ( .A(n445), .B(n437), .Y(n441) );
  clknd2d1_hd U257 ( .A(n214), .B(n427), .Y(n230) );
  clknd2d1_hd U258 ( .A(n434), .B(n431), .Y(N182) );
  clknd2d1_hd U259 ( .A(n430), .B(n433), .Y(n429) );
  clknd2d1_hd U260 ( .A(n457), .B(n456), .Y(N177) );
  clknd2d1_hd U261 ( .A(n212), .B(n408), .Y(n281) );
  clknd2d1_hd U262 ( .A(n288), .B(n287), .Y(n286) );
  clknd2d1_hd U263 ( .A(a_s), .B(n285), .Y(n287) );
  clknd2d1_hd U264 ( .A(a_m[3]), .B(n292), .Y(n291) );
  clknd2d1_hd U265 ( .A(n297), .B(n296), .Y(n295) );
  clknd2d1_hd U266 ( .A(a_s), .B(n294), .Y(n296) );
  clknd2d1_hd U267 ( .A(a_m[5]), .B(n301), .Y(n300) );
  clknd2d1_hd U268 ( .A(n306), .B(n305), .Y(n304) );
  clknd2d1_hd U269 ( .A(a_s), .B(n303), .Y(n305) );
  clknd2d1_hd U270 ( .A(a_m[7]), .B(n310), .Y(n309) );
  clknd2d1_hd U271 ( .A(n315), .B(n314), .Y(n313) );
  clknd2d1_hd U272 ( .A(a_s), .B(n312), .Y(n314) );
  clknd2d1_hd U273 ( .A(a_m[9]), .B(n319), .Y(n318) );
  clknd2d1_hd U274 ( .A(n324), .B(n323), .Y(n322) );
  clknd2d1_hd U275 ( .A(a_s), .B(n321), .Y(n323) );
  clknd2d1_hd U276 ( .A(a_m[11]), .B(n328), .Y(n327) );
  clknd2d1_hd U277 ( .A(n333), .B(n332), .Y(n331) );
  clknd2d1_hd U278 ( .A(a_s), .B(n330), .Y(n332) );
  clknd2d1_hd U279 ( .A(a_m[13]), .B(n337), .Y(n336) );
  clknd2d1_hd U280 ( .A(n342), .B(n341), .Y(n340) );
  clknd2d1_hd U281 ( .A(a_s), .B(n339), .Y(n341) );
  clknd2d1_hd U282 ( .A(a_m[15]), .B(n346), .Y(n345) );
  clknd2d1_hd U283 ( .A(n351), .B(n350), .Y(n349) );
  clknd2d1_hd U284 ( .A(a_s), .B(n348), .Y(n350) );
  clknd2d1_hd U285 ( .A(a_m[17]), .B(n355), .Y(n354) );
  clknd2d1_hd U286 ( .A(n360), .B(n359), .Y(n358) );
  clknd2d1_hd U287 ( .A(a_s), .B(n357), .Y(n359) );
  clknd2d1_hd U288 ( .A(a_m[19]), .B(n364), .Y(n363) );
  clknd2d1_hd U289 ( .A(n369), .B(n368), .Y(n367) );
  clknd2d1_hd U290 ( .A(a_s), .B(n366), .Y(n368) );
  clknd2d1_hd U291 ( .A(a_m[21]), .B(n373), .Y(n372) );
  clknd2d1_hd U292 ( .A(n378), .B(n377), .Y(n376) );
  clknd2d1_hd U293 ( .A(a_s), .B(n375), .Y(n377) );
  clknd2d1_hd U294 ( .A(a_m[23]), .B(n382), .Y(n381) );
  clknd2d1_hd U295 ( .A(n387), .B(n386), .Y(n385) );
  clknd2d1_hd U296 ( .A(a_s), .B(n384), .Y(n386) );
  clknd2d1_hd U297 ( .A(a_m[25]), .B(n391), .Y(n390) );
  clknd2d1_hd U298 ( .A(n396), .B(n395), .Y(n394) );
  clknd2d1_hd U299 ( .A(a_s), .B(n393), .Y(n395) );
  clknd2d1_hd U300 ( .A(a_m[27]), .B(n400), .Y(n399) );
  clknd2d1_hd U301 ( .A(n405), .B(n404), .Y(n403) );
  clknd2d1_hd U302 ( .A(a_s), .B(n402), .Y(n404) );
  clknd2d1_hd U303 ( .A(a_m[29]), .B(n410), .Y(n409) );
  clknd2d1_hd U304 ( .A(n416), .B(n415), .Y(n413) );
  clknd2d1_hd U305 ( .A(a_s), .B(n412), .Y(n415) );
  ivd4_hd U306 ( .A(n215), .Y(n113) );
  nr2d4_hd U307 ( .A(n225), .B(n223), .Y(n1) );
  clknd2d1_hd U308 ( .A(n236), .B(n231), .Y(n223) );
  scg2d1_hd U309 ( .A(N65), .B(n212), .C(n213), .D(z[0]), .Y(n172) );
  nr2d2_hd U310 ( .A(n470), .B(n280), .Y(n414) );
  or2d1_hd U311 ( .A(n279), .B(n278), .Y(n422) );
  or2d1_hd U312 ( .A(state[0]), .B(n227), .Y(RSOP_38_C1_CONTROL1) );
  or2d1_hd U313 ( .A(a_e[5]), .B(a_e[6]), .Y(n218) );
  nid2_hd U314 ( .A(n277), .Y(n211) );
  ivd1_hd U315 ( .A(a_m[1]), .Y(n284) );
  ivd2_hd U316 ( .A(n88), .Y(n275) );
  nd2d1_hd U317 ( .A(n459), .B(n88), .Y(n277) );
  scg20d2_hd U318 ( .A(n228), .B(n231), .C(n227), .Y(n88) );
  ivd2_hd U319 ( .A(n422), .Y(n213) );
  nr2d1_hd U320 ( .A(a_m[30]), .B(n412), .Y(n425) );
  nr2d1_hd U321 ( .A(a_m[28]), .B(n402), .Y(n407) );
  nr2d1_hd U322 ( .A(a_m[26]), .B(n393), .Y(n398) );
  nr2d1_hd U323 ( .A(a_m[24]), .B(n384), .Y(n389) );
  nr2d1_hd U324 ( .A(a_m[22]), .B(n375), .Y(n380) );
  nr2d1_hd U325 ( .A(a_m[20]), .B(n366), .Y(n371) );
  nr2d1_hd U326 ( .A(a_m[18]), .B(n357), .Y(n362) );
  nr2d1_hd U327 ( .A(a_m[16]), .B(n348), .Y(n353) );
  nr2d1_hd U328 ( .A(a_m[14]), .B(n339), .Y(n344) );
  nr2d1_hd U329 ( .A(a_m[12]), .B(n330), .Y(n335) );
  nr2d1_hd U330 ( .A(a_m[10]), .B(n321), .Y(n326) );
  nr2d1_hd U331 ( .A(a_m[8]), .B(n312), .Y(n317) );
  nr2d1_hd U332 ( .A(a_m[6]), .B(n303), .Y(n308) );
  nr2d1_hd U333 ( .A(a_m[4]), .B(n294), .Y(n299) );
  ivd1_hd U334 ( .A(a_m[3]), .Y(n239) );
  ivd1_hd U335 ( .A(N65), .Y(n238) );
  nr2d1_hd U336 ( .A(n228), .B(n470), .Y(n279) );
  ao22d1_hd U337 ( .A(n425), .B(n418), .C(n430), .D(n221), .Y(n228) );
  ivd1_hd U338 ( .A(a_m[7]), .Y(n241) );
  ivd1_hd U339 ( .A(a_m[5]), .Y(n240) );
  nr2d1_hd U340 ( .A(a_m[2]), .B(n285), .Y(n290) );
  ivd1_hd U341 ( .A(n459), .Y(n470) );
  nr2d1_hd U342 ( .A(n227), .B(n231), .Y(n459) );
  ivd2_hd U343 ( .A(RSOP_38_C1_CONTROL1), .Y(n214) );
  ivd1_hd U344 ( .A(a_s), .Y(n408) );
  scg20d1_hd U345 ( .A(a_e[8]), .B(n220), .C(n420), .Y(n229) );
  nr2d1_hd U346 ( .A(n458), .B(n454), .Y(n453) );
  ivd1_hd U347 ( .A(a_e[3]), .Y(n454) );
  ivd1_hd U348 ( .A(a_e[8]), .Y(n430) );
  ivd1_hd U349 ( .A(a_m[29]), .Y(n273) );
  ivd1_hd U350 ( .A(a_m[27]), .Y(n270) );
  ivd1_hd U351 ( .A(a_m[25]), .Y(n267) );
  ivd1_hd U352 ( .A(a_m[23]), .Y(n264) );
  ivd1_hd U353 ( .A(a_m[21]), .Y(n261) );
  ivd1_hd U354 ( .A(a_m[19]), .Y(n258) );
  ivd1_hd U355 ( .A(a_m[17]), .Y(n255) );
  ivd1_hd U356 ( .A(a_m[15]), .Y(n252) );
  ivd1_hd U357 ( .A(a_m[13]), .Y(n249) );
  ivd1_hd U358 ( .A(a_m[11]), .Y(n246) );
  ivd1_hd U359 ( .A(a_m[31]), .Y(n418) );
  ivd1_hd U360 ( .A(state[0]), .Y(n231) );
  ivd1_hd U361 ( .A(state[2]), .Y(n225) );
  scg6d1_hd U362 ( .A(n442), .B(n441), .C(n440), .Y(N180) );
  ivd1_hd U363 ( .A(a[29]), .Y(n437) );
  nd3d1_hd U364 ( .A(n232), .B(i_A_STB), .C(o_A_ACK), .Y(n215) );
  scg14d1_hd U365 ( .A(n213), .B(z[24]), .C(n388), .Y(n148) );
  ivd1_hd U366 ( .A(a_m[24]), .Y(n387) );
  scg14d1_hd U367 ( .A(n213), .B(z[20]), .C(n370), .Y(n152) );
  ivd1_hd U368 ( .A(a_m[20]), .Y(n369) );
  scg14d1_hd U369 ( .A(n213), .B(z[18]), .C(n361), .Y(n154) );
  ivd1_hd U370 ( .A(a_m[18]), .Y(n360) );
  scg14d1_hd U371 ( .A(n213), .B(z[6]), .C(n307), .Y(n166) );
  scg14d1_hd U372 ( .A(n213), .B(z[22]), .C(n379), .Y(n150) );
  ivd1_hd U373 ( .A(a_m[22]), .Y(n378) );
  ivd1_hd U374 ( .A(a_m[6]), .Y(n306) );
  scg14d1_hd U375 ( .A(n213), .B(z[9]), .C(n320), .Y(n163) );
  scg14d1_hd U376 ( .A(n213), .B(z[26]), .C(n397), .Y(n146) );
  ivd1_hd U377 ( .A(a_m[26]), .Y(n396) );
  scg14d1_hd U378 ( .A(n213), .B(z[12]), .C(n334), .Y(n160) );
  ivd1_hd U379 ( .A(a_m[12]), .Y(n333) );
  scg14d1_hd U380 ( .A(n213), .B(z[14]), .C(n343), .Y(n158) );
  ivd1_hd U381 ( .A(a_m[14]), .Y(n342) );
  scg14d1_hd U382 ( .A(n213), .B(z[28]), .C(n406), .Y(n144) );
  ivd1_hd U383 ( .A(a_m[28]), .Y(n405) );
  scg14d1_hd U384 ( .A(n213), .B(z[10]), .C(n325), .Y(n162) );
  ivd1_hd U385 ( .A(a_m[10]), .Y(n324) );
  scg14d1_hd U386 ( .A(n213), .B(z[16]), .C(n352), .Y(n156) );
  ivd1_hd U387 ( .A(a_m[16]), .Y(n351) );
  scg14d1_hd U388 ( .A(n213), .B(z[8]), .C(n316), .Y(n164) );
  ivd1_hd U389 ( .A(a_m[8]), .Y(n315) );
  scg14d1_hd U390 ( .A(n213), .B(z[30]), .C(n417), .Y(n142) );
  ivd1_hd U391 ( .A(a_m[30]), .Y(n416) );
  scg14d1_hd U392 ( .A(n213), .B(z[27]), .C(n401), .Y(n145) );
  scg14d1_hd U393 ( .A(n213), .B(z[4]), .C(n298), .Y(n168) );
  ivd1_hd U394 ( .A(a_m[4]), .Y(n297) );
  scg14d1_hd U395 ( .A(n213), .B(z[2]), .C(n289), .Y(n170) );
  ivd1_hd U396 ( .A(a_m[2]), .Y(n288) );
  scg14d1_hd U397 ( .A(n213), .B(z[29]), .C(n411), .Y(n143) );
  nr2d1_hd U398 ( .A(n229), .B(n419), .Y(n278) );
  ivd1_hd U399 ( .A(a_e[0]), .Y(n466) );
  nr3d1_hd U400 ( .A(a_e[7]), .B(a_e[5]), .C(a_e[6]), .Y(n220) );
  ivd1_hd U401 ( .A(a_m[9]), .Y(n243) );
  nd2bd1_hd U402 ( .AN(a[30]), .B(n442), .Y(n434) );
  nr2d1_hd U403 ( .A(state[2]), .B(n223), .Y(n232) );
  ivd1_hd U404 ( .A(state[1]), .Y(n236) );
  nr2d1_hd U405 ( .A(state[2]), .B(state[1]), .Y(n219) );
  ivd1_hd U406 ( .A(i_RST), .Y(n427) );
  scg20d1_hd U407 ( .A(n232), .B(o_A_ACK), .C(n222), .Y(n208) );
  nr2d1_hd U408 ( .A(a_e[1]), .B(n466), .Y(n465) );
  ivd1_hd U409 ( .A(a_e[4]), .Y(n216) );
  nd4d1_hd U410 ( .A(a_e[8]), .B(a_e[7]), .C(n465), .D(n216), .Y(n217) );
  nr4d1_hd U411 ( .A(a_e[2]), .B(a_e[3]), .C(n218), .D(n217), .Y(n420) );
  nr2d1_hd U412 ( .A(n459), .B(n278), .Y(n226) );
  nd3d1_hd U413 ( .A(a_e[0]), .B(a_e[1]), .C(a_e[2]), .Y(n458) );
  nr2d1_hd U414 ( .A(n279), .B(n222), .Y(n224) );
  nd3d1_hd U415 ( .A(n1), .B(i_Z_ACK), .C(o_Z_STB), .Y(n426) );
  nd4d1_hd U416 ( .A(n224), .B(n419), .C(n426), .D(RSOP_38_C1_CONTROL1), .Y(
        n237) );
  oa22d1_hd U417 ( .A(n226), .B(n233), .C(n225), .D(n237), .Y(n207) );
  scg13d1_hd U418 ( .A(n419), .B(i_RST), .C(n229), .Y(n235) );
  oa211d1_hd U419 ( .A(n237), .B(n231), .C(n235), .D(n230), .Y(n206) );
  nd2bd1_hd U420 ( .AN(n233), .B(n232), .Y(n234) );
  oa211d1_hd U421 ( .A(n237), .B(n236), .C(n235), .D(n234), .Y(n205) );
  oa21d1_hd U422 ( .A(n418), .B(n88), .C(RSOP_38_C1_CONTROL1), .Y(n204) );
  oa22d1_hd U423 ( .A(n284), .B(n277), .C(n238), .D(n88), .Y(n203) );
  oa22d1_hd U424 ( .A(n284), .B(n88), .C(n288), .D(n211), .Y(n202) );
  oa22d1_hd U425 ( .A(n239), .B(n277), .C(n288), .D(n88), .Y(n201) );
  oa22d1_hd U426 ( .A(n297), .B(n211), .C(n239), .D(n88), .Y(n200) );
  oa22d1_hd U427 ( .A(n240), .B(n277), .C(n297), .D(n88), .Y(n199) );
  oa22d1_hd U428 ( .A(n306), .B(n211), .C(n240), .D(n88), .Y(n198) );
  oa22d1_hd U429 ( .A(n241), .B(n211), .C(n306), .D(n88), .Y(n197) );
  oa22d1_hd U430 ( .A(n315), .B(n211), .C(n241), .D(n88), .Y(n196) );
  ao22d1_hd U431 ( .A(a_m[8]), .B(n275), .C(n214), .D(a[0]), .Y(n242) );
  oa21d1_hd U432 ( .A(n243), .B(n211), .C(n242), .Y(n195) );
  ao22d1_hd U433 ( .A(a_m[9]), .B(n275), .C(n214), .D(a[1]), .Y(n244) );
  oa21d1_hd U434 ( .A(n324), .B(n211), .C(n244), .Y(n194) );
  ao22d1_hd U435 ( .A(a_m[10]), .B(n275), .C(n214), .D(a[2]), .Y(n245) );
  oa21d1_hd U436 ( .A(n246), .B(n211), .C(n245), .Y(n193) );
  ao22d1_hd U437 ( .A(a_m[11]), .B(n275), .C(n214), .D(a[3]), .Y(n247) );
  oa21d1_hd U438 ( .A(n333), .B(n211), .C(n247), .Y(n192) );
  ao22d1_hd U439 ( .A(a_m[12]), .B(n275), .C(n214), .D(a[4]), .Y(n248) );
  oa21d1_hd U440 ( .A(n249), .B(n211), .C(n248), .Y(n191) );
  ao22d1_hd U441 ( .A(a_m[13]), .B(n275), .C(n214), .D(a[5]), .Y(n250) );
  oa21d1_hd U442 ( .A(n342), .B(n211), .C(n250), .Y(n190) );
  ao22d1_hd U443 ( .A(a_m[14]), .B(n275), .C(n214), .D(a[6]), .Y(n251) );
  oa21d1_hd U444 ( .A(n252), .B(n211), .C(n251), .Y(n189) );
  ao22d1_hd U445 ( .A(a_m[15]), .B(n275), .C(n214), .D(a[7]), .Y(n253) );
  oa21d1_hd U446 ( .A(n351), .B(n211), .C(n253), .Y(n188) );
  ao22d1_hd U447 ( .A(a_m[16]), .B(n275), .C(n214), .D(a[8]), .Y(n254) );
  oa21d1_hd U448 ( .A(n255), .B(n211), .C(n254), .Y(n187) );
  ao22d1_hd U449 ( .A(a_m[17]), .B(n275), .C(n214), .D(a[9]), .Y(n256) );
  oa21d1_hd U450 ( .A(n360), .B(n277), .C(n256), .Y(n186) );
  ao22d1_hd U451 ( .A(a_m[18]), .B(n275), .C(n214), .D(a[10]), .Y(n257) );
  oa21d1_hd U452 ( .A(n258), .B(n277), .C(n257), .Y(n185) );
  ao22d1_hd U453 ( .A(a_m[19]), .B(n275), .C(n214), .D(a[11]), .Y(n259) );
  oa21d1_hd U454 ( .A(n369), .B(n277), .C(n259), .Y(n184) );
  ao22d1_hd U455 ( .A(a_m[20]), .B(n275), .C(n214), .D(a[12]), .Y(n260) );
  oa21d1_hd U456 ( .A(n261), .B(n277), .C(n260), .Y(n183) );
  ao22d1_hd U457 ( .A(a_m[21]), .B(n275), .C(n214), .D(a[13]), .Y(n262) );
  oa21d1_hd U458 ( .A(n378), .B(n277), .C(n262), .Y(n182) );
  ao22d1_hd U459 ( .A(a_m[22]), .B(n275), .C(n214), .D(a[14]), .Y(n263) );
  oa21d1_hd U460 ( .A(n264), .B(n277), .C(n263), .Y(n181) );
  ao22d1_hd U461 ( .A(a_m[23]), .B(n275), .C(n214), .D(a[15]), .Y(n265) );
  oa21d1_hd U462 ( .A(n387), .B(n277), .C(n265), .Y(n180) );
  ao22d1_hd U463 ( .A(a_m[24]), .B(n275), .C(n214), .D(a[16]), .Y(n266) );
  oa21d1_hd U464 ( .A(n267), .B(n211), .C(n266), .Y(n179) );
  ao22d1_hd U465 ( .A(a_m[25]), .B(n275), .C(n214), .D(a[17]), .Y(n268) );
  oa21d1_hd U466 ( .A(n396), .B(n277), .C(n268), .Y(n178) );
  ao22d1_hd U467 ( .A(a_m[26]), .B(n275), .C(n214), .D(a[18]), .Y(n269) );
  oa21d1_hd U468 ( .A(n270), .B(n211), .C(n269), .Y(n177) );
  ao22d1_hd U469 ( .A(a_m[27]), .B(n275), .C(n214), .D(a[19]), .Y(n271) );
  oa21d1_hd U470 ( .A(n405), .B(n277), .C(n271), .Y(n176) );
  ao22d1_hd U471 ( .A(a_m[28]), .B(n275), .C(n214), .D(a[20]), .Y(n272) );
  oa21d1_hd U472 ( .A(n273), .B(n211), .C(n272), .Y(n175) );
  ao22d1_hd U473 ( .A(a_m[29]), .B(n275), .C(n214), .D(a[21]), .Y(n274) );
  oa21d1_hd U474 ( .A(n416), .B(n277), .C(n274), .Y(n174) );
  ao22d1_hd U475 ( .A(a_m[30]), .B(n275), .C(n214), .D(a[22]), .Y(n276) );
  oa21d1_hd U476 ( .A(n418), .B(n211), .C(n276), .Y(n173) );
  oa21d1_hd U477 ( .A(N65), .B(n424), .C(n281), .Y(n282) );
  ao22d1_hd U478 ( .A(a_m[1]), .B(n282), .C(n213), .D(z[1]), .Y(n283) );
  scg22d1_hd U479 ( .A(N65), .B(n284), .C(n424), .D(n283), .Y(n171) );
  oa211d1_hd U480 ( .A(n288), .B(n287), .C(n212), .D(n286), .Y(n289) );
  nr2d1_hd U481 ( .A(n408), .B(n290), .Y(n292) );
  oa211d1_hd U482 ( .A(a_m[3]), .B(n292), .C(n212), .D(n291), .Y(n293) );
  scg14d1_hd U483 ( .A(n213), .B(z[3]), .C(n293), .Y(n169) );
  oa211d1_hd U484 ( .A(n297), .B(n296), .C(n212), .D(n295), .Y(n298) );
  nr2d1_hd U485 ( .A(n408), .B(n299), .Y(n301) );
  oa211d1_hd U486 ( .A(a_m[5]), .B(n301), .C(n212), .D(n300), .Y(n302) );
  scg14d1_hd U487 ( .A(n213), .B(z[5]), .C(n302), .Y(n167) );
  oa211d1_hd U488 ( .A(n306), .B(n305), .C(n414), .D(n304), .Y(n307) );
  nr2d1_hd U489 ( .A(n408), .B(n308), .Y(n310) );
  oa211d1_hd U490 ( .A(a_m[7]), .B(n310), .C(n414), .D(n309), .Y(n311) );
  scg14d1_hd U491 ( .A(n213), .B(z[7]), .C(n311), .Y(n165) );
  oa211d1_hd U492 ( .A(n315), .B(n314), .C(n414), .D(n313), .Y(n316) );
  nr2d1_hd U493 ( .A(n408), .B(n317), .Y(n319) );
  oa211d1_hd U494 ( .A(a_m[9]), .B(n319), .C(n414), .D(n318), .Y(n320) );
  oa211d1_hd U495 ( .A(n324), .B(n323), .C(n414), .D(n322), .Y(n325) );
  nr2d1_hd U496 ( .A(n408), .B(n326), .Y(n328) );
  oa211d1_hd U497 ( .A(a_m[11]), .B(n328), .C(n414), .D(n327), .Y(n329) );
  scg14d1_hd U498 ( .A(n213), .B(z[11]), .C(n329), .Y(n161) );
  oa211d1_hd U499 ( .A(n333), .B(n332), .C(n414), .D(n331), .Y(n334) );
  nr2d1_hd U500 ( .A(n408), .B(n335), .Y(n337) );
  oa211d1_hd U501 ( .A(a_m[13]), .B(n337), .C(n414), .D(n336), .Y(n338) );
  scg14d1_hd U502 ( .A(n213), .B(z[13]), .C(n338), .Y(n159) );
  oa211d1_hd U503 ( .A(n342), .B(n341), .C(n414), .D(n340), .Y(n343) );
  nr2d1_hd U504 ( .A(n408), .B(n344), .Y(n346) );
  oa211d1_hd U505 ( .A(a_m[15]), .B(n346), .C(n414), .D(n345), .Y(n347) );
  scg14d1_hd U506 ( .A(n213), .B(z[15]), .C(n347), .Y(n157) );
  oa211d1_hd U507 ( .A(n351), .B(n350), .C(n414), .D(n349), .Y(n352) );
  nr2d1_hd U508 ( .A(n408), .B(n353), .Y(n355) );
  oa211d1_hd U509 ( .A(a_m[17]), .B(n355), .C(n212), .D(n354), .Y(n356) );
  scg14d1_hd U510 ( .A(n213), .B(z[17]), .C(n356), .Y(n155) );
  oa211d1_hd U511 ( .A(n360), .B(n359), .C(n414), .D(n358), .Y(n361) );
  nr2d1_hd U512 ( .A(n408), .B(n362), .Y(n364) );
  oa211d1_hd U513 ( .A(a_m[19]), .B(n364), .C(n212), .D(n363), .Y(n365) );
  scg14d1_hd U514 ( .A(n213), .B(z[19]), .C(n365), .Y(n153) );
  oa211d1_hd U515 ( .A(n369), .B(n368), .C(n414), .D(n367), .Y(n370) );
  nr2d1_hd U516 ( .A(n408), .B(n371), .Y(n373) );
  oa211d1_hd U517 ( .A(a_m[21]), .B(n373), .C(n212), .D(n372), .Y(n374) );
  scg14d1_hd U518 ( .A(n213), .B(z[21]), .C(n374), .Y(n151) );
  oa211d1_hd U519 ( .A(n378), .B(n377), .C(n414), .D(n376), .Y(n379) );
  nr2d1_hd U520 ( .A(n408), .B(n380), .Y(n382) );
  oa211d1_hd U521 ( .A(a_m[23]), .B(n382), .C(n212), .D(n381), .Y(n383) );
  scg14d1_hd U522 ( .A(n213), .B(z[23]), .C(n383), .Y(n149) );
  oa211d1_hd U523 ( .A(n387), .B(n386), .C(n414), .D(n385), .Y(n388) );
  nr2d1_hd U524 ( .A(n408), .B(n389), .Y(n391) );
  oa211d1_hd U525 ( .A(a_m[25]), .B(n391), .C(n212), .D(n390), .Y(n392) );
  scg14d1_hd U526 ( .A(n213), .B(z[25]), .C(n392), .Y(n147) );
  oa211d1_hd U527 ( .A(n396), .B(n395), .C(n414), .D(n394), .Y(n397) );
  nr2d1_hd U528 ( .A(n408), .B(n398), .Y(n400) );
  oa211d1_hd U529 ( .A(a_m[27]), .B(n400), .C(n212), .D(n399), .Y(n401) );
  oa211d1_hd U530 ( .A(n405), .B(n404), .C(n414), .D(n403), .Y(n406) );
  nr2d1_hd U531 ( .A(n408), .B(n407), .Y(n410) );
  oa211d1_hd U532 ( .A(a_m[29]), .B(n410), .C(n212), .D(n409), .Y(n411) );
  oa211d1_hd U533 ( .A(n416), .B(n415), .C(n414), .D(n413), .Y(n417) );
  oa22d1_hd U534 ( .A(n420), .B(n419), .C(n470), .D(n418), .Y(n421) );
  ao22d1_hd U535 ( .A(n213), .B(z[31]), .C(n421), .D(n422), .Y(n423) );
  oa21d1_hd U536 ( .A(n425), .B(n424), .C(n423), .Y(n141) );
  oa211d1_hd U537 ( .A(n1), .B(o_Z_STB), .C(n427), .D(n426), .Y(n428) );
  ivd1_hd U538 ( .A(n428), .Y(n140) );
  ivd1_hd U539 ( .A(a[25]), .Y(n462) );
  nr2d1_hd U540 ( .A(n467), .B(n462), .Y(n461) );
  ivd1_hd U541 ( .A(a[27]), .Y(n450) );
  nr2d1_hd U542 ( .A(n455), .B(n450), .Y(n449) );
  nr2d1_hd U543 ( .A(n445), .B(n437), .Y(n432) );
  nr2d1_hd U544 ( .A(n432), .B(RSOP_38_C1_CONTROL1), .Y(n442) );
  ivd1_hd U545 ( .A(a_e[6]), .Y(n439) );
  ivd1_hd U546 ( .A(n448), .Y(n444) );
  nr2d1_hd U547 ( .A(n439), .B(n443), .Y(n438) );
  oa211d1_hd U548 ( .A(n430), .B(n433), .C(n459), .D(n429), .Y(n431) );
  oa211d1_hd U549 ( .A(a_e[7]), .B(n438), .C(n459), .D(n433), .Y(n435) );
  oa211d1_hd U550 ( .A(RSOP_38_C1_CONTROL1), .B(n436), .C(n435), .D(n434), .Y(
        N181) );
  ao211d1_hd U551 ( .A(n439), .B(n443), .C(n438), .D(n470), .Y(n440) );
  oa211d1_hd U552 ( .A(n444), .B(a_e[5]), .C(n459), .D(n443), .Y(n447) );
  oa211d1_hd U553 ( .A(n449), .B(a[28]), .C(n214), .D(n445), .Y(n446) );
  oa211d1_hd U554 ( .A(n453), .B(a_e[4]), .C(n459), .D(n448), .Y(n452) );
  scg17d1_hd U555 ( .A(n455), .B(n450), .C(n449), .D(n214), .Y(n451) );
  scg17d1_hd U556 ( .A(n458), .B(n454), .C(n453), .D(n459), .Y(n457) );
  oa211d1_hd U557 ( .A(n461), .B(a[26]), .C(n214), .D(n455), .Y(n456) );
  nr2bd1_hd U558 ( .AN(a_e[1]), .B(n466), .Y(n460) );
  oa211d1_hd U559 ( .A(n460), .B(a_e[2]), .C(n459), .D(n458), .Y(n464) );
  scg17d1_hd U560 ( .A(n467), .B(n462), .C(n461), .D(n214), .Y(n463) );
  ao21d1_hd U561 ( .A(a_e[1]), .B(n466), .C(n465), .Y(n469) );
  oa211d1_hd U562 ( .A(a[23]), .B(a[24]), .C(n214), .D(n467), .Y(n468) );
  oa21d1_hd U563 ( .A(n469), .B(n470), .C(n468), .Y(N175) );
  oa22d1_hd U564 ( .A(a_e[0]), .B(n470), .C(a[23]), .D(RSOP_38_C1_CONTROL1), 
        .Y(N174) );
endmodule

