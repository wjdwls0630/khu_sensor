
module float_multiplier ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N34, a_s, b_s, N35, round_bit, sticky, z_s, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201,
         N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212,
         N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         C82_DATA2_1, C82_DATA2_2, C82_DATA2_3, C82_DATA2_4, C82_DATA2_5,
         C82_DATA2_6, C81_DATA2_1, C81_DATA2_2, C81_DATA2_3, C81_DATA2_4,
         C81_DATA2_5, C81_DATA2_6, net908, n10, n14, n20, n29, n34, n36, n104,
         n105, n110, n138, n141, n146, n148, n151, n155, n156, n157, n158,
         n160, n161, n171, n172, n173, n174, n177, n179, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, DP_OP_116J2_127_7148_n3,
         DP_OP_116J2_127_7148_n4, DP_OP_116J2_127_7148_n5,
         DP_OP_116J2_127_7148_n6, DP_OP_116J2_127_7148_n7,
         DP_OP_116J2_127_7148_n8, DP_OP_113J2_124_6892_n3,
         DP_OP_113J2_124_6892_n4, DP_OP_113J2_124_6892_n5,
         DP_OP_113J2_124_6892_n6, DP_OP_113J2_124_6892_n7,
         DP_OP_113J2_124_6892_n8, C1_Z_6, C1_Z_5, C1_Z_4, C1_Z_3, C1_Z_2,
         C1_Z_1, mult_x_1_n879, mult_x_1_n878, mult_x_1_n877, mult_x_1_n876,
         mult_x_1_n875, mult_x_1_n874, mult_x_1_n873, mult_x_1_n872,
         mult_x_1_n871, mult_x_1_n870, mult_x_1_n869, mult_x_1_n868,
         mult_x_1_n867, mult_x_1_n866, mult_x_1_n865, mult_x_1_n864,
         mult_x_1_n863, mult_x_1_n862, mult_x_1_n861, mult_x_1_n860,
         mult_x_1_n859, mult_x_1_n858, mult_x_1_n857, mult_x_1_n856,
         mult_x_1_n855, mult_x_1_n854, mult_x_1_n852, mult_x_1_n851,
         mult_x_1_n850, mult_x_1_n849, mult_x_1_n848, mult_x_1_n847,
         mult_x_1_n846, mult_x_1_n845, mult_x_1_n844, mult_x_1_n843,
         mult_x_1_n842, mult_x_1_n841, mult_x_1_n840, mult_x_1_n839,
         mult_x_1_n838, mult_x_1_n837, mult_x_1_n836, mult_x_1_n835,
         mult_x_1_n834, mult_x_1_n833, mult_x_1_n832, mult_x_1_n831,
         mult_x_1_n830, mult_x_1_n829, mult_x_1_n828, mult_x_1_n827,
         mult_x_1_n825, mult_x_1_n824, mult_x_1_n823, mult_x_1_n822,
         mult_x_1_n821, mult_x_1_n820, mult_x_1_n819, mult_x_1_n818,
         mult_x_1_n817, mult_x_1_n816, mult_x_1_n815, mult_x_1_n814,
         mult_x_1_n813, mult_x_1_n812, mult_x_1_n811, mult_x_1_n810,
         mult_x_1_n809, mult_x_1_n808, mult_x_1_n807, mult_x_1_n806,
         mult_x_1_n805, mult_x_1_n804, mult_x_1_n803, mult_x_1_n802,
         mult_x_1_n801, mult_x_1_n800, mult_x_1_n798, mult_x_1_n797,
         mult_x_1_n796, mult_x_1_n795, mult_x_1_n794, mult_x_1_n793,
         mult_x_1_n792, mult_x_1_n791, mult_x_1_n790, mult_x_1_n789,
         mult_x_1_n788, mult_x_1_n787, mult_x_1_n786, mult_x_1_n785,
         mult_x_1_n784, mult_x_1_n783, mult_x_1_n782, mult_x_1_n781,
         mult_x_1_n780, mult_x_1_n779, mult_x_1_n778, mult_x_1_n777,
         mult_x_1_n776, mult_x_1_n775, mult_x_1_n774, mult_x_1_n773,
         mult_x_1_n771, mult_x_1_n770, mult_x_1_n769, mult_x_1_n768,
         mult_x_1_n767, mult_x_1_n766, mult_x_1_n765, mult_x_1_n764,
         mult_x_1_n763, mult_x_1_n762, mult_x_1_n761, mult_x_1_n760,
         mult_x_1_n759, mult_x_1_n758, mult_x_1_n757, mult_x_1_n756,
         mult_x_1_n755, mult_x_1_n754, mult_x_1_n753, mult_x_1_n752,
         mult_x_1_n751, mult_x_1_n750, mult_x_1_n749, mult_x_1_n748,
         mult_x_1_n747, mult_x_1_n746, mult_x_1_n744, mult_x_1_n743,
         mult_x_1_n742, mult_x_1_n741, mult_x_1_n740, mult_x_1_n739,
         mult_x_1_n738, mult_x_1_n737, mult_x_1_n736, mult_x_1_n735,
         mult_x_1_n734, mult_x_1_n733, mult_x_1_n732, mult_x_1_n731,
         mult_x_1_n730, mult_x_1_n729, mult_x_1_n728, mult_x_1_n727,
         mult_x_1_n726, mult_x_1_n725, mult_x_1_n724, mult_x_1_n723,
         mult_x_1_n722, mult_x_1_n721, mult_x_1_n720, mult_x_1_n719,
         mult_x_1_n717, mult_x_1_n716, mult_x_1_n715, mult_x_1_n714,
         mult_x_1_n713, mult_x_1_n712, mult_x_1_n711, mult_x_1_n710,
         mult_x_1_n709, mult_x_1_n708, mult_x_1_n707, mult_x_1_n706,
         mult_x_1_n705, mult_x_1_n704, mult_x_1_n703, mult_x_1_n702,
         mult_x_1_n701, mult_x_1_n700, mult_x_1_n699, mult_x_1_n698,
         mult_x_1_n697, mult_x_1_n696, mult_x_1_n695, mult_x_1_n694,
         mult_x_1_n693, mult_x_1_n692, mult_x_1_n690, mult_x_1_n689,
         mult_x_1_n688, mult_x_1_n687, mult_x_1_n686, mult_x_1_n685,
         mult_x_1_n684, mult_x_1_n683, mult_x_1_n682, mult_x_1_n681,
         mult_x_1_n680, mult_x_1_n679, mult_x_1_n678, mult_x_1_n677,
         mult_x_1_n676, mult_x_1_n675, mult_x_1_n674, mult_x_1_n673,
         mult_x_1_n672, mult_x_1_n671, mult_x_1_n670, mult_x_1_n669,
         mult_x_1_n668, mult_x_1_n667, mult_x_1_n666, mult_x_1_n665,
         mult_x_1_n663, mult_x_1_n662, mult_x_1_n661, mult_x_1_n660,
         mult_x_1_n659, mult_x_1_n658, mult_x_1_n657, mult_x_1_n656,
         mult_x_1_n655, mult_x_1_n654, mult_x_1_n653, mult_x_1_n652,
         mult_x_1_n651, mult_x_1_n650, mult_x_1_n649, mult_x_1_n648,
         mult_x_1_n647, mult_x_1_n646, mult_x_1_n645, mult_x_1_n644,
         mult_x_1_n643, mult_x_1_n642, mult_x_1_n641, mult_x_1_n640,
         mult_x_1_n639, mult_x_1_n638, mult_x_1_n637, mult_x_1_n636,
         mult_x_1_n635, mult_x_1_n634, mult_x_1_n633, mult_x_1_n632,
         mult_x_1_n631, mult_x_1_n630, mult_x_1_n629, mult_x_1_n628,
         mult_x_1_n627, mult_x_1_n626, mult_x_1_n625, mult_x_1_n624,
         mult_x_1_n623, mult_x_1_n622, mult_x_1_n621, mult_x_1_n620,
         mult_x_1_n619, mult_x_1_n618, mult_x_1_n617, mult_x_1_n616,
         mult_x_1_n591, mult_x_1_n590, mult_x_1_n589, mult_x_1_n588,
         mult_x_1_n587, mult_x_1_n586, mult_x_1_n583, mult_x_1_n581,
         mult_x_1_n580, mult_x_1_n577, mult_x_1_n575, mult_x_1_n574,
         mult_x_1_n571, mult_x_1_n569, mult_x_1_n567, mult_x_1_n566,
         mult_x_1_n565, mult_x_1_n564, mult_x_1_n563, mult_x_1_n562,
         mult_x_1_n561, mult_x_1_n560, mult_x_1_n559, mult_x_1_n558,
         mult_x_1_n557, mult_x_1_n556, mult_x_1_n555, mult_x_1_n554,
         mult_x_1_n553, mult_x_1_n552, mult_x_1_n551, mult_x_1_n550,
         mult_x_1_n549, mult_x_1_n548, mult_x_1_n547, mult_x_1_n546,
         mult_x_1_n545, mult_x_1_n544, mult_x_1_n543, mult_x_1_n542,
         mult_x_1_n541, mult_x_1_n540, mult_x_1_n539, mult_x_1_n538,
         mult_x_1_n537, mult_x_1_n536, mult_x_1_n535, mult_x_1_n534,
         mult_x_1_n533, mult_x_1_n532, mult_x_1_n531, mult_x_1_n530,
         mult_x_1_n529, mult_x_1_n528, mult_x_1_n527, mult_x_1_n526,
         mult_x_1_n525, mult_x_1_n524, mult_x_1_n523, mult_x_1_n522,
         mult_x_1_n521, mult_x_1_n520, mult_x_1_n519, mult_x_1_n518,
         mult_x_1_n517, mult_x_1_n516, mult_x_1_n515, mult_x_1_n514,
         mult_x_1_n513, mult_x_1_n512, mult_x_1_n511, mult_x_1_n510,
         mult_x_1_n509, mult_x_1_n508, mult_x_1_n507, mult_x_1_n506,
         mult_x_1_n505, mult_x_1_n504, mult_x_1_n503, mult_x_1_n502,
         mult_x_1_n501, mult_x_1_n500, mult_x_1_n499, mult_x_1_n498,
         mult_x_1_n497, mult_x_1_n496, mult_x_1_n495, mult_x_1_n494,
         mult_x_1_n493, mult_x_1_n492, mult_x_1_n491, mult_x_1_n490,
         mult_x_1_n489, mult_x_1_n488, mult_x_1_n487, mult_x_1_n486,
         mult_x_1_n485, mult_x_1_n484, mult_x_1_n483, mult_x_1_n482,
         mult_x_1_n481, mult_x_1_n480, mult_x_1_n479, mult_x_1_n478,
         mult_x_1_n477, mult_x_1_n476, mult_x_1_n475, mult_x_1_n474,
         mult_x_1_n473, mult_x_1_n472, mult_x_1_n471, mult_x_1_n470,
         mult_x_1_n469, mult_x_1_n468, mult_x_1_n467, mult_x_1_n466,
         mult_x_1_n465, mult_x_1_n464, mult_x_1_n463, mult_x_1_n462,
         mult_x_1_n461, mult_x_1_n460, mult_x_1_n459, mult_x_1_n458,
         mult_x_1_n457, mult_x_1_n456, mult_x_1_n455, mult_x_1_n454,
         mult_x_1_n453, mult_x_1_n452, mult_x_1_n451, mult_x_1_n450,
         mult_x_1_n449, mult_x_1_n448, mult_x_1_n447, mult_x_1_n446,
         mult_x_1_n445, mult_x_1_n444, mult_x_1_n443, mult_x_1_n442,
         mult_x_1_n441, mult_x_1_n440, mult_x_1_n439, mult_x_1_n438,
         mult_x_1_n437, mult_x_1_n436, mult_x_1_n435, mult_x_1_n434,
         mult_x_1_n433, mult_x_1_n432, mult_x_1_n431, mult_x_1_n430,
         mult_x_1_n429, mult_x_1_n428, mult_x_1_n427, mult_x_1_n426,
         mult_x_1_n425, mult_x_1_n424, mult_x_1_n423, mult_x_1_n422,
         mult_x_1_n421, mult_x_1_n420, mult_x_1_n419, mult_x_1_n418,
         mult_x_1_n417, mult_x_1_n416, mult_x_1_n415, mult_x_1_n414,
         mult_x_1_n413, mult_x_1_n412, mult_x_1_n411, mult_x_1_n410,
         mult_x_1_n409, mult_x_1_n408, mult_x_1_n407, mult_x_1_n406,
         mult_x_1_n405, mult_x_1_n404, mult_x_1_n403, mult_x_1_n402,
         mult_x_1_n401, mult_x_1_n400, mult_x_1_n399, mult_x_1_n398,
         mult_x_1_n397, mult_x_1_n396, mult_x_1_n395, mult_x_1_n394,
         mult_x_1_n393, mult_x_1_n392, mult_x_1_n391, mult_x_1_n390,
         mult_x_1_n389, mult_x_1_n388, mult_x_1_n387, mult_x_1_n386,
         mult_x_1_n385, mult_x_1_n384, mult_x_1_n383, mult_x_1_n382,
         mult_x_1_n381, mult_x_1_n380, mult_x_1_n379, mult_x_1_n378,
         mult_x_1_n377, mult_x_1_n376, mult_x_1_n375, mult_x_1_n374,
         mult_x_1_n373, mult_x_1_n372, mult_x_1_n371, mult_x_1_n370,
         mult_x_1_n369, mult_x_1_n368, mult_x_1_n367, mult_x_1_n366,
         mult_x_1_n365, mult_x_1_n364, mult_x_1_n363, mult_x_1_n362,
         mult_x_1_n361, mult_x_1_n360, mult_x_1_n359, mult_x_1_n358,
         mult_x_1_n357, mult_x_1_n356, mult_x_1_n355, mult_x_1_n354,
         mult_x_1_n353, mult_x_1_n352, mult_x_1_n351, mult_x_1_n350,
         mult_x_1_n349, mult_x_1_n348, mult_x_1_n347, mult_x_1_n346,
         mult_x_1_n345, mult_x_1_n344, mult_x_1_n343, mult_x_1_n342,
         mult_x_1_n341, mult_x_1_n340, mult_x_1_n339, mult_x_1_n338,
         mult_x_1_n337, mult_x_1_n336, mult_x_1_n335, mult_x_1_n334,
         mult_x_1_n333, mult_x_1_n332, mult_x_1_n331, mult_x_1_n330,
         mult_x_1_n329, mult_x_1_n328, mult_x_1_n327, mult_x_1_n326,
         mult_x_1_n325, mult_x_1_n324, mult_x_1_n323, mult_x_1_n322,
         mult_x_1_n321, mult_x_1_n320, mult_x_1_n319, mult_x_1_n318,
         mult_x_1_n317, mult_x_1_n316, mult_x_1_n315, mult_x_1_n314,
         mult_x_1_n313, mult_x_1_n312, mult_x_1_n311, mult_x_1_n310,
         mult_x_1_n309, mult_x_1_n308, mult_x_1_n307, mult_x_1_n306,
         mult_x_1_n305, mult_x_1_n304, mult_x_1_n303, mult_x_1_n302,
         mult_x_1_n301, mult_x_1_n300, mult_x_1_n299, mult_x_1_n298,
         mult_x_1_n297, mult_x_1_n296, mult_x_1_n295, mult_x_1_n294,
         mult_x_1_n293, mult_x_1_n292, mult_x_1_n291, mult_x_1_n290,
         mult_x_1_n289, mult_x_1_n288, mult_x_1_n287, mult_x_1_n286,
         mult_x_1_n285, mult_x_1_n284, mult_x_1_n283, mult_x_1_n282,
         mult_x_1_n281, mult_x_1_n280, mult_x_1_n279, mult_x_1_n278,
         mult_x_1_n277, mult_x_1_n276, mult_x_1_n275, mult_x_1_n274,
         mult_x_1_n273, mult_x_1_n272, mult_x_1_n271, mult_x_1_n270,
         mult_x_1_n269, mult_x_1_n268, mult_x_1_n267, mult_x_1_n265,
         mult_x_1_n264, mult_x_1_n263, mult_x_1_n262, mult_x_1_n261,
         mult_x_1_n260, mult_x_1_n259, mult_x_1_n258, mult_x_1_n257,
         mult_x_1_n256, mult_x_1_n255, mult_x_1_n254, mult_x_1_n253,
         mult_x_1_n252, mult_x_1_n251, mult_x_1_n250, mult_x_1_n249,
         mult_x_1_n248, mult_x_1_n247, mult_x_1_n246, mult_x_1_n245,
         mult_x_1_n244, mult_x_1_n243, mult_x_1_n242, mult_x_1_n241,
         mult_x_1_n240, mult_x_1_n239, mult_x_1_n238, mult_x_1_n237,
         mult_x_1_n236, mult_x_1_n235, mult_x_1_n234, mult_x_1_n233,
         mult_x_1_n232, mult_x_1_n231, mult_x_1_n230, mult_x_1_n229,
         mult_x_1_n228, mult_x_1_n227, mult_x_1_n226, mult_x_1_n225,
         mult_x_1_n224, mult_x_1_n223, mult_x_1_n222, mult_x_1_n221,
         mult_x_1_n220, mult_x_1_n219, mult_x_1_n218, mult_x_1_n217,
         mult_x_1_n216, mult_x_1_n215, mult_x_1_n214, mult_x_1_n213,
         mult_x_1_n211, mult_x_1_n210, mult_x_1_n209, mult_x_1_n208,
         mult_x_1_n207, mult_x_1_n206, mult_x_1_n205, mult_x_1_n204,
         mult_x_1_n203, mult_x_1_n202, mult_x_1_n201, mult_x_1_n200,
         mult_x_1_n199, mult_x_1_n198, mult_x_1_n197, mult_x_1_n196,
         mult_x_1_n195, mult_x_1_n194, mult_x_1_n193, mult_x_1_n192,
         mult_x_1_n191, mult_x_1_n190, mult_x_1_n189, mult_x_1_n188,
         mult_x_1_n187, mult_x_1_n186, mult_x_1_n185, mult_x_1_n184,
         mult_x_1_n183, mult_x_1_n181, mult_x_1_n180, mult_x_1_n178,
         mult_x_1_n177, mult_x_1_n176, mult_x_1_n175, mult_x_1_n174,
         mult_x_1_n173, mult_x_1_n172, mult_x_1_n171, mult_x_1_n170,
         mult_x_1_n169, mult_x_1_n168, mult_x_1_n167, mult_x_1_n166,
         mult_x_1_n165, mult_x_1_n164, mult_x_1_n163, mult_x_1_n162,
         mult_x_1_n161, mult_x_1_n160, mult_x_1_n159, mult_x_1_n158,
         mult_x_1_n157, mult_x_1_n156, mult_x_1_n155, mult_x_1_n154,
         mult_x_1_n153, mult_x_1_n152, mult_x_1_n151, mult_x_1_n150,
         mult_x_1_n149, mult_x_1_n148, mult_x_1_n147, mult_x_1_n146,
         mult_x_1_n145, mult_x_1_n144, mult_x_1_n143, mult_x_1_n142,
         mult_x_1_n141, mult_x_1_n140, mult_x_1_n139, mult_x_1_n138,
         mult_x_1_n137, mult_x_1_n136, mult_x_1_n135, mult_x_1_n134,
         mult_x_1_n133, mult_x_1_n132, DP_OP_125J2_130_6300_I3,
         DP_OP_125J2_130_6300_I5, DP_OP_125J2_130_6300_n54,
         DP_OP_125J2_130_6300_n43, DP_OP_125J2_130_6300_n42,
         DP_OP_125J2_130_6300_n41, DP_OP_125J2_130_6300_n40,
         DP_OP_125J2_130_6300_n39, DP_OP_125J2_130_6300_n38,
         DP_OP_125J2_130_6300_n37, DP_OP_125J2_130_6300_n36,
         DP_OP_125J2_130_6300_n35, DP_OP_125J2_130_6300_n34,
         DP_OP_125J2_130_6300_n33, DP_OP_125J2_130_6300_n32,
         DP_OP_125J2_130_6300_n31, DP_OP_125J2_130_6300_n30,
         DP_OP_125J2_130_6300_n29, DP_OP_125J2_130_6300_n28,
         DP_OP_125J2_130_6300_n27, DP_OP_125J2_130_6300_n26,
         DP_OP_125J2_130_6300_n25, DP_OP_125J2_130_6300_n20,
         DP_OP_125J2_130_6300_n19, DP_OP_125J2_130_6300_n18,
         DP_OP_125J2_130_6300_n17, DP_OP_125J2_130_6300_n16,
         DP_OP_125J2_130_6300_n15, DP_OP_125J2_130_6300_n14,
         DP_OP_125J2_130_6300_n13, DP_OP_125J2_130_6300_n12,
         DP_OP_125J2_130_6300_n11, DP_OP_125J2_130_6300_n10,
         DP_OP_125J2_130_6300_n9, DP_OP_125J2_130_6300_n8,
         DP_OP_125J2_130_6300_n7, DP_OP_125J2_130_6300_n6,
         DP_OP_125J2_130_6300_n5, DP_OP_125J2_130_6300_n4,
         DP_OP_125J2_130_6300_n3, DP_OP_125J2_130_6300_n2,
         DP_OP_125J2_130_6300_n1, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [23:0] a_m;
  wire   [9:0] b_e;
  wire   [23:0] b_m;
  wire   [49:2] product;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ao211d1_hd U246 ( .A(n20), .B(n155), .C(i_RST), .D(n1167), .Y(n350) );
  oa22d1_hd U247 ( .A(n156), .B(n157), .C(n1221), .D(n158), .Y(n351) );
  oa22d1_hd U249 ( .A(n160), .B(n157), .C(n462), .D(n158), .Y(n352) );
  oa22d1_hd U250 ( .A(n161), .B(n157), .C(n34), .D(n158), .Y(n353) );
  oa22d1_hd U267 ( .A(n171), .B(n157), .C(n1220), .D(n158), .Y(n357) );
  nd4d1_hd U269 ( .A(n160), .B(n172), .C(n173), .D(n174), .Y(n158) );
  ao211d1_hd U270 ( .A(n29), .B(n36), .C(i_RST), .D(n1167), .Y(n174) );
  ao211d1_hd U281 ( .A(n1165), .B(n177), .C(i_RST), .D(n179), .Y(n358) );
  ivd1_hd U364 ( .A(i_RST), .Y(N34) );
  fad1_hd DP_OP_116J2_127_7148_U6 ( .A(n478), .B(n1213), .CI(
        DP_OP_116J2_127_7148_n4), .CO(DP_OP_116J2_127_7148_n3), .S(C82_DATA2_6) );
  fad1_hd DP_OP_116J2_127_7148_U7 ( .A(n480), .B(n1212), .CI(
        DP_OP_116J2_127_7148_n5), .CO(DP_OP_116J2_127_7148_n4), .S(C82_DATA2_5) );
  fad1_hd DP_OP_116J2_127_7148_U8 ( .A(n480), .B(n1211), .CI(
        DP_OP_116J2_127_7148_n6), .CO(DP_OP_116J2_127_7148_n5), .S(C82_DATA2_4) );
  fad1_hd DP_OP_116J2_127_7148_U9 ( .A(n478), .B(n1210), .CI(
        DP_OP_116J2_127_7148_n7), .CO(DP_OP_116J2_127_7148_n6), .S(C82_DATA2_3) );
  fad1_hd DP_OP_116J2_127_7148_U10 ( .A(n480), .B(n1209), .CI(
        DP_OP_116J2_127_7148_n8), .CO(DP_OP_116J2_127_7148_n7), .S(C82_DATA2_2) );
  fad1_hd DP_OP_116J2_127_7148_U11 ( .A(n478), .B(n1208), .CI(n1207), .CO(
        DP_OP_116J2_127_7148_n8), .S(C82_DATA2_1) );
  fad1_hd DP_OP_113J2_124_6892_U6 ( .A(n481), .B(C1_Z_6), .CI(
        DP_OP_113J2_124_6892_n4), .CO(DP_OP_113J2_124_6892_n3), .S(C81_DATA2_6) );
  fad1_hd DP_OP_113J2_124_6892_U7 ( .A(n479), .B(C1_Z_5), .CI(
        DP_OP_113J2_124_6892_n5), .CO(DP_OP_113J2_124_6892_n4), .S(C81_DATA2_5) );
  fad1_hd DP_OP_113J2_124_6892_U8 ( .A(n479), .B(C1_Z_4), .CI(
        DP_OP_113J2_124_6892_n6), .CO(DP_OP_113J2_124_6892_n5), .S(C81_DATA2_4) );
  fad1_hd DP_OP_113J2_124_6892_U9 ( .A(n481), .B(C1_Z_3), .CI(
        DP_OP_113J2_124_6892_n7), .CO(DP_OP_113J2_124_6892_n6), .S(C81_DATA2_3) );
  fad1_hd DP_OP_113J2_124_6892_U10 ( .A(n479), .B(C1_Z_2), .CI(
        DP_OP_113J2_124_6892_n8), .CO(DP_OP_113J2_124_6892_n7), .S(C81_DATA2_2) );
  fad1_hd DP_OP_113J2_124_6892_U11 ( .A(n481), .B(C1_Z_1), .CI(n1206), .CO(
        DP_OP_113J2_124_6892_n8), .S(C81_DATA2_1) );
  had1_hd mult_x_1_U362 ( .A(n917), .B(mult_x_1_n771), .CO(mult_x_1_n530), .S(
        mult_x_1_n531) );
  fad1_hd mult_x_1_U361 ( .A(mult_x_1_n795), .B(mult_x_1_n531), .CI(
        mult_x_1_n536), .CO(mult_x_1_n528), .S(mult_x_1_n529) );
  fad1_hd mult_x_1_U357 ( .A(mult_x_1_n794), .B(mult_x_1_n523), .CI(
        mult_x_1_n528), .CO(mult_x_1_n520), .S(mult_x_1_n521) );
  fad1_hd mult_x_1_U353 ( .A(mult_x_1_n793), .B(mult_x_1_n515), .CI(
        mult_x_1_n520), .CO(mult_x_1_n512), .S(mult_x_1_n513) );
  had1_hd mult_x_1_U350 ( .A(n910), .B(mult_x_1_n744), .CO(mult_x_1_n506), .S(
        mult_x_1_n507) );
  fad1_hd mult_x_1_U349 ( .A(mult_x_1_n768), .B(mult_x_1_n507), .CI(
        mult_x_1_n514), .CO(mult_x_1_n504), .S(mult_x_1_n505) );
  fad1_hd mult_x_1_U348 ( .A(mult_x_1_n792), .B(mult_x_1_n505), .CI(
        mult_x_1_n512), .CO(mult_x_1_n502), .S(mult_x_1_n503) );
  had1_hd mult_x_1_U345 ( .A(mult_x_1_n743), .B(mult_x_1_n506), .CO(
        mult_x_1_n496), .S(mult_x_1_n497) );
  fad1_hd mult_x_1_U344 ( .A(mult_x_1_n767), .B(mult_x_1_n497), .CI(
        mult_x_1_n504), .CO(mult_x_1_n494), .S(mult_x_1_n495) );
  fad1_hd mult_x_1_U343 ( .A(mult_x_1_n791), .B(mult_x_1_n495), .CI(
        mult_x_1_n502), .CO(mult_x_1_n492), .S(mult_x_1_n493) );
  had1_hd mult_x_1_U340 ( .A(mult_x_1_n742), .B(mult_x_1_n496), .CO(
        mult_x_1_n486), .S(mult_x_1_n487) );
  fad1_hd mult_x_1_U339 ( .A(mult_x_1_n766), .B(mult_x_1_n487), .CI(
        mult_x_1_n494), .CO(mult_x_1_n484), .S(mult_x_1_n485) );
  fad1_hd mult_x_1_U338 ( .A(mult_x_1_n790), .B(mult_x_1_n485), .CI(
        mult_x_1_n492), .CO(mult_x_1_n482), .S(mult_x_1_n483) );
  had1_hd mult_x_1_U335 ( .A(n903), .B(mult_x_1_n717), .CO(mult_x_1_n476), .S(
        mult_x_1_n477) );
  fad1_hd mult_x_1_U334 ( .A(mult_x_1_n741), .B(mult_x_1_n477), .CI(
        mult_x_1_n486), .CO(mult_x_1_n474), .S(mult_x_1_n475) );
  fad1_hd mult_x_1_U333 ( .A(mult_x_1_n765), .B(mult_x_1_n475), .CI(
        mult_x_1_n484), .CO(mult_x_1_n472), .S(mult_x_1_n473) );
  fad1_hd mult_x_1_U332 ( .A(mult_x_1_n789), .B(mult_x_1_n473), .CI(
        mult_x_1_n482), .CO(mult_x_1_n470), .S(mult_x_1_n471) );
  had1_hd mult_x_1_U329 ( .A(mult_x_1_n716), .B(mult_x_1_n476), .CO(
        mult_x_1_n464), .S(mult_x_1_n465) );
  fad1_hd mult_x_1_U328 ( .A(mult_x_1_n740), .B(mult_x_1_n465), .CI(
        mult_x_1_n474), .CO(mult_x_1_n462), .S(mult_x_1_n463) );
  fad1_hd mult_x_1_U327 ( .A(mult_x_1_n764), .B(mult_x_1_n463), .CI(
        mult_x_1_n472), .CO(mult_x_1_n460), .S(mult_x_1_n461) );
  fad1_hd mult_x_1_U326 ( .A(mult_x_1_n788), .B(mult_x_1_n461), .CI(
        mult_x_1_n470), .CO(mult_x_1_n458), .S(mult_x_1_n459) );
  had1_hd mult_x_1_U323 ( .A(mult_x_1_n715), .B(mult_x_1_n464), .CO(
        mult_x_1_n452), .S(mult_x_1_n453) );
  fad1_hd mult_x_1_U322 ( .A(mult_x_1_n739), .B(mult_x_1_n453), .CI(
        mult_x_1_n462), .CO(mult_x_1_n450), .S(mult_x_1_n451) );
  fad1_hd mult_x_1_U321 ( .A(mult_x_1_n763), .B(mult_x_1_n451), .CI(
        mult_x_1_n460), .CO(mult_x_1_n448), .S(mult_x_1_n449) );
  fad1_hd mult_x_1_U320 ( .A(mult_x_1_n787), .B(mult_x_1_n449), .CI(
        mult_x_1_n458), .CO(mult_x_1_n446), .S(mult_x_1_n447) );
  had1_hd mult_x_1_U317 ( .A(n896), .B(mult_x_1_n690), .CO(mult_x_1_n440), .S(
        mult_x_1_n441) );
  fad1_hd mult_x_1_U316 ( .A(mult_x_1_n714), .B(mult_x_1_n441), .CI(
        mult_x_1_n452), .CO(mult_x_1_n438), .S(mult_x_1_n439) );
  fad1_hd mult_x_1_U315 ( .A(mult_x_1_n738), .B(mult_x_1_n439), .CI(
        mult_x_1_n450), .CO(mult_x_1_n436), .S(mult_x_1_n437) );
  fad1_hd mult_x_1_U314 ( .A(mult_x_1_n762), .B(mult_x_1_n437), .CI(
        mult_x_1_n448), .CO(mult_x_1_n434), .S(mult_x_1_n435) );
  fad1_hd mult_x_1_U313 ( .A(mult_x_1_n786), .B(mult_x_1_n435), .CI(
        mult_x_1_n446), .CO(mult_x_1_n432), .S(mult_x_1_n433) );
  had1_hd mult_x_1_U310 ( .A(mult_x_1_n689), .B(mult_x_1_n440), .CO(
        mult_x_1_n426), .S(mult_x_1_n427) );
  fad1_hd mult_x_1_U309 ( .A(mult_x_1_n713), .B(mult_x_1_n427), .CI(
        mult_x_1_n438), .CO(mult_x_1_n424), .S(mult_x_1_n425) );
  fad1_hd mult_x_1_U308 ( .A(mult_x_1_n737), .B(mult_x_1_n425), .CI(
        mult_x_1_n436), .CO(mult_x_1_n422), .S(mult_x_1_n423) );
  fad1_hd mult_x_1_U307 ( .A(mult_x_1_n761), .B(mult_x_1_n423), .CI(
        mult_x_1_n434), .CO(mult_x_1_n420), .S(mult_x_1_n421) );
  fad1_hd mult_x_1_U306 ( .A(mult_x_1_n785), .B(mult_x_1_n421), .CI(
        mult_x_1_n432), .CO(mult_x_1_n418), .S(mult_x_1_n419) );
  had1_hd mult_x_1_U303 ( .A(mult_x_1_n688), .B(mult_x_1_n426), .CO(
        mult_x_1_n412), .S(mult_x_1_n413) );
  fad1_hd mult_x_1_U302 ( .A(mult_x_1_n712), .B(mult_x_1_n413), .CI(
        mult_x_1_n424), .CO(mult_x_1_n410), .S(mult_x_1_n411) );
  fad1_hd mult_x_1_U301 ( .A(mult_x_1_n736), .B(mult_x_1_n411), .CI(
        mult_x_1_n422), .CO(mult_x_1_n408), .S(mult_x_1_n409) );
  fad1_hd mult_x_1_U300 ( .A(mult_x_1_n760), .B(mult_x_1_n409), .CI(
        mult_x_1_n420), .CO(mult_x_1_n406), .S(mult_x_1_n407) );
  fad1_hd mult_x_1_U299 ( .A(mult_x_1_n784), .B(mult_x_1_n407), .CI(
        mult_x_1_n418), .CO(mult_x_1_n404), .S(mult_x_1_n405) );
  fad1_hd mult_x_1_U296 ( .A(mult_x_1_n687), .B(mult_x_1_n591), .CI(
        mult_x_1_n412), .CO(mult_x_1_n398), .S(mult_x_1_n399) );
  fad1_hd mult_x_1_U295 ( .A(mult_x_1_n711), .B(mult_x_1_n399), .CI(
        mult_x_1_n410), .CO(mult_x_1_n396), .S(mult_x_1_n397) );
  fad1_hd mult_x_1_U294 ( .A(mult_x_1_n735), .B(mult_x_1_n397), .CI(
        mult_x_1_n408), .CO(mult_x_1_n394), .S(mult_x_1_n395) );
  fad1_hd mult_x_1_U293 ( .A(mult_x_1_n759), .B(mult_x_1_n395), .CI(
        mult_x_1_n406), .CO(mult_x_1_n392), .S(mult_x_1_n393) );
  fad1_hd mult_x_1_U292 ( .A(mult_x_1_n783), .B(mult_x_1_n393), .CI(
        mult_x_1_n404), .CO(mult_x_1_n390), .S(mult_x_1_n391) );
  fad1_hd mult_x_1_U289 ( .A(mult_x_1_n686), .B(mult_x_1_n590), .CI(
        mult_x_1_n398), .CO(mult_x_1_n384), .S(mult_x_1_n385) );
  fad1_hd mult_x_1_U288 ( .A(mult_x_1_n710), .B(mult_x_1_n385), .CI(
        mult_x_1_n396), .CO(mult_x_1_n382), .S(mult_x_1_n383) );
  fad1_hd mult_x_1_U287 ( .A(mult_x_1_n734), .B(mult_x_1_n383), .CI(
        mult_x_1_n394), .CO(mult_x_1_n380), .S(mult_x_1_n381) );
  fad1_hd mult_x_1_U286 ( .A(mult_x_1_n758), .B(mult_x_1_n381), .CI(
        mult_x_1_n392), .CO(mult_x_1_n378), .S(mult_x_1_n379) );
  fad1_hd mult_x_1_U282 ( .A(mult_x_1_n589), .B(n945), .CI(mult_x_1_n685), 
        .CO(mult_x_1_n370), .S(mult_x_1_n371) );
  fad1_hd mult_x_1_U281 ( .A(mult_x_1_n371), .B(mult_x_1_n384), .CI(
        mult_x_1_n709), .CO(mult_x_1_n368), .S(mult_x_1_n369) );
  fad1_hd mult_x_1_U280 ( .A(mult_x_1_n369), .B(mult_x_1_n382), .CI(
        mult_x_1_n733), .CO(mult_x_1_n366), .S(mult_x_1_n367) );
  fad1_hd mult_x_1_U279 ( .A(mult_x_1_n367), .B(mult_x_1_n380), .CI(
        mult_x_1_n757), .CO(mult_x_1_n364), .S(mult_x_1_n365) );
  fad1_hd mult_x_1_U278 ( .A(mult_x_1_n365), .B(mult_x_1_n378), .CI(
        mult_x_1_n781), .CO(mult_x_1_n362), .S(mult_x_1_n363) );
  fad1_hd mult_x_1_U275 ( .A(mult_x_1_n588), .B(n945), .CI(mult_x_1_n684), 
        .CO(mult_x_1_n356), .S(mult_x_1_n357) );
  fad1_hd mult_x_1_U274 ( .A(mult_x_1_n357), .B(mult_x_1_n370), .CI(
        mult_x_1_n708), .CO(mult_x_1_n354), .S(mult_x_1_n355) );
  fad1_hd mult_x_1_U273 ( .A(mult_x_1_n355), .B(mult_x_1_n368), .CI(
        mult_x_1_n366), .CO(mult_x_1_n352), .S(mult_x_1_n353) );
  fad1_hd mult_x_1_U272 ( .A(mult_x_1_n353), .B(mult_x_1_n732), .CI(
        mult_x_1_n364), .CO(mult_x_1_n350), .S(mult_x_1_n351) );
  fad1_hd mult_x_1_U268 ( .A(mult_x_1_n587), .B(n945), .CI(mult_x_1_n683), 
        .CO(mult_x_1_n342), .S(mult_x_1_n343) );
  fad1_hd mult_x_1_U267 ( .A(mult_x_1_n343), .B(mult_x_1_n356), .CI(
        mult_x_1_n354), .CO(mult_x_1_n340), .S(mult_x_1_n341) );
  fad1_hd mult_x_1_U266 ( .A(mult_x_1_n341), .B(mult_x_1_n707), .CI(
        mult_x_1_n352), .CO(mult_x_1_n338), .S(mult_x_1_n339) );
  fad1_hd mult_x_1_U265 ( .A(mult_x_1_n339), .B(mult_x_1_n731), .CI(
        mult_x_1_n350), .CO(mult_x_1_n336), .S(mult_x_1_n337) );
  fad1_hd mult_x_1_U261 ( .A(n933), .B(n940), .CI(mult_x_1_n586), .CO(
        mult_x_1_n328), .S(mult_x_1_n329) );
  fad1_hd mult_x_1_U260 ( .A(mult_x_1_n342), .B(mult_x_1_n329), .CI(
        mult_x_1_n682), .CO(mult_x_1_n326), .S(mult_x_1_n327) );
  fad1_hd mult_x_1_U259 ( .A(mult_x_1_n706), .B(mult_x_1_n327), .CI(
        mult_x_1_n340), .CO(mult_x_1_n324), .S(mult_x_1_n325) );
  fad1_hd mult_x_1_U258 ( .A(mult_x_1_n338), .B(mult_x_1_n325), .CI(
        mult_x_1_n730), .CO(mult_x_1_n322), .S(mult_x_1_n323) );
  fad1_hd mult_x_1_U253 ( .A(mult_x_1_n328), .B(mult_x_1_n315), .CI(
        mult_x_1_n681), .CO(mult_x_1_n313), .S(mult_x_1_n314) );
  fad1_hd mult_x_1_U252 ( .A(mult_x_1_n314), .B(mult_x_1_n326), .CI(
        mult_x_1_n705), .CO(mult_x_1_n311), .S(mult_x_1_n312) );
  fad1_hd mult_x_1_U251 ( .A(mult_x_1_n312), .B(mult_x_1_n324), .CI(
        mult_x_1_n729), .CO(mult_x_1_n309), .S(mult_x_1_n310) );
  fad1_hd mult_x_1_U246 ( .A(mult_x_1_n302), .B(n878), .CI(mult_x_1_n313), 
        .CO(mult_x_1_n300), .S(mult_x_1_n301) );
  fad1_hd mult_x_1_U245 ( .A(mult_x_1_n301), .B(mult_x_1_n680), .CI(
        mult_x_1_n704), .CO(mult_x_1_n298), .S(mult_x_1_n299) );
  fad1_hd mult_x_1_U244 ( .A(mult_x_1_n299), .B(mult_x_1_n311), .CI(
        mult_x_1_n309), .CO(mult_x_1_n296), .S(mult_x_1_n297) );
  fad1_hd mult_x_1_U240 ( .A(n879), .B(n925), .CI(mult_x_1_n583), .CO(
        mult_x_1_n288), .S(mult_x_1_n289) );
  fad1_hd mult_x_1_U239 ( .A(mult_x_1_n679), .B(mult_x_1_n289), .CI(
        mult_x_1_n300), .CO(mult_x_1_n286), .S(mult_x_1_n287) );
  fad1_hd mult_x_1_U238 ( .A(mult_x_1_n298), .B(mult_x_1_n287), .CI(
        mult_x_1_n703), .CO(mult_x_1_n284), .S(mult_x_1_n285) );
  fad1_hd mult_x_1_U233 ( .A(mult_x_1_n288), .B(mult_x_1_n277), .CI(
        mult_x_1_n678), .CO(mult_x_1_n275), .S(mult_x_1_n276) );
  fad1_hd mult_x_1_U232 ( .A(mult_x_1_n276), .B(mult_x_1_n286), .CI(
        mult_x_1_n702), .CO(mult_x_1_n273), .S(mult_x_1_n274) );
  fad1_hd mult_x_1_U227 ( .A(mult_x_1_n277), .B(mult_x_1_n581), .CI(
        mult_x_1_n677), .CO(mult_x_1_n264), .S(mult_x_1_n265) );
  fad1_hd mult_x_1_U226 ( .A(mult_x_1_n265), .B(mult_x_1_n275), .CI(
        mult_x_1_n273), .CO(mult_x_1_n262), .S(mult_x_1_n263) );
  fad1_hd mult_x_1_U222 ( .A(mult_x_1_n580), .B(n919), .CI(n880), .CO(
        mult_x_1_n254), .S(mult_x_1_n255) );
  fad1_hd mult_x_1_U221 ( .A(mult_x_1_n264), .B(mult_x_1_n255), .CI(
        mult_x_1_n676), .CO(mult_x_1_n252), .S(mult_x_1_n253) );
  fad1_hd mult_x_1_U216 ( .A(mult_x_1_n254), .B(mult_x_1_n245), .CI(
        mult_x_1_n675), .CO(mult_x_1_n243), .S(mult_x_1_n244) );
  fad1_hd mult_x_1_U211 ( .A(mult_x_1_n236), .B(n881), .CI(mult_x_1_n243), 
        .CO(mult_x_1_n234), .S(mult_x_1_n235) );
  fad1_hd mult_x_1_U207 ( .A(n882), .B(n912), .CI(mult_x_1_n577), .CO(
        mult_x_1_n226), .S(mult_x_1_n227) );
  fad1_hd mult_x_1_U202 ( .A(mult_x_1_n226), .B(mult_x_1_n219), .CI(
        mult_x_1_n672), .CO(mult_x_1_n217), .S(mult_x_1_n218) );
  fad1_hd mult_x_1_U198 ( .A(mult_x_1_n219), .B(mult_x_1_n575), .CI(
        mult_x_1_n671), .CO(mult_x_1_n210), .S(mult_x_1_n211) );
  fad1_hd mult_x_1_U195 ( .A(mult_x_1_n574), .B(n905), .CI(n883), .CO(
        mult_x_1_n204), .S(mult_x_1_n205) );
  had1_hd DP_OP_125J2_130_6300_U32 ( .A(b_e[0]), .B(a_e[0]), .CO(
        DP_OP_125J2_130_6300_n20), .S(DP_OP_125J2_130_6300_n34) );
  fad1_hd DP_OP_125J2_130_6300_U31 ( .A(a_e[1]), .B(b_e[1]), .CI(
        DP_OP_125J2_130_6300_n20), .CO(DP_OP_125J2_130_6300_n19), .S(
        DP_OP_125J2_130_6300_n35) );
  fad1_hd DP_OP_125J2_130_6300_U30 ( .A(a_e[2]), .B(b_e[2]), .CI(
        DP_OP_125J2_130_6300_n19), .CO(DP_OP_125J2_130_6300_n18), .S(
        DP_OP_125J2_130_6300_n36) );
  fad1_hd DP_OP_125J2_130_6300_U29 ( .A(a_e[3]), .B(b_e[3]), .CI(
        DP_OP_125J2_130_6300_n18), .CO(DP_OP_125J2_130_6300_n17), .S(
        DP_OP_125J2_130_6300_n37) );
  fad1_hd DP_OP_125J2_130_6300_U28 ( .A(a_e[4]), .B(b_e[4]), .CI(
        DP_OP_125J2_130_6300_n17), .CO(DP_OP_125J2_130_6300_n16), .S(
        DP_OP_125J2_130_6300_n38) );
  fad1_hd DP_OP_125J2_130_6300_U27 ( .A(a_e[5]), .B(b_e[5]), .CI(
        DP_OP_125J2_130_6300_n16), .CO(DP_OP_125J2_130_6300_n15), .S(
        DP_OP_125J2_130_6300_n39) );
  fad1_hd DP_OP_125J2_130_6300_U26 ( .A(a_e[6]), .B(b_e[6]), .CI(
        DP_OP_125J2_130_6300_n15), .CO(DP_OP_125J2_130_6300_n14), .S(
        DP_OP_125J2_130_6300_n40) );
  fad1_hd DP_OP_125J2_130_6300_U25 ( .A(a_e[7]), .B(b_e[7]), .CI(
        DP_OP_125J2_130_6300_n14), .CO(DP_OP_125J2_130_6300_n13), .S(
        DP_OP_125J2_130_6300_n41) );
  fad1_hd DP_OP_125J2_130_6300_U24 ( .A(a_e[8]), .B(b_e[8]), .CI(
        DP_OP_125J2_130_6300_n13), .CO(DP_OP_125J2_130_6300_n12), .S(
        DP_OP_125J2_130_6300_n42) );
  ivd1_hd DP_OP_125J2_130_6300_U11 ( .A(DP_OP_125J2_130_6300_n10), .Y(N466) );
  fad1_hd DP_OP_125J2_130_6300_U10 ( .A(DP_OP_125J2_130_6300_n10), .B(n573), 
        .CI(DP_OP_125J2_130_6300_n25), .CO(DP_OP_125J2_130_6300_n9), .S(N467)
         );
  fad1_hd DP_OP_125J2_130_6300_U9 ( .A(DP_OP_125J2_130_6300_n26), .B(n571), 
        .CI(DP_OP_125J2_130_6300_n9), .CO(DP_OP_125J2_130_6300_n8), .S(N468)
         );
  fad1_hd DP_OP_125J2_130_6300_U8 ( .A(DP_OP_125J2_130_6300_n27), .B(n572), 
        .CI(DP_OP_125J2_130_6300_n8), .CO(DP_OP_125J2_130_6300_n7), .S(N469)
         );
  fad1_hd DP_OP_125J2_130_6300_U7 ( .A(DP_OP_125J2_130_6300_n28), .B(n573), 
        .CI(DP_OP_125J2_130_6300_n7), .CO(DP_OP_125J2_130_6300_n6), .S(N470)
         );
  fad1_hd DP_OP_125J2_130_6300_U6 ( .A(DP_OP_125J2_130_6300_n29), .B(n572), 
        .CI(DP_OP_125J2_130_6300_n6), .CO(DP_OP_125J2_130_6300_n5), .S(N471)
         );
  fad1_hd DP_OP_125J2_130_6300_U5 ( .A(DP_OP_125J2_130_6300_n30), .B(n573), 
        .CI(DP_OP_125J2_130_6300_n5), .CO(DP_OP_125J2_130_6300_n4), .S(N472)
         );
  fad1_hd DP_OP_125J2_130_6300_U4 ( .A(DP_OP_125J2_130_6300_n31), .B(n571), 
        .CI(DP_OP_125J2_130_6300_n4), .CO(DP_OP_125J2_130_6300_n3), .S(N473)
         );
  fad1_hd DP_OP_125J2_130_6300_U3 ( .A(DP_OP_125J2_130_6300_n32), .B(n573), 
        .CI(DP_OP_125J2_130_6300_n3), .CO(DP_OP_125J2_130_6300_n2), .S(N474)
         );
  fds2d1_hd a_e_reg_7_ ( .CRN(n141), .D(n138), .CK(i_CLK), .Q(n10), .QN(a_e[7]) );
  fds2d1_hd b_e_reg_7_ ( .CRN(n151), .D(n148), .CK(i_CLK), .Q(n14), .QN(b_e[7]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n319), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n356), .CK(i_CLK), .Q(b_e[9]) );
  fad1_hd mult_x_1_U215 ( .A(mult_x_1_n244), .B(mult_x_1_n252), .CI(
        mult_x_1_n699), .CO(mult_x_1_n241), .S(mult_x_1_n242) );
  fad1_hd mult_x_1_U231 ( .A(mult_x_1_n274), .B(mult_x_1_n284), .CI(
        mult_x_1_n726), .CO(mult_x_1_n271), .S(mult_x_1_n272) );
  fad1_hd mult_x_1_U250 ( .A(mult_x_1_n310), .B(mult_x_1_n322), .CI(
        mult_x_1_n753), .CO(mult_x_1_n307), .S(mult_x_1_n308) );
  fad1_hd mult_x_1_U271 ( .A(mult_x_1_n351), .B(mult_x_1_n756), .CI(
        mult_x_1_n780), .CO(mult_x_1_n348), .S(mult_x_1_n349) );
  fad1_hd mult_x_1_U186 ( .A(mult_x_1_n571), .B(n898), .CI(n885), .CO(
        mult_x_1_n188), .S(mult_x_1_n189) );
  fad1_hd mult_x_1_U206 ( .A(mult_x_1_n673), .B(mult_x_1_n227), .CI(
        mult_x_1_n234), .CO(mult_x_1_n224), .S(mult_x_1_n225) );
  fad1_hd mult_x_1_U210 ( .A(mult_x_1_n235), .B(mult_x_1_n674), .CI(
        mult_x_1_n698), .CO(mult_x_1_n232), .S(mult_x_1_n233) );
  fad1_hd mult_x_1_U220 ( .A(mult_x_1_n700), .B(mult_x_1_n253), .CI(
        mult_x_1_n262), .CO(mult_x_1_n250), .S(mult_x_1_n251) );
  fad1_hd mult_x_1_U225 ( .A(mult_x_1_n263), .B(mult_x_1_n701), .CI(
        mult_x_1_n725), .CO(mult_x_1_n260), .S(mult_x_1_n261) );
  fad1_hd mult_x_1_U237 ( .A(mult_x_1_n727), .B(mult_x_1_n285), .CI(
        mult_x_1_n296), .CO(mult_x_1_n282), .S(mult_x_1_n283) );
  fad1_hd mult_x_1_U243 ( .A(mult_x_1_n297), .B(mult_x_1_n728), .CI(
        mult_x_1_n752), .CO(mult_x_1_n294), .S(mult_x_1_n295) );
  fad1_hd mult_x_1_U257 ( .A(mult_x_1_n754), .B(mult_x_1_n323), .CI(
        mult_x_1_n336), .CO(mult_x_1_n320), .S(mult_x_1_n321) );
  fad1_hd mult_x_1_U264 ( .A(mult_x_1_n337), .B(mult_x_1_n755), .CI(
        mult_x_1_n779), .CO(mult_x_1_n334), .S(mult_x_1_n335) );
  had1_hd mult_x_1_U358 ( .A(mult_x_1_n770), .B(mult_x_1_n530), .CO(
        mult_x_1_n522), .S(mult_x_1_n523) );
  had1_hd mult_x_1_U354 ( .A(mult_x_1_n769), .B(mult_x_1_n522), .CO(
        mult_x_1_n514), .S(mult_x_1_n515) );
  had1_hd mult_x_1_U371 ( .A(n924), .B(mult_x_1_n798), .CO(mult_x_1_n548), .S(
        mult_x_1_n549) );
  had1_hd mult_x_1_U368 ( .A(mult_x_1_n797), .B(mult_x_1_n548), .CO(
        mult_x_1_n542), .S(mult_x_1_n543) );
  had1_hd mult_x_1_U365 ( .A(mult_x_1_n796), .B(mult_x_1_n542), .CO(
        mult_x_1_n536), .S(mult_x_1_n537) );
  fad1_hd mult_x_1_U285 ( .A(mult_x_1_n782), .B(mult_x_1_n379), .CI(
        mult_x_1_n390), .CO(mult_x_1_n376), .S(mult_x_1_n377) );
  had1_hd mult_x_1_U377 ( .A(n931), .B(mult_x_1_n825), .CO(mult_x_1_n560), .S(
        mult_x_1_n561) );
  fad1_hd mult_x_1_U370 ( .A(mult_x_1_n822), .B(mult_x_1_n549), .CI(
        mult_x_1_n552), .CO(mult_x_1_n546), .S(mult_x_1_n547) );
  fad1_hd mult_x_1_U367 ( .A(mult_x_1_n821), .B(mult_x_1_n543), .CI(
        mult_x_1_n546), .CO(mult_x_1_n540), .S(mult_x_1_n541) );
  fad1_hd mult_x_1_U364 ( .A(mult_x_1_n820), .B(mult_x_1_n537), .CI(
        mult_x_1_n540), .CO(mult_x_1_n534), .S(mult_x_1_n535) );
  fad1_hd mult_x_1_U360 ( .A(mult_x_1_n819), .B(mult_x_1_n529), .CI(
        mult_x_1_n534), .CO(mult_x_1_n526), .S(mult_x_1_n527) );
  fad1_hd mult_x_1_U356 ( .A(mult_x_1_n818), .B(mult_x_1_n521), .CI(
        mult_x_1_n526), .CO(mult_x_1_n518), .S(mult_x_1_n519) );
  fad1_hd mult_x_1_U352 ( .A(mult_x_1_n817), .B(mult_x_1_n513), .CI(
        mult_x_1_n518), .CO(mult_x_1_n510), .S(mult_x_1_n511) );
  fad1_hd mult_x_1_U347 ( .A(mult_x_1_n816), .B(mult_x_1_n503), .CI(
        mult_x_1_n510), .CO(mult_x_1_n500), .S(mult_x_1_n501) );
  fad1_hd mult_x_1_U342 ( .A(mult_x_1_n815), .B(mult_x_1_n493), .CI(
        mult_x_1_n500), .CO(mult_x_1_n490), .S(mult_x_1_n491) );
  fad1_hd mult_x_1_U337 ( .A(mult_x_1_n814), .B(mult_x_1_n483), .CI(
        mult_x_1_n490), .CO(mult_x_1_n480), .S(mult_x_1_n481) );
  fad1_hd mult_x_1_U331 ( .A(mult_x_1_n813), .B(mult_x_1_n471), .CI(
        mult_x_1_n480), .CO(mult_x_1_n468), .S(mult_x_1_n469) );
  fad1_hd mult_x_1_U325 ( .A(mult_x_1_n812), .B(mult_x_1_n459), .CI(
        mult_x_1_n468), .CO(mult_x_1_n456), .S(mult_x_1_n457) );
  fad1_hd mult_x_1_U319 ( .A(mult_x_1_n811), .B(mult_x_1_n447), .CI(
        mult_x_1_n456), .CO(mult_x_1_n444), .S(mult_x_1_n445) );
  fad1_hd mult_x_1_U312 ( .A(mult_x_1_n810), .B(mult_x_1_n433), .CI(
        mult_x_1_n444), .CO(mult_x_1_n430), .S(mult_x_1_n431) );
  fad1_hd mult_x_1_U305 ( .A(mult_x_1_n809), .B(mult_x_1_n419), .CI(
        mult_x_1_n430), .CO(mult_x_1_n416), .S(mult_x_1_n417) );
  fad1_hd mult_x_1_U298 ( .A(mult_x_1_n808), .B(mult_x_1_n405), .CI(
        mult_x_1_n416), .CO(mult_x_1_n402), .S(mult_x_1_n403) );
  fad1_hd mult_x_1_U291 ( .A(mult_x_1_n807), .B(mult_x_1_n391), .CI(
        mult_x_1_n402), .CO(mult_x_1_n388), .S(mult_x_1_n389) );
  had1_hd mult_x_1_U380 ( .A(n938), .B(mult_x_1_n852), .CO(mult_x_1_n566), .S(
        mult_x_1_n567) );
  fad1_hd mult_x_1_U376 ( .A(mult_x_1_n849), .B(mult_x_1_n561), .CI(
        mult_x_1_n562), .CO(mult_x_1_n558), .S(mult_x_1_n559) );
  had1_hd mult_x_1_U179 ( .A(n945), .B(mult_x_1_n879), .CO(mult_x_1_n178), .S(
        N176) );
  fad1_hd mult_x_1_U176 ( .A(mult_x_1_n876), .B(mult_x_1_n567), .CI(
        mult_x_1_n176), .CO(mult_x_1_n175), .S(N179) );
  fad1_hd mult_x_1_U175 ( .A(mult_x_1_n875), .B(mult_x_1_n565), .CI(
        mult_x_1_n175), .CO(mult_x_1_n174), .S(N180) );
  fad1_hd mult_x_1_U174 ( .A(mult_x_1_n874), .B(mult_x_1_n563), .CI(
        mult_x_1_n174), .CO(mult_x_1_n173), .S(N181) );
  fad1_hd mult_x_1_U197 ( .A(mult_x_1_n211), .B(mult_x_1_n217), .CI(
        mult_x_1_n215), .CO(mult_x_1_n208), .S(mult_x_1_n209) );
  fad1_hd mult_x_1_U205 ( .A(mult_x_1_n697), .B(mult_x_1_n225), .CI(
        mult_x_1_n232), .CO(mult_x_1_n222), .S(mult_x_1_n223) );
  fad1_hd mult_x_1_U214 ( .A(mult_x_1_n242), .B(mult_x_1_n250), .CI(
        mult_x_1_n723), .CO(mult_x_1_n239), .S(mult_x_1_n240) );
  fad1_hd mult_x_1_U209 ( .A(mult_x_1_n233), .B(mult_x_1_n241), .CI(
        mult_x_1_n239), .CO(mult_x_1_n230), .S(mult_x_1_n231) );
  fad1_hd mult_x_1_U219 ( .A(mult_x_1_n724), .B(mult_x_1_n251), .CI(
        mult_x_1_n260), .CO(mult_x_1_n248), .S(mult_x_1_n249) );
  fad1_hd mult_x_1_U230 ( .A(mult_x_1_n272), .B(mult_x_1_n282), .CI(
        mult_x_1_n750), .CO(mult_x_1_n269), .S(mult_x_1_n270) );
  fad1_hd mult_x_1_U224 ( .A(mult_x_1_n261), .B(mult_x_1_n271), .CI(
        mult_x_1_n269), .CO(mult_x_1_n258), .S(mult_x_1_n259) );
  fad1_hd mult_x_1_U236 ( .A(mult_x_1_n751), .B(mult_x_1_n283), .CI(
        mult_x_1_n294), .CO(mult_x_1_n280), .S(mult_x_1_n281) );
  fad1_hd mult_x_1_U249 ( .A(mult_x_1_n308), .B(mult_x_1_n320), .CI(
        mult_x_1_n777), .CO(mult_x_1_n305), .S(mult_x_1_n306) );
  fad1_hd mult_x_1_U242 ( .A(mult_x_1_n295), .B(mult_x_1_n307), .CI(
        mult_x_1_n305), .CO(mult_x_1_n292), .S(mult_x_1_n293) );
  fad1_hd mult_x_1_U256 ( .A(mult_x_1_n778), .B(mult_x_1_n321), .CI(
        mult_x_1_n334), .CO(mult_x_1_n318), .S(mult_x_1_n319) );
  fad1_hd mult_x_1_U277 ( .A(mult_x_1_n363), .B(mult_x_1_n376), .CI(
        mult_x_1_n805), .CO(mult_x_1_n360), .S(mult_x_1_n361) );
  fad1_hd mult_x_1_U270 ( .A(mult_x_1_n349), .B(mult_x_1_n362), .CI(
        mult_x_1_n360), .CO(mult_x_1_n346), .S(mult_x_1_n347) );
  fad1_hd mult_x_1_U269 ( .A(mult_x_1_n347), .B(mult_x_1_n804), .CI(
        mult_x_1_n828), .CO(mult_x_1_n344), .S(mult_x_1_n345) );
  had1_hd mult_x_1_U375 ( .A(mult_x_1_n824), .B(mult_x_1_n560), .CO(
        mult_x_1_n556), .S(mult_x_1_n557) );
  had1_hd mult_x_1_U373 ( .A(mult_x_1_n823), .B(mult_x_1_n556), .CO(
        mult_x_1_n552), .S(mult_x_1_n553) );
  fad1_hd mult_x_1_U284 ( .A(mult_x_1_n806), .B(mult_x_1_n377), .CI(
        mult_x_1_n388), .CO(mult_x_1_n374), .S(mult_x_1_n375) );
  fad1_hd mult_x_1_U276 ( .A(mult_x_1_n361), .B(mult_x_1_n374), .CI(
        mult_x_1_n829), .CO(mult_x_1_n358), .S(mult_x_1_n359) );
  had1_hd mult_x_1_U379 ( .A(mult_x_1_n851), .B(mult_x_1_n566), .CO(
        mult_x_1_n564), .S(mult_x_1_n565) );
  had1_hd mult_x_1_U378 ( .A(mult_x_1_n850), .B(mult_x_1_n564), .CO(
        mult_x_1_n562), .S(mult_x_1_n563) );
  fad1_hd mult_x_1_U374 ( .A(mult_x_1_n848), .B(mult_x_1_n557), .CI(
        mult_x_1_n558), .CO(mult_x_1_n554), .S(mult_x_1_n555) );
  fad1_hd mult_x_1_U372 ( .A(mult_x_1_n847), .B(mult_x_1_n553), .CI(
        mult_x_1_n554), .CO(mult_x_1_n550), .S(mult_x_1_n551) );
  fad1_hd mult_x_1_U366 ( .A(mult_x_1_n845), .B(mult_x_1_n541), .CI(
        mult_x_1_n544), .CO(mult_x_1_n538), .S(mult_x_1_n539) );
  fad1_hd mult_x_1_U363 ( .A(mult_x_1_n844), .B(mult_x_1_n535), .CI(
        mult_x_1_n538), .CO(mult_x_1_n532), .S(mult_x_1_n533) );
  fad1_hd mult_x_1_U359 ( .A(mult_x_1_n843), .B(mult_x_1_n527), .CI(
        mult_x_1_n532), .CO(mult_x_1_n524), .S(mult_x_1_n525) );
  fad1_hd mult_x_1_U355 ( .A(mult_x_1_n842), .B(mult_x_1_n519), .CI(
        mult_x_1_n524), .CO(mult_x_1_n516), .S(mult_x_1_n517) );
  fad1_hd mult_x_1_U351 ( .A(mult_x_1_n841), .B(mult_x_1_n511), .CI(
        mult_x_1_n516), .CO(mult_x_1_n508), .S(mult_x_1_n509) );
  fad1_hd mult_x_1_U346 ( .A(mult_x_1_n840), .B(mult_x_1_n501), .CI(
        mult_x_1_n508), .CO(mult_x_1_n498), .S(mult_x_1_n499) );
  fad1_hd mult_x_1_U341 ( .A(mult_x_1_n839), .B(mult_x_1_n491), .CI(
        mult_x_1_n498), .CO(mult_x_1_n488), .S(mult_x_1_n489) );
  fad1_hd mult_x_1_U336 ( .A(mult_x_1_n838), .B(mult_x_1_n481), .CI(
        mult_x_1_n488), .CO(mult_x_1_n478), .S(mult_x_1_n479) );
  fad1_hd mult_x_1_U318 ( .A(mult_x_1_n835), .B(mult_x_1_n445), .CI(
        mult_x_1_n454), .CO(mult_x_1_n442), .S(mult_x_1_n443) );
  fad1_hd mult_x_1_U311 ( .A(mult_x_1_n834), .B(mult_x_1_n431), .CI(
        mult_x_1_n442), .CO(mult_x_1_n428), .S(mult_x_1_n429) );
  fad1_hd mult_x_1_U304 ( .A(mult_x_1_n833), .B(mult_x_1_n417), .CI(
        mult_x_1_n428), .CO(mult_x_1_n414), .S(mult_x_1_n415) );
  fad1_hd mult_x_1_U297 ( .A(mult_x_1_n832), .B(mult_x_1_n403), .CI(
        mult_x_1_n414), .CO(mult_x_1_n400), .S(mult_x_1_n401) );
  fad1_hd mult_x_1_U290 ( .A(mult_x_1_n831), .B(mult_x_1_n389), .CI(
        mult_x_1_n400), .CO(mult_x_1_n386), .S(mult_x_1_n387) );
  fad1_hd mult_x_1_U283 ( .A(mult_x_1_n830), .B(mult_x_1_n375), .CI(
        mult_x_1_n386), .CO(mult_x_1_n372), .S(mult_x_1_n373) );
  had1_hd mult_x_1_U178 ( .A(mult_x_1_n878), .B(mult_x_1_n178), .CO(
        mult_x_1_n177), .S(N177) );
  had1_hd mult_x_1_U177 ( .A(mult_x_1_n877), .B(mult_x_1_n177), .CO(
        mult_x_1_n176), .S(N178) );
  fad1_hd mult_x_1_U173 ( .A(mult_x_1_n873), .B(mult_x_1_n559), .CI(
        mult_x_1_n173), .CO(mult_x_1_n172), .S(N182) );
  fad1_hd mult_x_1_U169 ( .A(mult_x_1_n869), .B(mult_x_1_n539), .CI(
        mult_x_1_n169), .CO(mult_x_1_n168), .S(N186) );
  fad1_hd mult_x_1_U168 ( .A(mult_x_1_n868), .B(mult_x_1_n533), .CI(
        mult_x_1_n168), .CO(mult_x_1_n167), .S(N187) );
  fad1_hd mult_x_1_U167 ( .A(mult_x_1_n867), .B(mult_x_1_n525), .CI(
        mult_x_1_n167), .CO(mult_x_1_n166), .S(N188) );
  fad1_hd mult_x_1_U166 ( .A(mult_x_1_n866), .B(mult_x_1_n517), .CI(
        mult_x_1_n166), .CO(mult_x_1_n165), .S(N189) );
  fad1_hd mult_x_1_U165 ( .A(mult_x_1_n865), .B(mult_x_1_n509), .CI(
        mult_x_1_n165), .CO(mult_x_1_n164), .S(N190) );
  fad1_hd mult_x_1_U164 ( .A(mult_x_1_n864), .B(mult_x_1_n499), .CI(
        mult_x_1_n164), .CO(mult_x_1_n163), .S(N191) );
  fad1_hd mult_x_1_U163 ( .A(mult_x_1_n863), .B(mult_x_1_n489), .CI(
        mult_x_1_n163), .CO(mult_x_1_n162), .S(N192) );
  fad1_hd mult_x_1_U194 ( .A(mult_x_1_n670), .B(mult_x_1_n205), .CI(
        mult_x_1_n210), .CO(mult_x_1_n202), .S(mult_x_1_n203) );
  fad1_hd mult_x_1_U201 ( .A(mult_x_1_n218), .B(mult_x_1_n224), .CI(
        mult_x_1_n696), .CO(mult_x_1_n215), .S(mult_x_1_n216) );
  fad1_hd mult_x_1_U218 ( .A(mult_x_1_n258), .B(mult_x_1_n249), .CI(
        mult_x_1_n748), .CO(mult_x_1_n246), .S(mult_x_1_n247) );
  fad1_hd mult_x_1_U229 ( .A(mult_x_1_n270), .B(mult_x_1_n280), .CI(
        mult_x_1_n774), .CO(mult_x_1_n267), .S(mult_x_1_n268) );
  fad1_hd mult_x_1_U223 ( .A(mult_x_1_n259), .B(mult_x_1_n749), .CI(
        mult_x_1_n773), .CO(mult_x_1_n256), .S(mult_x_1_n257) );
  fad1_hd mult_x_1_U159 ( .A(mult_x_1_n859), .B(mult_x_1_n443), .CI(
        mult_x_1_n159), .CO(mult_x_1_n158), .S(N196) );
  fad1_hd mult_x_1_U158 ( .A(mult_x_1_n858), .B(mult_x_1_n429), .CI(
        mult_x_1_n158), .CO(mult_x_1_n157), .S(N197) );
  fad1_hd mult_x_1_U157 ( .A(mult_x_1_n857), .B(mult_x_1_n415), .CI(
        mult_x_1_n157), .CO(mult_x_1_n156), .S(N198) );
  fad1_hd mult_x_1_U156 ( .A(mult_x_1_n856), .B(mult_x_1_n401), .CI(
        mult_x_1_n156), .CO(mult_x_1_n155), .S(N199) );
  fad1_hd mult_x_1_U155 ( .A(mult_x_1_n855), .B(mult_x_1_n387), .CI(
        mult_x_1_n155), .CO(mult_x_1_n154), .S(N200) );
  fad1_hd mult_x_1_U154 ( .A(mult_x_1_n373), .B(mult_x_1_n854), .CI(
        mult_x_1_n154), .CO(mult_x_1_n153), .S(N201) );
  fad1_hd mult_x_1_U153 ( .A(mult_x_1_n359), .B(mult_x_1_n372), .CI(
        mult_x_1_n153), .CO(mult_x_1_n152), .S(N202) );
  fad1_hd mult_x_1_U181 ( .A(mult_x_1_n185), .B(mult_x_1_n569), .CI(
        mult_x_1_n665), .CO(mult_x_1_n180), .S(mult_x_1_n181) );
  fad1_hd mult_x_1_U183 ( .A(mult_x_1_n188), .B(mult_x_1_n185), .CI(
        mult_x_1_n666), .CO(mult_x_1_n183), .S(mult_x_1_n184) );
  fad1_hd mult_x_1_U188 ( .A(mult_x_1_n194), .B(n884), .CI(mult_x_1_n197), 
        .CO(mult_x_1_n192), .S(mult_x_1_n193) );
  fad1_hd mult_x_1_U204 ( .A(mult_x_1_n230), .B(mult_x_1_n223), .CI(
        mult_x_1_n721), .CO(mult_x_1_n220), .S(mult_x_1_n221) );
  fad1_hd mult_x_1_U213 ( .A(mult_x_1_n240), .B(mult_x_1_n248), .CI(
        mult_x_1_n747), .CO(mult_x_1_n237), .S(mult_x_1_n238) );
  fad1_hd mult_x_1_U208 ( .A(mult_x_1_n231), .B(mult_x_1_n722), .CI(
        mult_x_1_n746), .CO(mult_x_1_n228), .S(mult_x_1_n229) );
  fad1_hd mult_x_1_U185 ( .A(mult_x_1_n192), .B(mult_x_1_n189), .CI(
        mult_x_1_n667), .CO(mult_x_1_n186), .S(mult_x_1_n187) );
  fad1_hd mult_x_1_U187 ( .A(mult_x_1_n193), .B(mult_x_1_n668), .CI(
        mult_x_1_n692), .CO(mult_x_1_n190), .S(mult_x_1_n191) );
  fad1_hd mult_x_1_U191 ( .A(mult_x_1_n204), .B(mult_x_1_n199), .CI(
        mult_x_1_n669), .CO(mult_x_1_n197), .S(mult_x_1_n198) );
  fad1_hd mult_x_1_U190 ( .A(mult_x_1_n198), .B(mult_x_1_n202), .CI(
        mult_x_1_n693), .CO(mult_x_1_n195), .S(mult_x_1_n196) );
  fad1_hd mult_x_1_U193 ( .A(mult_x_1_n208), .B(mult_x_1_n203), .CI(
        mult_x_1_n694), .CO(mult_x_1_n200), .S(mult_x_1_n201) );
  fad1_hd mult_x_1_U196 ( .A(mult_x_1_n209), .B(mult_x_1_n695), .CI(
        mult_x_1_n719), .CO(mult_x_1_n206), .S(mult_x_1_n207) );
  fad1_hd mult_x_1_U200 ( .A(mult_x_1_n216), .B(mult_x_1_n222), .CI(
        mult_x_1_n720), .CO(mult_x_1_n213), .S(mult_x_1_n214) );
  fad1_hd mult_x_1_U1162 ( .A(n1031), .B(n1026), .CI(mult_x_1_n633), .CO(
        mult_x_1_n632), .S(mult_x_1_n657) );
  fad1_hd mult_x_1_U1163 ( .A(n1036), .B(n1031), .CI(mult_x_1_n634), .CO(
        mult_x_1_n633), .S(mult_x_1_n658) );
  fad1_hd mult_x_1_U1164 ( .A(n1041), .B(n1036), .CI(mult_x_1_n635), .CO(
        mult_x_1_n634), .S(mult_x_1_n659) );
  fad1_hd mult_x_1_U1165 ( .A(n1046), .B(n1041), .CI(mult_x_1_n636), .CO(
        mult_x_1_n635), .S(mult_x_1_n660) );
  fad1_hd mult_x_1_U1166 ( .A(n1051), .B(n1046), .CI(mult_x_1_n637), .CO(
        mult_x_1_n636), .S(mult_x_1_n661) );
  fad1_hd mult_x_1_U1167 ( .A(n1056), .B(n1051), .CI(mult_x_1_n638), .CO(
        mult_x_1_n637), .S(mult_x_1_n662) );
  had1_hd mult_x_1_U1168 ( .A(n1056), .B(n483), .CO(mult_x_1_n638), .S(
        mult_x_1_n663) );
  xo2d1_hd DP_OP_125J2_130_6300_U23 ( .A(a_e[9]), .B(b_e[9]), .Y(
        DP_OP_125J2_130_6300_n11) );
  scg2d1_hd DP_OP_125J2_130_6300_U20 ( .A(DP_OP_125J2_130_6300_n35), .B(n580), 
        .C(n467), .D(z_e[1]), .Y(DP_OP_125J2_130_6300_n25) );
  scg2d1_hd DP_OP_125J2_130_6300_U19 ( .A(DP_OP_125J2_130_6300_n36), .B(n580), 
        .C(n466), .D(z_e[2]), .Y(DP_OP_125J2_130_6300_n26) );
  scg2d1_hd DP_OP_125J2_130_6300_U18 ( .A(DP_OP_125J2_130_6300_n37), .B(n580), 
        .C(n467), .D(z_e[3]), .Y(DP_OP_125J2_130_6300_n27) );
  scg2d1_hd DP_OP_125J2_130_6300_U17 ( .A(DP_OP_125J2_130_6300_n38), .B(n581), 
        .C(n466), .D(z_e[4]), .Y(DP_OP_125J2_130_6300_n28) );
  scg2d1_hd DP_OP_125J2_130_6300_U16 ( .A(DP_OP_125J2_130_6300_n39), .B(n581), 
        .C(n467), .D(z_e[5]), .Y(DP_OP_125J2_130_6300_n29) );
  scg2d1_hd DP_OP_125J2_130_6300_U15 ( .A(DP_OP_125J2_130_6300_n40), .B(n581), 
        .C(n466), .D(z_e[6]), .Y(DP_OP_125J2_130_6300_n30) );
  scg2d1_hd DP_OP_125J2_130_6300_U14 ( .A(DP_OP_125J2_130_6300_n41), .B(n581), 
        .C(n467), .D(z_e[7]), .Y(DP_OP_125J2_130_6300_n31) );
  scg2d1_hd DP_OP_125J2_130_6300_U13 ( .A(DP_OP_125J2_130_6300_n42), .B(n581), 
        .C(n466), .D(z_e[8]), .Y(DP_OP_125J2_130_6300_n32) );
  scg2d1_hd DP_OP_125J2_130_6300_U21 ( .A(DP_OP_125J2_130_6300_n34), .B(n580), 
        .C(n466), .D(z_e[0]), .Y(DP_OP_125J2_130_6300_n10) );
  scg2d1_hd DP_OP_125J2_130_6300_U12 ( .A(DP_OP_125J2_130_6300_n43), .B(n581), 
        .C(n467), .D(z_e[9]), .Y(DP_OP_125J2_130_6300_n33) );
  xo2d1_hd DP_OP_125J2_130_6300_U22 ( .A(DP_OP_125J2_130_6300_n12), .B(
        DP_OP_125J2_130_6300_n11), .Y(DP_OP_125J2_130_6300_n43) );
  xo2d1_hd DP_OP_125J2_130_6300_U1 ( .A(DP_OP_125J2_130_6300_n1), .B(
        DP_OP_125J2_130_6300_n2), .Y(N475) );
  fad1_hd mult_x_1_U235 ( .A(mult_x_1_n292), .B(mult_x_1_n281), .CI(
        mult_x_1_n775), .CO(mult_x_1_n278), .S(mult_x_1_n279) );
  fad1_hd mult_x_1_U241 ( .A(mult_x_1_n293), .B(mult_x_1_n776), .CI(
        mult_x_1_n800), .CO(mult_x_1_n290), .S(mult_x_1_n291) );
  fad1_hd mult_x_1_U263 ( .A(mult_x_1_n335), .B(mult_x_1_n348), .CI(
        mult_x_1_n346), .CO(mult_x_1_n332), .S(mult_x_1_n333) );
  fad1_hd mult_x_1_U262 ( .A(mult_x_1_n333), .B(mult_x_1_n803), .CI(
        mult_x_1_n827), .CO(mult_x_1_n330), .S(mult_x_1_n331) );
  fad1_hd mult_x_1_U255 ( .A(mult_x_1_n332), .B(mult_x_1_n319), .CI(
        mult_x_1_n802), .CO(mult_x_1_n316), .S(mult_x_1_n317) );
  fad1_hd mult_x_1_U248 ( .A(mult_x_1_n306), .B(mult_x_1_n318), .CI(
        mult_x_1_n801), .CO(mult_x_1_n303), .S(mult_x_1_n304) );
  fad1_hd mult_x_1_U1150 ( .A(n971), .B(n966), .CI(mult_x_1_n621), .CO(
        mult_x_1_n620), .S(mult_x_1_n645) );
  fad1_hd mult_x_1_U1149 ( .A(n966), .B(n961), .CI(mult_x_1_n620), .CO(
        mult_x_1_n619), .S(mult_x_1_n644) );
  fad1_hd mult_x_1_U1148 ( .A(n961), .B(n956), .CI(mult_x_1_n619), .CO(
        mult_x_1_n618), .S(mult_x_1_n643) );
  fad1_hd mult_x_1_U1147 ( .A(n956), .B(n486), .CI(mult_x_1_n618), .CO(
        mult_x_1_n617), .S(mult_x_1_n642) );
  fad1_hd mult_x_1_U1154 ( .A(n991), .B(n986), .CI(mult_x_1_n625), .CO(
        mult_x_1_n624), .S(mult_x_1_n649) );
  fad1_hd mult_x_1_U1153 ( .A(n986), .B(n981), .CI(mult_x_1_n624), .CO(
        mult_x_1_n623), .S(mult_x_1_n648) );
  fad1_hd mult_x_1_U1152 ( .A(n981), .B(n976), .CI(mult_x_1_n623), .CO(
        mult_x_1_n622), .S(mult_x_1_n647) );
  fad1_hd mult_x_1_U1151 ( .A(n976), .B(n971), .CI(mult_x_1_n622), .CO(
        mult_x_1_n621), .S(mult_x_1_n646) );
  fd1qd1_hd b_m_reg_0_ ( .D(n308), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n358), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd a_m_reg_0_ ( .D(n349), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n310), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n355), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n350), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd sticky_reg ( .D(n283), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd b_m_reg_21_ ( .D(n309), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n306), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n290), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n291), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n292), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n295), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n296), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n299), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n305), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n294), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n332), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n344), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n329), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n336), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n346), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n331), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n330), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n333), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n337), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n340), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd z_reg_22_ ( .D(n238), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd z_reg_28_ ( .D(n232), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n234), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_29_ ( .D(n231), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_24_ ( .D(n236), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n237), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n289), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n297), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n298), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n302), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n301), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n287), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd z_reg_27_ ( .D(n233), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n235), .CK(i_CLK), .Q(z[25]) );
  fd1qd1_hd z_reg_30_ ( .D(n230), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n338), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n304), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n293), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n303), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n307), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n300), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd z_reg_17_ ( .D(n243), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n244), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_20_ ( .D(n240), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_18_ ( .D(n242), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_15_ ( .D(n245), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n246), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n335), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n339), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n342), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n343), .CK(i_CLK), .Q(a_m[6]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n354), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n341), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd z_reg_1_ ( .D(n259), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_0_ ( .D(n260), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_21_ ( .D(n239), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_2_ ( .D(n258), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n345), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n334), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n348), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n347), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd z_reg_31_ ( .D(n229), .CK(i_CLK), .Q(z[31]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n288), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n328), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n326), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n317), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd z_reg_13_ ( .D(n247), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n248), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_9_ ( .D(n251), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n252), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_5_ ( .D(n255), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_4_ ( .D(n256), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_19_ ( .D(n241), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_11_ ( .D(n249), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n250), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_7_ ( .D(n253), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n254), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_3_ ( .D(n257), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd round_bit_reg ( .D(n284), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd b_e_reg_0_ ( .D(n327), .CK(i_CLK), .Q(b_e[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n318), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n325), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n316), .CK(i_CLK), .Q(a_e[2]) );
  fd1qd1_hd state_reg_3_ ( .D(n357), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd state_reg_2_ ( .D(n351), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_0_ ( .D(n353), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd state_reg_1_ ( .D(n352), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n315), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n324), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n323), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n314), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n282), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n322), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n313), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n281), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n285), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n312), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n321), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n262), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n276), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n264), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n280), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n268), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n272), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n261), .CK(i_CLK), .Q(z_m[22]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n270), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n266), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n274), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n278), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n269), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n265), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n277), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n273), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n275), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n267), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n279), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n271), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n263), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n286), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n320), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n311), .CK(i_CLK), .Q(a_e[8]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n380), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n380), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n370), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n1165), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n386), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n384), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n373), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n386), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n374), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n379), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n379), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n378), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n369), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n372), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n384), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n1168), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n371), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1165), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n370), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n380), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd product_reg_2_ ( .D(N176), .E(n383), .CK(i_CLK), .Q(product[2])
         );
  fd1eqd1_hd z_s_reg ( .D(N35), .E(n383), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n370), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n369), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n369), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n379), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n378), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n370), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n370), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n369), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n380), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n378), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n378), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n369), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n386), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n1167), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n374), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n1168), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n372), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n379), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n380), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n380), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n370), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n1165), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n379), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n379), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n378), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n369), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1332), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1332), .CK(i_CLK), .Q(a_s) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n385), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n385), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n385), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n371), .CK(i_CLK), .Q(b[28]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n385), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n374), .CK(i_CLK), .Q(b[26]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n1169), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n371), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n1166), .CK(i_CLK), .Q(b[23]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n1168), .CK(i_CLK), .Q(b[22]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n1166), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n1167), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n384), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n373), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n1169), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n385), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n372), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n374), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n1169), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n372), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n1166), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n384), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n368), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n1167), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n368), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n372), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n1169), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n1169), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n386), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n373), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n368), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n373), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n368), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n368), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n373), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n373), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n368), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n384), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n1166), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n371), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd guard_reg ( .D(n104), .E(n105), .CK(i_CLK), .Q(net908) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n1168), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n374), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n374), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n386), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n1167), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n1168), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n371), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n1166), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n385), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n386), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd product_reg_3_ ( .D(N177), .E(n381), .CK(i_CLK), .Q(product[3])
         );
  fd1eqd1_hd product_reg_4_ ( .D(N178), .E(n377), .CK(i_CLK), .Q(product[4])
         );
  fd1eqd1_hd product_reg_5_ ( .D(N179), .E(n376), .CK(i_CLK), .Q(product[5])
         );
  fd1eqd1_hd product_reg_6_ ( .D(N180), .E(n383), .CK(i_CLK), .Q(product[6])
         );
  fd1eqd1_hd product_reg_7_ ( .D(N181), .E(n1128), .CK(i_CLK), .Q(product[7])
         );
  fd1eqd1_hd product_reg_8_ ( .D(N182), .E(n375), .CK(i_CLK), .Q(product[8])
         );
  fd1eqd1_hd z_e_reg_7_ ( .D(N473), .E(n469), .CK(i_CLK), .Q(z_e[7]) );
  fd1eqd1_hd z_e_reg_6_ ( .D(N472), .E(n468), .CK(i_CLK), .Q(z_e[6]) );
  fd1eqd1_hd z_e_reg_5_ ( .D(N471), .E(n468), .CK(i_CLK), .Q(z_e[5]) );
  fd1eqd1_hd z_e_reg_4_ ( .D(N470), .E(n469), .CK(i_CLK), .Q(z_e[4]) );
  fd1eqd1_hd z_e_reg_3_ ( .D(N469), .E(n469), .CK(i_CLK), .Q(z_e[3]) );
  fd1eqd1_hd z_e_reg_2_ ( .D(N468), .E(n469), .CK(i_CLK), .Q(z_e[2]) );
  fd1eqd1_hd z_e_reg_1_ ( .D(N467), .E(n468), .CK(i_CLK), .Q(z_e[1]) );
  fd1eqd1_hd z_e_reg_0_ ( .D(N466), .E(n468), .CK(i_CLK), .Q(z_e[0]) );
  fd1eqd1_hd z_e_reg_8_ ( .D(N474), .E(n468), .CK(i_CLK), .Q(z_e[8]) );
  fd1eqd1_hd product_reg_9_ ( .D(N183), .E(n375), .CK(i_CLK), .Q(product[9])
         );
  fd1eqd1_hd z_e_reg_9_ ( .D(N475), .E(n469), .CK(i_CLK), .Q(z_e[9]) );
  fd1eqd1_hd product_reg_10_ ( .D(N184), .E(n1214), .CK(i_CLK), .Q(product[10]) );
  fd1eqd1_hd product_reg_11_ ( .D(N185), .E(n1129), .CK(i_CLK), .Q(product[11]) );
  fd1eqd1_hd product_reg_12_ ( .D(N186), .E(n381), .CK(i_CLK), .Q(product[12])
         );
  fd1eqd1_hd product_reg_13_ ( .D(N187), .E(n376), .CK(i_CLK), .Q(product[13])
         );
  fd1eqd1_hd product_reg_14_ ( .D(N188), .E(n1129), .CK(i_CLK), .Q(product[14]) );
  fd1eqd1_hd product_reg_15_ ( .D(N189), .E(n1128), .CK(i_CLK), .Q(product[15]) );
  fd1eqd1_hd product_reg_16_ ( .D(N190), .E(n1129), .CK(i_CLK), .Q(product[16]) );
  fd1eqd1_hd product_reg_17_ ( .D(N191), .E(n377), .CK(i_CLK), .Q(product[17])
         );
  fd1eqd1_hd product_reg_18_ ( .D(N192), .E(n376), .CK(i_CLK), .Q(product[18])
         );
  fd1eqd1_hd product_reg_19_ ( .D(N193), .E(n1128), .CK(i_CLK), .Q(product[19]) );
  fd1eqd1_hd product_reg_20_ ( .D(N194), .E(DP_OP_125J2_130_6300_I3), .CK(
        i_CLK), .Q(product[20]) );
  fd1eqd1_hd product_reg_21_ ( .D(N195), .E(n381), .CK(i_CLK), .Q(product[21])
         );
  fd1eqd1_hd product_reg_22_ ( .D(N196), .E(n375), .CK(i_CLK), .Q(product[22])
         );
  fd1eqd1_hd product_reg_23_ ( .D(N197), .E(n383), .CK(i_CLK), .Q(product[23])
         );
  fd1eqd1_hd product_reg_24_ ( .D(N198), .E(n1214), .CK(i_CLK), .Q(product[24]) );
  fd1eqd1_hd product_reg_25_ ( .D(N199), .E(DP_OP_125J2_130_6300_I3), .CK(
        i_CLK), .Q(product[25]) );
  fd1eqd1_hd product_reg_26_ ( .D(N200), .E(n376), .CK(i_CLK), .Q(product[26])
         );
  fd1eqd1_hd product_reg_27_ ( .D(N201), .E(n377), .CK(i_CLK), .Q(product[27])
         );
  fd1eqd1_hd product_reg_28_ ( .D(N202), .E(n377), .CK(i_CLK), .Q(product[28])
         );
  fd1eqd1_hd product_reg_29_ ( .D(N203), .E(n1127), .CK(i_CLK), .Q(product[29]) );
  fd1eqd1_hd product_reg_30_ ( .D(N204), .E(n381), .CK(i_CLK), .Q(product[30])
         );
  fd1eqd1_hd product_reg_31_ ( .D(N205), .E(n377), .CK(i_CLK), .Q(product[31])
         );
  fd1eqd1_hd product_reg_32_ ( .D(N206), .E(n1214), .CK(i_CLK), .Q(product[32]) );
  fd1eqd1_hd product_reg_33_ ( .D(N207), .E(n1129), .CK(i_CLK), .Q(product[33]) );
  fd1eqd1_hd product_reg_34_ ( .D(N208), .E(n1127), .CK(i_CLK), .Q(product[34]) );
  fd1eqd1_hd product_reg_35_ ( .D(N209), .E(n375), .CK(i_CLK), .Q(product[35])
         );
  fd1eqd1_hd product_reg_36_ ( .D(N210), .E(n375), .CK(i_CLK), .Q(product[36])
         );
  fd1eqd1_hd product_reg_37_ ( .D(N211), .E(n1129), .CK(i_CLK), .Q(product[37]) );
  fd1eqd1_hd product_reg_38_ ( .D(N212), .E(n1127), .CK(i_CLK), .Q(product[38]) );
  fd1eqd1_hd product_reg_39_ ( .D(N213), .E(n1127), .CK(i_CLK), .Q(product[39]) );
  fd1eqd1_hd product_reg_40_ ( .D(N214), .E(n376), .CK(i_CLK), .Q(product[40])
         );
  fd1eqd1_hd product_reg_41_ ( .D(N215), .E(n1128), .CK(i_CLK), .Q(product[41]) );
  fd1eqd1_hd product_reg_42_ ( .D(N216), .E(n1128), .CK(i_CLK), .Q(product[42]) );
  fd1eqd1_hd product_reg_43_ ( .D(N217), .E(n580), .CK(i_CLK), .Q(product[43])
         );
  fd1eqd1_hd product_reg_44_ ( .D(N218), .E(n377), .CK(i_CLK), .Q(product[44])
         );
  fd1eqd1_hd product_reg_45_ ( .D(N219), .E(n376), .CK(i_CLK), .Q(product[45])
         );
  fd1eqd1_hd product_reg_46_ ( .D(N220), .E(n383), .CK(i_CLK), .Q(product[46])
         );
  fd1eqd1_hd product_reg_47_ ( .D(N221), .E(DP_OP_125J2_130_6300_I3), .CK(
        i_CLK), .Q(product[47]) );
  fd1eqd1_hd product_reg_48_ ( .D(N222), .E(n383), .CK(i_CLK), .Q(product[48])
         );
  fd1eqd1_hd product_reg_49_ ( .D(N223), .E(n375), .CK(i_CLK), .Q(product[49])
         );
  fad2_hd U367 ( .A(mult_x_1_n184), .B(mult_x_1_n186), .CI(mult_x_1_n134), 
        .CO(mult_x_1_n133), .S(N221) );
  fad2_hd U368 ( .A(mult_x_1_n344), .B(mult_x_1_n331), .CI(mult_x_1_n151), 
        .CO(mult_x_1_n150), .S(N204) );
  fad2_hd U369 ( .A(mult_x_1_n330), .B(mult_x_1_n317), .CI(mult_x_1_n150), 
        .CO(mult_x_1_n149), .S(N205) );
  fad2_hd U370 ( .A(mult_x_1_n862), .B(mult_x_1_n479), .CI(mult_x_1_n162), 
        .CO(mult_x_1_n161), .S(N193) );
  fad2_hd U371 ( .A(mult_x_1_n861), .B(mult_x_1_n467), .CI(mult_x_1_n161), 
        .CO(mult_x_1_n160), .S(N194) );
  fad1_hd U372 ( .A(mult_x_1_n837), .B(mult_x_1_n469), .CI(mult_x_1_n478), 
        .CO(mult_x_1_n466), .S(mult_x_1_n467) );
  fad2_hd U373 ( .A(mult_x_1_n237), .B(mult_x_1_n229), .CI(mult_x_1_n142), 
        .CO(mult_x_1_n141), .S(N213) );
  fad2_hd U374 ( .A(mult_x_1_n860), .B(mult_x_1_n455), .CI(mult_x_1_n160), 
        .CO(mult_x_1_n159), .S(N195) );
  fad2_hd U375 ( .A(mult_x_1_n871), .B(mult_x_1_n551), .CI(mult_x_1_n171), 
        .CO(mult_x_1_n170), .S(N184) );
  ao22d1_hd U376 ( .A(n945), .B(n863), .C(a_m[1]), .D(n940), .Y(n831) );
  clknd2d1_hd U377 ( .A(n453), .B(n1123), .Y(n828) );
  nr2d1_hd U378 ( .A(n831), .B(n387), .Y(n857) );
  ivd1_hd U379 ( .A(a_m[2]), .Y(n939) );
  fad1_hd U380 ( .A(mult_x_1_n836), .B(mult_x_1_n457), .CI(mult_x_1_n466), 
        .CO(mult_x_1_n454), .S(mult_x_1_n455) );
  fad1_hd U381 ( .A(mult_x_1_n846), .B(mult_x_1_n547), .CI(mult_x_1_n550), 
        .CO(mult_x_1_n544), .S(mult_x_1_n545) );
  ivd1_hd U382 ( .A(n939), .Y(n945) );
  fad2_hd U383 ( .A(mult_x_1_n183), .B(mult_x_1_n181), .CI(mult_x_1_n133), 
        .CO(mult_x_1_n132), .S(N222) );
  fad1_hd U384 ( .A(mult_x_1_n228), .B(mult_x_1_n221), .CI(mult_x_1_n141), 
        .CO(mult_x_1_n140), .S(N214) );
  fad1_hd U385 ( .A(mult_x_1_n345), .B(mult_x_1_n358), .CI(mult_x_1_n152), 
        .CO(mult_x_1_n151), .S(N203) );
  fad1_hd U386 ( .A(mult_x_1_n870), .B(mult_x_1_n545), .CI(mult_x_1_n170), 
        .CO(mult_x_1_n169), .S(N185) );
  fad4_hd U387 ( .A(mult_x_1_n872), .B(mult_x_1_n555), .CI(mult_x_1_n172), 
        .CO(mult_x_1_n171), .S(N183) );
  nid1_hd U388 ( .A(n751), .Y(n1093) );
  nid1_hd U389 ( .A(n786), .Y(n1101) );
  clknd2d1_hd U390 ( .A(n453), .B(n1106), .Y(n759) );
  nid1_hd U391 ( .A(n855), .Y(n1121) );
  nid1_hd U392 ( .A(n1063), .Y(n1064) );
  clknd2d1_hd U393 ( .A(n892), .B(n1026), .Y(mult_x_1_n302) );
  clknd2d1_hd U394 ( .A(n891), .B(n1031), .Y(mult_x_1_n315) );
  clknd2d1_hd U395 ( .A(n891), .B(n1018), .Y(mult_x_1_n277) );
  nid1_hd U396 ( .A(n1059), .Y(n1061) );
  clknd2d1_hd U397 ( .A(n891), .B(n998), .Y(mult_x_1_n236) );
  clknd2d1_hd U398 ( .A(n891), .B(n1003), .Y(mult_x_1_n245) );
  nid1_hd U399 ( .A(n1074), .Y(n1072) );
  nid1_hd U400 ( .A(n1082), .Y(n1080) );
  ivd1_hd U401 ( .A(n887), .Y(n896) );
  ivd1_hd U402 ( .A(n898), .Y(n903) );
  clknd2d1_hd U403 ( .A(n891), .B(n986), .Y(mult_x_1_n219) );
  nid1_hd U404 ( .A(n904), .Y(n905) );
  ivd1_hd U405 ( .A(n905), .Y(n910) );
  nid1_hd U406 ( .A(n611), .Y(n1062) );
  nid1_hd U407 ( .A(n1066), .Y(n1065) );
  nid1_hd U408 ( .A(n911), .Y(n912) );
  ivd1_hd U409 ( .A(n912), .Y(n917) );
  nid1_hd U410 ( .A(n918), .Y(n919) );
  nid1_hd U411 ( .A(n1078), .Y(n1076) );
  nid1_hd U412 ( .A(n1090), .Y(n1088) );
  nid1_hd U413 ( .A(n1086), .Y(n1084) );
  ivd1_hd U414 ( .A(n919), .Y(n924) );
  nid1_hd U415 ( .A(n897), .Y(n898) );
  ao22d1_hd U416 ( .A(n903), .B(n876), .C(a_m[21]), .D(n898), .Y(n615) );
  nid1_hd U417 ( .A(n1062), .Y(n1059) );
  clknd2d1_hd U418 ( .A(n890), .B(n966), .Y(mult_x_1_n194) );
  clknd2d1_hd U419 ( .A(n891), .B(n971), .Y(mult_x_1_n199) );
  nid1_hd U420 ( .A(n1074), .Y(n1071) );
  nid1_hd U421 ( .A(n1066), .Y(n1063) );
  nid1_hd U422 ( .A(n1082), .Y(n1079) );
  nid1_hd U423 ( .A(n648), .Y(n1074) );
  nid1_hd U424 ( .A(n1090), .Y(n1087) );
  nid1_hd U425 ( .A(n683), .Y(n1082) );
  nid1_hd U426 ( .A(n1098), .Y(n1095) );
  nid1_hd U427 ( .A(n718), .Y(n1090) );
  nid1_hd U428 ( .A(n753), .Y(n1098) );
  nid1_hd U429 ( .A(n994), .Y(n996) );
  nid1_hd U430 ( .A(n1102), .Y(n1100) );
  nid1_hd U431 ( .A(n999), .Y(n1001) );
  ivd1_hd U432 ( .A(n926), .Y(n931) );
  nid1_hd U433 ( .A(n886), .Y(n887) );
  nid1_hd U434 ( .A(n612), .Y(n1066) );
  nr2bd1_hd U435 ( .AN(n615), .B(n583), .Y(n611) );
  clknd2d1_hd U436 ( .A(mult_x_1_n640), .B(n612), .Y(n585) );
  clknd2d1_hd U437 ( .A(n892), .B(n956), .Y(mult_x_1_n185) );
  nr2bd1_hd U438 ( .AN(n588), .B(n615), .Y(n612) );
  nid1_hd U439 ( .A(n1059), .Y(n1060) );
  clknd2d1_hd U440 ( .A(n453), .B(n1073), .Y(n619) );
  nid1_hd U441 ( .A(n1071), .Y(n1073) );
  nid1_hd U442 ( .A(n1070), .Y(n1067) );
  clknd2d1_hd U443 ( .A(mult_x_1_n640), .B(n1081), .Y(n654) );
  nid1_hd U444 ( .A(n1079), .Y(n1081) );
  nid1_hd U445 ( .A(n1078), .Y(n1075) );
  clknd2d1_hd U446 ( .A(n453), .B(n1089), .Y(n689) );
  nid1_hd U447 ( .A(n1087), .Y(n1089) );
  nid1_hd U448 ( .A(n1086), .Y(n1083) );
  clknd2d1_hd U449 ( .A(mult_x_1_n640), .B(n1097), .Y(n724) );
  nid1_hd U450 ( .A(n1094), .Y(n1091) );
  nid1_hd U451 ( .A(n1102), .Y(n1099) );
  clknd2d1_hd U452 ( .A(n951), .B(n1110), .Y(n795) );
  clknd2d1_hd U453 ( .A(mult_x_1_n640), .B(n1114), .Y(n794) );
  ivd1_hd U454 ( .A(n485), .Y(n486) );
  nid1_hd U455 ( .A(n957), .Y(n954) );
  nid1_hd U456 ( .A(b_m[21]), .Y(n958) );
  nid1_hd U457 ( .A(b_m[20]), .Y(n963) );
  nid1_hd U458 ( .A(b_m[19]), .Y(n968) );
  nid1_hd U459 ( .A(b_m[18]), .Y(n973) );
  nid1_hd U460 ( .A(n993), .Y(n989) );
  nid1_hd U461 ( .A(b_m[17]), .Y(n978) );
  nid1_hd U462 ( .A(b_m[16]), .Y(n983) );
  nid1_hd U463 ( .A(b_m[15]), .Y(n988) );
  nid1_hd U464 ( .A(n1004), .Y(n1006) );
  nid1_hd U465 ( .A(n1023), .Y(n1020) );
  nid1_hd U466 ( .A(n1107), .Y(n1109) );
  nid1_hd U467 ( .A(b_m[8]), .Y(n1023) );
  nid1_hd U468 ( .A(b_m[7]), .Y(n1028) );
  nid1_hd U469 ( .A(n1107), .Y(n1110) );
  nid1_hd U470 ( .A(b_m[5]), .Y(n1038) );
  nid1_hd U471 ( .A(n823), .Y(n1114) );
  nid1_hd U472 ( .A(b_m[4]), .Y(n1043) );
  nid1_hd U473 ( .A(b_m[1]), .Y(n1058) );
  nid1_hd U474 ( .A(b_m[2]), .Y(n1053) );
  clknd2d1_hd U475 ( .A(n831), .B(n388), .Y(n856) );
  clknd2d1_hd U476 ( .A(state[0]), .B(n1219), .Y(n1368) );
  clknd2d1_hd U477 ( .A(state[2]), .B(n1304), .Y(n1172) );
  nid1_hd U478 ( .A(n1140), .Y(n1131) );
  clknd2d1_hd U479 ( .A(state[1]), .B(n1303), .Y(n1258) );
  clknd2d1_hd U480 ( .A(n1254), .B(n1253), .Y(n1364) );
  clknd2d1_hd U481 ( .A(z_e[8]), .B(z_e[7]), .Y(n1365) );
  clknd2d1_hd U482 ( .A(n34), .B(n1219), .Y(n1394) );
  clknd2d1_hd U483 ( .A(state[1]), .B(n1304), .Y(n1290) );
  nid1_hd U484 ( .A(n1140), .Y(n1130) );
  clknd2d1_hd U485 ( .A(n950), .B(n611), .Y(n584) );
  clknd2d1_hd U486 ( .A(n950), .B(n1069), .Y(n620) );
  clknd2d1_hd U487 ( .A(n950), .B(n1077), .Y(n655) );
  clknd2d1_hd U488 ( .A(n950), .B(n1085), .Y(n690) );
  clknd2d1_hd U489 ( .A(n950), .B(n1093), .Y(n725) );
  clknd2d1_hd U490 ( .A(n950), .B(n1101), .Y(n760) );
  ivd1_hd U491 ( .A(n947), .Y(n952) );
  nid1_hd U492 ( .A(n958), .Y(n956) );
  nid1_hd U493 ( .A(n967), .Y(n964) );
  nid1_hd U494 ( .A(n958), .Y(n955) );
  nid1_hd U495 ( .A(n963), .Y(n961) );
  nid1_hd U496 ( .A(n968), .Y(n966) );
  nid1_hd U497 ( .A(n972), .Y(n969) );
  nid1_hd U498 ( .A(n963), .Y(n960) );
  nid1_hd U499 ( .A(n973), .Y(n971) );
  nid1_hd U500 ( .A(n977), .Y(n974) );
  nid1_hd U501 ( .A(n968), .Y(n965) );
  nid1_hd U502 ( .A(n978), .Y(n976) );
  nid1_hd U503 ( .A(n982), .Y(n979) );
  nid1_hd U504 ( .A(n973), .Y(n970) );
  nid1_hd U505 ( .A(n983), .Y(n981) );
  nid1_hd U506 ( .A(n978), .Y(n975) );
  nid1_hd U507 ( .A(n987), .Y(n984) );
  nid1_hd U508 ( .A(n988), .Y(n986) );
  nid1_hd U509 ( .A(n983), .Y(n980) );
  nid1_hd U510 ( .A(n993), .Y(n991) );
  nid1_hd U511 ( .A(n988), .Y(n985) );
  nid1_hd U512 ( .A(b_m[13]), .Y(n998) );
  nid1_hd U513 ( .A(n993), .Y(n990) );
  nid1_hd U514 ( .A(b_m[12]), .Y(n1003) );
  nid1_hd U515 ( .A(b_m[11]), .Y(n1008) );
  nid1_hd U516 ( .A(b_m[10]), .Y(n1013) );
  nid1_hd U517 ( .A(b_m[9]), .Y(n1018) );
  nid1_hd U518 ( .A(n1023), .Y(n1019) );
  nid1_hd U519 ( .A(n1023), .Y(n1022) );
  nid1_hd U520 ( .A(n1028), .Y(n1026) );
  nid1_hd U521 ( .A(n1023), .Y(n1021) );
  nid1_hd U522 ( .A(n1033), .Y(n1031) );
  nid1_hd U523 ( .A(n1028), .Y(n1025) );
  nid1_hd U524 ( .A(DP_OP_125J2_130_6300_I3), .Y(n581) );
  nid1_hd U525 ( .A(n1038), .Y(n1036) );
  nid1_hd U526 ( .A(n1043), .Y(n1041) );
  nid1_hd U527 ( .A(n1038), .Y(n1035) );
  nid1_hd U528 ( .A(n1048), .Y(n1046) );
  nid1_hd U529 ( .A(n1043), .Y(n1040) );
  nid1_hd U530 ( .A(n1058), .Y(n1055) );
  nid1_hd U531 ( .A(n1053), .Y(n1051) );
  nid1_hd U532 ( .A(n1048), .Y(n1045) );
  nid1_hd U533 ( .A(n1118), .Y(n1117) );
  nid1_hd U534 ( .A(n1058), .Y(n1056) );
  nid1_hd U535 ( .A(n1053), .Y(n1050) );
  nid1_hd U536 ( .A(n1118), .Y(n1115) );
  nid1_hd U537 ( .A(n1057), .Y(n1054) );
  nid1_hd U538 ( .A(n1122), .Y(n1119) );
  clknd2d1_hd U539 ( .A(n572), .B(n1373), .Y(n1378) );
  clknd2d1_hd U540 ( .A(z_m[21]), .B(n1478), .Y(n1488) );
  clknd2d1_hd U541 ( .A(n477), .B(n1437), .Y(n1442) );
  clknd2d1_hd U542 ( .A(n475), .B(n1452), .Y(n1457) );
  clknd2d1_hd U543 ( .A(n475), .B(n1407), .Y(n1412) );
  clknd2d1_hd U544 ( .A(n476), .B(n1469), .Y(n1473) );
  nid1_hd U545 ( .A(n1154), .Y(n1155) );
  clknd2d1_hd U546 ( .A(n476), .B(n1422), .Y(n1427) );
  nid1_hd U547 ( .A(n1149), .Y(n1150) );
  clknd2d1_hd U548 ( .A(n477), .B(n1380), .Y(n1400) );
  nid1_hd U549 ( .A(n1484), .Y(n1156) );
  nid1_hd U550 ( .A(n1483), .Y(n1149) );
  clknd2d1_hd U551 ( .A(n407), .B(n1400), .Y(n1403) );
  clknd2d1_hd U552 ( .A(N34), .B(n158), .Y(n157) );
  clknd2d1_hd U553 ( .A(n518), .B(a_e[0]), .Y(n1189) );
  clknd2d1_hd U554 ( .A(n575), .B(b_e[0]), .Y(n1173) );
  nid1_hd U555 ( .A(n1153), .Y(n1151) );
  nid1_hd U556 ( .A(b_m[4]), .Y(n1042) );
  nid1_hd U557 ( .A(n1139), .Y(n1132) );
  nid1_hd U558 ( .A(b_m[6]), .Y(n1032) );
  nid1_hd U559 ( .A(b_m[5]), .Y(n1037) );
  nid1_hd U560 ( .A(b_m[10]), .Y(n1009) );
  nid1_hd U561 ( .A(b_m[19]), .Y(n967) );
  clknd2d1_hd U562 ( .A(n1278), .B(n1277), .Y(n1283) );
  clknd2d1_hd U563 ( .A(n1263), .B(n1262), .Y(n1266) );
  clknd2d1_hd U564 ( .A(n1270), .B(n1269), .Y(n1273) );
  clknd2d1_hd U565 ( .A(n1293), .B(n1257), .Y(n1252) );
  nid1_hd U566 ( .A(n1327), .Y(n1142) );
  nid1_hd U567 ( .A(n1139), .Y(n1134) );
  nid1_hd U568 ( .A(n1327), .Y(n1141) );
  nid1_hd U569 ( .A(n1139), .Y(n1133) );
  nid1_hd U570 ( .A(n1327), .Y(n1143) );
  nid1_hd U571 ( .A(b_m[3]), .Y(n1047) );
  nid1_hd U572 ( .A(n1132), .Y(n1136) );
  nid1_hd U573 ( .A(b_m[9]), .Y(n1014) );
  nid1_hd U574 ( .A(n1361), .Y(n1146) );
  nid1_hd U575 ( .A(b_m[11]), .Y(n1004) );
  nid1_hd U576 ( .A(b_m[12]), .Y(n999) );
  nid1_hd U577 ( .A(b_m[13]), .Y(n994) );
  nid1_hd U578 ( .A(n1139), .Y(n1137) );
  nid1_hd U579 ( .A(n1361), .Y(n1147) );
  nid1_hd U580 ( .A(b_m[15]), .Y(n987) );
  nid1_hd U581 ( .A(b_m[16]), .Y(n982) );
  nid1_hd U582 ( .A(b_m[17]), .Y(n977) );
  nid1_hd U583 ( .A(b_m[18]), .Y(n972) );
  nid1_hd U584 ( .A(n1361), .Y(n1148) );
  nid1_hd U585 ( .A(n1139), .Y(n1138) );
  nid1_hd U586 ( .A(b_m[2]), .Y(n1052) );
  nid1_hd U587 ( .A(n957), .Y(n953) );
  nid1_hd U588 ( .A(n1132), .Y(n1135) );
  clknd2d1_hd U589 ( .A(state[1]), .B(n1218), .Y(n1398) );
  clknd2d1_hd U590 ( .A(n1151), .B(n1394), .Y(n1395) );
  nid1_hd U591 ( .A(n1215), .Y(n1139) );
  nid1_hd U592 ( .A(n1327), .Y(n1144) );
  nid1_hd U593 ( .A(n1361), .Y(n1145) );
  clknd2d1_hd U594 ( .A(n1181), .B(n1180), .Y(n1185) );
  clknd2d1_hd U595 ( .A(n1193), .B(n1192), .Y(n1195) );
  clknd2d1_hd U596 ( .A(n947), .B(n956), .Y(n860) );
  fad1_hd U597 ( .A(mult_x_1_n190), .B(mult_x_1_n187), .CI(mult_x_1_n135), 
        .CO(mult_x_1_n134), .S(N220) );
  fad1_hd U598 ( .A(mult_x_1_n195), .B(mult_x_1_n191), .CI(mult_x_1_n136), 
        .CO(mult_x_1_n135), .S(N219) );
  fad1_hd U599 ( .A(mult_x_1_n196), .B(mult_x_1_n200), .CI(mult_x_1_n137), 
        .CO(mult_x_1_n136), .S(N218) );
  nid1_hd U600 ( .A(DP_OP_125J2_130_6300_I3), .Y(n580) );
  fad1_hd U601 ( .A(mult_x_1_n206), .B(mult_x_1_n201), .CI(mult_x_1_n138), 
        .CO(mult_x_1_n137), .S(N217) );
  fad1_hd U602 ( .A(mult_x_1_n213), .B(mult_x_1_n207), .CI(mult_x_1_n139), 
        .CO(mult_x_1_n138), .S(N216) );
  fad1_hd U603 ( .A(mult_x_1_n214), .B(mult_x_1_n220), .CI(mult_x_1_n140), 
        .CO(mult_x_1_n139), .S(N215) );
  fad1_hd U604 ( .A(mult_x_1_n238), .B(mult_x_1_n246), .CI(mult_x_1_n143), 
        .CO(mult_x_1_n142), .S(N212) );
  fad1_hd U605 ( .A(mult_x_1_n256), .B(mult_x_1_n247), .CI(mult_x_1_n144), 
        .CO(mult_x_1_n143), .S(N211) );
  fad1_hd U606 ( .A(mult_x_1_n267), .B(mult_x_1_n257), .CI(mult_x_1_n145), 
        .CO(mult_x_1_n144), .S(N210) );
  fad1_hd U607 ( .A(mult_x_1_n268), .B(mult_x_1_n278), .CI(mult_x_1_n146), 
        .CO(mult_x_1_n145), .S(N209) );
  fad1_hd U608 ( .A(mult_x_1_n290), .B(mult_x_1_n279), .CI(mult_x_1_n147), 
        .CO(mult_x_1_n146), .S(N208) );
  fad1_hd U609 ( .A(mult_x_1_n303), .B(mult_x_1_n291), .CI(mult_x_1_n148), 
        .CO(mult_x_1_n147), .S(N207) );
  fad1_hd U610 ( .A(mult_x_1_n304), .B(mult_x_1_n316), .CI(mult_x_1_n149), 
        .CO(mult_x_1_n148), .S(N206) );
  nid1_hd U611 ( .A(n1128), .Y(n1127) );
  clknd2d1_hd U612 ( .A(n951), .B(n1121), .Y(n829) );
  nid1_hd U613 ( .A(n1129), .Y(DP_OP_125J2_130_6300_I3) );
  nid1_hd U614 ( .A(n1214), .Y(n1129) );
  nid1_hd U615 ( .A(n1214), .Y(n1128) );
  clknd2d1_hd U616 ( .A(n1393), .B(n1378), .Y(n105) );
  nid1_hd U617 ( .A(n146), .Y(n368) );
  nid1_hd U618 ( .A(n372), .Y(n1166) );
  nid1_hd U619 ( .A(n1166), .Y(n1169) );
  nid1_hd U620 ( .A(n384), .Y(n385) );
  nid1_hd U621 ( .A(n1168), .Y(n1167) );
  nid1_hd U622 ( .A(n1214), .Y(n383) );
  nid1_hd U623 ( .A(n1169), .Y(n1168) );
  nid1_hd U624 ( .A(n146), .Y(n372) );
  nid1_hd U625 ( .A(n146), .Y(n374) );
  nid1_hd U626 ( .A(n146), .Y(n373) );
  nid1_hd U627 ( .A(n371), .Y(n386) );
  clknd2d1_hd U628 ( .A(n1202), .B(a_e[8]), .Y(n1196) );
  clknd2d1_hd U629 ( .A(n1186), .B(b_e[8]), .Y(n1187) );
  clknd2d1_hd U630 ( .A(n1404), .B(n474), .Y(n1405) );
  clknd2d1_hd U631 ( .A(n472), .B(n1402), .Y(n1401) );
  clknd2d1_hd U632 ( .A(n1202), .B(a_e[1]), .Y(n1191) );
  clknd2d1_hd U633 ( .A(n1186), .B(b_e[1]), .Y(n1179) );
  clknd2d1_hd U634 ( .A(n1163), .B(n1286), .Y(n1287) );
  clknd2d1_hd U635 ( .A(z_e[7]), .B(n1283), .Y(n1281) );
  clknd2d1_hd U636 ( .A(n1285), .B(n1265), .Y(n235) );
  clknd2d1_hd U637 ( .A(n1285), .B(n1272), .Y(n233) );
  clknd2d1_hd U638 ( .A(n1162), .B(z[23]), .Y(n1259) );
  clknd2d1_hd U639 ( .A(n1162), .B(z[24]), .Y(n1260) );
  clknd2d1_hd U640 ( .A(n1285), .B(n1280), .Y(n231) );
  clknd2d1_hd U641 ( .A(n1162), .B(z[26]), .Y(n1267) );
  clknd2d1_hd U642 ( .A(n1162), .B(z[28]), .Y(n1274) );
  clknd2d1_hd U643 ( .A(a_m[22]), .B(n519), .Y(n1299) );
  clknd2d1_hd U644 ( .A(n1300), .B(a_m[23]), .Y(n1298) );
  clknd2d1_hd U645 ( .A(n575), .B(n488), .Y(n1337) );
  clknd2d1_hd U646 ( .A(n1339), .B(b_m[23]), .Y(n1336) );
  clknd2d1_hd U647 ( .A(n1186), .B(b_e[9]), .Y(n1176) );
  clknd2d1_hd U648 ( .A(n574), .B(b_e[9]), .Y(n1175) );
  clknd2d1_hd U649 ( .A(n1202), .B(a_e[9]), .Y(n1203) );
  clknd2d1_hd U650 ( .A(n517), .B(a_e[9]), .Y(n1201) );
  clknd2d1_hd U651 ( .A(n1330), .B(n1297), .Y(n148) );
  clknd2d1_hd U652 ( .A(n1330), .B(n1331), .Y(n138) );
  fad1_hd U653 ( .A(n1003), .B(n998), .CI(mult_x_1_n627), .CO(mult_x_1_n626), 
        .S(mult_x_1_n651) );
  fad1_hd U654 ( .A(n1008), .B(n1003), .CI(mult_x_1_n628), .CO(mult_x_1_n627), 
        .S(mult_x_1_n652) );
  fad1_hd U655 ( .A(n1013), .B(n1008), .CI(mult_x_1_n629), .CO(mult_x_1_n628), 
        .S(mult_x_1_n653) );
  fad1_hd U656 ( .A(n1018), .B(n1013), .CI(mult_x_1_n630), .CO(mult_x_1_n629), 
        .S(mult_x_1_n654) );
  fad1_hd U657 ( .A(n1022), .B(n1018), .CI(mult_x_1_n631), .CO(mult_x_1_n630), 
        .S(mult_x_1_n655) );
  fad1_hd U658 ( .A(n1026), .B(n1022), .CI(mult_x_1_n632), .CO(mult_x_1_n631), 
        .S(mult_x_1_n656) );
  had1_hd U659 ( .A(n952), .B(mult_x_1_n616), .CO(mult_x_1_n639), .S(
        mult_x_1_n640) );
  fad1_hd U660 ( .A(n998), .B(n991), .CI(mult_x_1_n626), .CO(mult_x_1_n625), 
        .S(mult_x_1_n650) );
  ivd1_hd U661 ( .A(a_m[23]), .Y(n886) );
  ivd1_hd U662 ( .A(n359), .Y(n369) );
  ivd1_hd U663 ( .A(n359), .Y(n370) );
  nid1_hd U664 ( .A(n146), .Y(n371) );
  scg12d1_hd U665 ( .A(o_AB_ACK), .B(i_AB_STB), .C(n155), .Y(n146) );
  ivd1_hd U666 ( .A(n381), .Y(n382) );
  ivd1_hd U667 ( .A(n382), .Y(n375) );
  ivd1_hd U668 ( .A(n382), .Y(n376) );
  ivd1_hd U669 ( .A(n382), .Y(n377) );
  or3d1_hd U670 ( .A(n1220), .B(n34), .C(n1289), .Y(n359) );
  ivd1_hd U671 ( .A(n359), .Y(n378) );
  ivd1_hd U672 ( .A(n359), .Y(n379) );
  ivd1_hd U673 ( .A(n359), .Y(n380) );
  nr3d1_hd U674 ( .A(n1291), .B(n463), .C(n1221), .Y(n381) );
  nid1_hd U675 ( .A(n146), .Y(n384) );
  nid1_hd U676 ( .A(b_m[6]), .Y(n1033) );
  ivd1_hd U677 ( .A(a_m[20]), .Y(n897) );
  ivd1_hd U678 ( .A(mult_x_1_n640), .Y(n452) );
  ivd1_hd U679 ( .A(mult_x_1_n641), .Y(n408) );
  ivd1_hd U680 ( .A(mult_x_1_n642), .Y(n448) );
  nid1_hd U681 ( .A(b_m[14]), .Y(n993) );
  xo3d1_hd U682 ( .A(mult_x_1_n180), .B(mult_x_1_n132), .C(n861), .Y(N223) );
  ivd1_hd U683 ( .A(n452), .Y(n453) );
  ivd1_hd U684 ( .A(n408), .Y(n409) );
  ivd1_hd U685 ( .A(n448), .Y(n449) );
  fad1_hd U686 ( .A(n487), .B(n952), .CI(mult_x_1_n617), .CO(mult_x_1_n616), 
        .S(mult_x_1_n641) );
  ivd1_hd U687 ( .A(n446), .Y(n447) );
  ivd1_hd U688 ( .A(mult_x_1_n643), .Y(n450) );
  ivd1_hd U689 ( .A(mult_x_1_n644), .Y(n446) );
  ivd1_hd U690 ( .A(mult_x_1_n645), .Y(n444) );
  ivd1_hd U691 ( .A(mult_x_1_n646), .Y(n442) );
  ivd1_hd U692 ( .A(mult_x_1_n647), .Y(n440) );
  nid1_hd U693 ( .A(n821), .Y(n1108) );
  nid1_hd U694 ( .A(n925), .Y(n926) );
  nid1_hd U695 ( .A(n886), .Y(n888) );
  nid1_hd U696 ( .A(n946), .Y(n947) );
  ivd1_hd U697 ( .A(a_m[8]), .Y(n925) );
  ivd1_hd U698 ( .A(a_m[17]), .Y(n904) );
  ivd1_hd U699 ( .A(a_m[14]), .Y(n911) );
  xo2d1_hd U700 ( .A(n944), .B(n830), .Y(mult_x_1_n855) );
  xo2d1_hd U701 ( .A(n930), .B(n762), .Y(mult_x_1_n801) );
  xo2d1_hd U702 ( .A(n916), .B(n692), .Y(mult_x_1_n747) );
  xo2d1_hd U703 ( .A(n923), .B(n727), .Y(mult_x_1_n774) );
  xo2d1_hd U704 ( .A(n937), .B(n797), .Y(mult_x_1_n828) );
  xo2d1_hd U705 ( .A(n906), .B(n659), .Y(mult_x_1_n721) );
  xo2d1_hd U706 ( .A(n920), .B(n729), .Y(mult_x_1_n775) );
  xo2d1_hd U707 ( .A(n913), .B(n694), .Y(mult_x_1_n748) );
  xo2d1_hd U708 ( .A(n934), .B(n799), .Y(mult_x_1_n829) );
  xo2d1_hd U709 ( .A(a_m[2]), .B(n832), .Y(mult_x_1_n856) );
  xo2d1_hd U710 ( .A(n927), .B(n764), .Y(mult_x_1_n802) );
  xo2d1_hd U711 ( .A(n906), .B(n660), .Y(mult_x_1_n722) );
  xo2d1_hd U712 ( .A(n941), .B(n833), .Y(mult_x_1_n857) );
  xo2d1_hd U713 ( .A(n913), .B(n695), .Y(mult_x_1_n749) );
  xo2d1_hd U714 ( .A(n934), .B(n800), .Y(mult_x_1_n830) );
  xo2d1_hd U715 ( .A(n920), .B(n730), .Y(mult_x_1_n776) );
  xo2d1_hd U716 ( .A(n927), .B(n765), .Y(mult_x_1_n803) );
  xo2d1_hd U717 ( .A(n899), .B(n625), .Y(mult_x_1_n695) );
  nid1_hd U718 ( .A(mult_x_1_n639), .Y(n525) );
  xo2d1_hd U719 ( .A(n927), .B(n766), .Y(mult_x_1_n804) );
  xo2d1_hd U720 ( .A(n934), .B(n801), .Y(mult_x_1_n831) );
  xo2d1_hd U721 ( .A(n920), .B(n731), .Y(mult_x_1_n777) );
  xo2d1_hd U722 ( .A(n899), .B(n627), .Y(mult_x_1_n697) );
  xo2d1_hd U723 ( .A(n906), .B(n662), .Y(mult_x_1_n724) );
  xo2d1_hd U724 ( .A(n920), .B(n732), .Y(mult_x_1_n778) );
  xo2d1_hd U725 ( .A(n913), .B(n697), .Y(mult_x_1_n751) );
  xo2d1_hd U726 ( .A(n927), .B(n767), .Y(mult_x_1_n805) );
  xo2d1_hd U727 ( .A(n934), .B(n802), .Y(mult_x_1_n832) );
  ivd1_hd U728 ( .A(n450), .Y(n451) );
  xo2d1_hd U729 ( .A(n928), .B(n768), .Y(mult_x_1_n806) );
  xo2d1_hd U730 ( .A(n928), .B(n769), .Y(mult_x_1_n807) );
  xo2d1_hd U731 ( .A(n921), .B(n734), .Y(mult_x_1_n780) );
  xo2d1_hd U732 ( .A(n928), .B(n770), .Y(mult_x_1_n808) );
  ivd1_hd U733 ( .A(n444), .Y(n445) );
  xo2d1_hd U734 ( .A(n921), .B(n735), .Y(mult_x_1_n781) );
  xo2d1_hd U735 ( .A(n921), .B(n736), .Y(mult_x_1_n782) );
  ivd1_hd U736 ( .A(n442), .Y(n443) );
  xo2d1_hd U737 ( .A(n921), .B(n737), .Y(mult_x_1_n783) );
  ivd1_hd U738 ( .A(mult_x_1_n648), .Y(n436) );
  xo2d1_hd U739 ( .A(n915), .B(n704), .Y(mult_x_1_n758) );
  xo2d1_hd U740 ( .A(n922), .B(n739), .Y(mult_x_1_n785) );
  xo2d1_hd U741 ( .A(n922), .B(n740), .Y(mult_x_1_n786) );
  ivd1_hd U742 ( .A(mult_x_1_n649), .Y(n438) );
  xo2d1_hd U743 ( .A(n922), .B(n741), .Y(mult_x_1_n787) );
  or2d1_hd U744 ( .A(n658), .B(n685), .Y(n682) );
  nd3d1_hd U745 ( .A(n588), .B(n615), .C(n583), .Y(n586) );
  nid1_hd U746 ( .A(n823), .Y(n1113) );
  or2d1_hd U747 ( .A(n588), .B(n615), .Y(n613) );
  nd3d1_hd U748 ( .A(n658), .B(n685), .C(n653), .Y(n656) );
  nd3d1_hd U749 ( .A(n693), .B(n720), .C(n688), .Y(n691) );
  or2d1_hd U750 ( .A(n693), .B(n720), .Y(n717) );
  nr2bd1_hd U751 ( .AN(n693), .B(n720), .Y(n718) );
  nd3d1_hd U752 ( .A(n623), .B(n650), .C(n618), .Y(n621) );
  xo2d1_hd U753 ( .A(n944), .B(n859), .Y(mult_x_1_n879) );
  nd3d1_hd U754 ( .A(n728), .B(n755), .C(n723), .Y(n726) );
  or2d1_hd U755 ( .A(n728), .B(n755), .Y(n752) );
  nd3d1_hd U756 ( .A(n763), .B(n790), .C(n758), .Y(n761) );
  or2d1_hd U757 ( .A(n623), .B(n650), .Y(n647) );
  nid1_hd U758 ( .A(n853), .Y(n1118) );
  nd3d1_hd U759 ( .A(n798), .B(n825), .C(n793), .Y(n796) );
  nid1_hd U760 ( .A(n932), .Y(n933) );
  ivd1_hd U761 ( .A(a_m[11]), .Y(n918) );
  nid1_hd U762 ( .A(b_m[3]), .Y(n1048) );
  nid1_hd U763 ( .A(b_m[0]), .Y(n579) );
  ivd1_hd U764 ( .A(a_m[5]), .Y(n932) );
  ivd1_hd U765 ( .A(b_m[22]), .Y(n485) );
  xo2d1_hd U766 ( .A(n909), .B(n657), .Y(mult_x_1_n720) );
  xo2d1_hd U767 ( .A(n902), .B(n622), .Y(mult_x_1_n693) );
  xo2d1_hd U768 ( .A(n892), .B(n587), .Y(mult_x_1_n666) );
  xo2d1_hd U769 ( .A(n899), .B(n624), .Y(mult_x_1_n694) );
  xo2d1_hd U770 ( .A(n617), .B(n897), .Y(mult_x_1_n692) );
  xo2d1_hd U771 ( .A(n652), .B(n904), .Y(mult_x_1_n719) );
  xo2d1_hd U772 ( .A(n892), .B(n589), .Y(mult_x_1_n667) );
  xo2d1_hd U773 ( .A(n582), .B(n886), .Y(mult_x_1_n665) );
  xo2d1_hd U774 ( .A(n827), .B(n939), .Y(mult_x_1_n854) );
  xo2d1_hd U775 ( .A(n687), .B(n911), .Y(mult_x_1_n746) );
  xo2d1_hd U776 ( .A(n722), .B(n918), .Y(mult_x_1_n773) );
  xo2d1_hd U777 ( .A(n757), .B(n926), .Y(mult_x_1_n800) );
  xo2d1_hd U778 ( .A(n792), .B(n932), .Y(mult_x_1_n827) );
  xo2d1_hd U779 ( .A(n892), .B(n590), .Y(mult_x_1_n668) );
  xo2d1_hd U780 ( .A(n893), .B(n591), .Y(mult_x_1_n669) );
  xo2d1_hd U781 ( .A(n913), .B(n696), .Y(mult_x_1_n750) );
  xo2d1_hd U782 ( .A(n899), .B(n626), .Y(mult_x_1_n696) );
  xo2d1_hd U783 ( .A(n906), .B(n661), .Y(mult_x_1_n723) );
  xo2d1_hd U784 ( .A(n941), .B(n834), .Y(mult_x_1_n858) );
  xo2d1_hd U785 ( .A(n943), .B(n835), .Y(mult_x_1_n859) );
  xo2d1_hd U786 ( .A(n893), .B(n592), .Y(mult_x_1_n670) );
  xo2d1_hd U787 ( .A(n900), .B(n628), .Y(mult_x_1_n698) );
  xo2d1_hd U788 ( .A(n914), .B(n698), .Y(mult_x_1_n752) );
  xo2d1_hd U789 ( .A(n907), .B(n663), .Y(mult_x_1_n725) );
  xo2d1_hd U790 ( .A(n921), .B(n733), .Y(mult_x_1_n779) );
  xo2d1_hd U791 ( .A(n935), .B(n803), .Y(mult_x_1_n833) );
  xo2d1_hd U792 ( .A(n893), .B(n593), .Y(mult_x_1_n671) );
  xo2d1_hd U793 ( .A(n941), .B(n836), .Y(mult_x_1_n860) );
  xo2d1_hd U794 ( .A(n900), .B(n629), .Y(mult_x_1_n699) );
  xo2d1_hd U795 ( .A(n941), .B(n837), .Y(mult_x_1_n861) );
  xo2d1_hd U796 ( .A(n935), .B(n804), .Y(mult_x_1_n834) );
  xo2d1_hd U797 ( .A(n893), .B(n594), .Y(mult_x_1_n672) );
  xo2d1_hd U798 ( .A(n914), .B(n699), .Y(mult_x_1_n753) );
  xo2d1_hd U799 ( .A(n907), .B(n664), .Y(mult_x_1_n726) );
  xo2d1_hd U800 ( .A(n893), .B(n595), .Y(mult_x_1_n673) );
  xo2d1_hd U801 ( .A(n900), .B(n630), .Y(mult_x_1_n700) );
  xo2d1_hd U802 ( .A(n941), .B(n838), .Y(mult_x_1_n862) );
  xo2d1_hd U803 ( .A(n914), .B(n700), .Y(mult_x_1_n754) );
  xo2d1_hd U804 ( .A(n907), .B(n665), .Y(mult_x_1_n727) );
  xo2d1_hd U805 ( .A(n935), .B(n805), .Y(mult_x_1_n835) );
  xo2d1_hd U806 ( .A(n941), .B(n839), .Y(mult_x_1_n863) );
  xo2d1_hd U807 ( .A(n935), .B(n806), .Y(mult_x_1_n836) );
  xo2d1_hd U808 ( .A(n928), .B(n771), .Y(mult_x_1_n809) );
  xo2d1_hd U809 ( .A(n907), .B(n666), .Y(mult_x_1_n728) );
  xo2d1_hd U810 ( .A(n914), .B(n701), .Y(mult_x_1_n755) );
  xo2d1_hd U811 ( .A(n900), .B(n631), .Y(mult_x_1_n701) );
  xo2d1_hd U812 ( .A(n894), .B(n596), .Y(mult_x_1_n674) );
  xo2d1_hd U813 ( .A(n907), .B(n667), .Y(mult_x_1_n729) );
  xo2d1_hd U814 ( .A(n914), .B(n702), .Y(mult_x_1_n756) );
  xo2d1_hd U815 ( .A(n928), .B(n772), .Y(mult_x_1_n810) );
  xo2d1_hd U816 ( .A(n900), .B(n632), .Y(mult_x_1_n702) );
  xo2d1_hd U817 ( .A(n894), .B(n597), .Y(mult_x_1_n675) );
  xo2d1_hd U818 ( .A(n942), .B(n840), .Y(mult_x_1_n864) );
  xo2d1_hd U819 ( .A(n935), .B(n807), .Y(mult_x_1_n837) );
  xo2d1_hd U820 ( .A(n894), .B(n598), .Y(mult_x_1_n676) );
  xo2d1_hd U821 ( .A(n935), .B(n808), .Y(mult_x_1_n838) );
  xo2d1_hd U822 ( .A(n921), .B(n738), .Y(mult_x_1_n784) );
  xo2d1_hd U823 ( .A(n914), .B(n703), .Y(mult_x_1_n757) );
  xo2d1_hd U824 ( .A(n942), .B(n841), .Y(mult_x_1_n865) );
  xo2d1_hd U825 ( .A(n928), .B(n773), .Y(mult_x_1_n811) );
  xo2d1_hd U826 ( .A(n900), .B(n633), .Y(mult_x_1_n703) );
  xo2d1_hd U827 ( .A(n907), .B(n668), .Y(mult_x_1_n730) );
  xo2d1_hd U828 ( .A(n929), .B(n774), .Y(mult_x_1_n812) );
  xo2d1_hd U829 ( .A(n1175), .B(n1184), .Y(n1177) );
  xo2d1_hd U830 ( .A(n1201), .B(n1200), .Y(n1204) );
  xo2d1_hd U831 ( .A(n893), .B(n599), .Y(mult_x_1_n677) );
  xo2d1_hd U832 ( .A(n901), .B(n634), .Y(mult_x_1_n704) );
  xo2d1_hd U833 ( .A(n936), .B(n809), .Y(mult_x_1_n839) );
  xo2d1_hd U834 ( .A(n908), .B(n669), .Y(mult_x_1_n731) );
  xo2d1_hd U835 ( .A(n942), .B(n842), .Y(mult_x_1_n866) );
  xo2d1_hd U836 ( .A(n929), .B(n775), .Y(mult_x_1_n813) );
  xo2d1_hd U837 ( .A(n894), .B(n600), .Y(mult_x_1_n678) );
  xo2d1_hd U838 ( .A(n908), .B(n670), .Y(mult_x_1_n732) );
  xo2d1_hd U839 ( .A(n915), .B(n705), .Y(mult_x_1_n759) );
  xo2d1_hd U840 ( .A(n936), .B(n810), .Y(mult_x_1_n840) );
  xo2d1_hd U841 ( .A(n901), .B(n635), .Y(mult_x_1_n705) );
  xo2d1_hd U842 ( .A(n942), .B(n843), .Y(mult_x_1_n867) );
  xo2d1_hd U843 ( .A(n936), .B(n811), .Y(mult_x_1_n841) );
  xo2d1_hd U844 ( .A(n915), .B(n706), .Y(mult_x_1_n760) );
  xo2d1_hd U845 ( .A(n901), .B(n636), .Y(mult_x_1_n706) );
  xo2d1_hd U846 ( .A(n894), .B(n601), .Y(mult_x_1_n679) );
  xo2d1_hd U847 ( .A(n929), .B(n776), .Y(mult_x_1_n814) );
  xo2d1_hd U848 ( .A(n908), .B(n671), .Y(mult_x_1_n733) );
  xo2d1_hd U849 ( .A(n942), .B(n844), .Y(mult_x_1_n868) );
  xo2d1_hd U850 ( .A(n908), .B(n672), .Y(mult_x_1_n734) );
  xo2d1_hd U851 ( .A(n915), .B(n707), .Y(mult_x_1_n761) );
  xo2d1_hd U852 ( .A(n942), .B(n845), .Y(mult_x_1_n869) );
  xo2d1_hd U853 ( .A(n936), .B(n812), .Y(mult_x_1_n842) );
  xo2d1_hd U854 ( .A(n922), .B(n742), .Y(mult_x_1_n788) );
  xo2d1_hd U855 ( .A(n901), .B(n637), .Y(mult_x_1_n707) );
  xo2d1_hd U856 ( .A(n929), .B(n777), .Y(mult_x_1_n815) );
  xo2d1_hd U857 ( .A(n895), .B(n602), .Y(mult_x_1_n680) );
  xo2d1_hd U858 ( .A(n943), .B(n846), .Y(mult_x_1_n870) );
  xo2d1_hd U859 ( .A(n915), .B(n708), .Y(mult_x_1_n762) );
  xo2d1_hd U860 ( .A(n929), .B(n778), .Y(mult_x_1_n816) );
  xo2d1_hd U861 ( .A(n922), .B(n743), .Y(mult_x_1_n789) );
  xo2d1_hd U862 ( .A(n895), .B(n603), .Y(mult_x_1_n681) );
  xo2d1_hd U863 ( .A(n936), .B(n813), .Y(mult_x_1_n843) );
  xo2d1_hd U864 ( .A(n908), .B(n673), .Y(mult_x_1_n735) );
  xo2d1_hd U865 ( .A(n901), .B(n638), .Y(mult_x_1_n708) );
  xo2d1_hd U866 ( .A(n902), .B(n639), .Y(mult_x_1_n709) );
  xo2d1_hd U867 ( .A(n937), .B(n814), .Y(mult_x_1_n844) );
  xo2d1_hd U868 ( .A(n943), .B(n847), .Y(mult_x_1_n871) );
  xo2d1_hd U869 ( .A(n916), .B(n709), .Y(mult_x_1_n763) );
  xo2d1_hd U870 ( .A(n923), .B(n744), .Y(mult_x_1_n790) );
  xo2d1_hd U871 ( .A(n909), .B(n674), .Y(mult_x_1_n736) );
  xo2d1_hd U872 ( .A(n895), .B(n604), .Y(mult_x_1_n682) );
  xo2d1_hd U873 ( .A(n930), .B(n779), .Y(mult_x_1_n817) );
  xo2d1_hd U874 ( .A(n923), .B(n745), .Y(mult_x_1_n791) );
  xo2d1_hd U875 ( .A(n902), .B(n640), .Y(mult_x_1_n710) );
  xo2d1_hd U876 ( .A(n895), .B(n605), .Y(mult_x_1_n683) );
  xo2d1_hd U877 ( .A(n930), .B(n780), .Y(mult_x_1_n818) );
  xo2d1_hd U878 ( .A(n937), .B(n815), .Y(mult_x_1_n845) );
  xo2d1_hd U879 ( .A(n943), .B(n848), .Y(mult_x_1_n872) );
  xo2d1_hd U880 ( .A(n909), .B(n675), .Y(mult_x_1_n737) );
  xo2d1_hd U881 ( .A(n916), .B(n710), .Y(mult_x_1_n764) );
  xo2d1_hd U882 ( .A(n916), .B(n711), .Y(mult_x_1_n765) );
  xo2d1_hd U883 ( .A(n909), .B(n676), .Y(mult_x_1_n738) );
  xo2d1_hd U884 ( .A(n937), .B(n816), .Y(mult_x_1_n846) );
  xo2d1_hd U885 ( .A(n923), .B(n746), .Y(mult_x_1_n792) );
  xo2d1_hd U886 ( .A(n902), .B(n641), .Y(mult_x_1_n711) );
  xo2d1_hd U887 ( .A(n895), .B(n606), .Y(mult_x_1_n684) );
  xo2d1_hd U888 ( .A(n930), .B(n781), .Y(mult_x_1_n819) );
  xo2d1_hd U889 ( .A(n943), .B(n849), .Y(mult_x_1_n873) );
  or2d1_hd U890 ( .A(n460), .B(n1368), .Y(n1468) );
  xo2d1_hd U891 ( .A(n895), .B(n607), .Y(mult_x_1_n685) );
  xo2d1_hd U892 ( .A(n943), .B(n850), .Y(mult_x_1_n874) );
  xo2d1_hd U893 ( .A(n901), .B(n642), .Y(mult_x_1_n712) );
  xo2d1_hd U894 ( .A(n936), .B(n817), .Y(mult_x_1_n847) );
  xo2d1_hd U895 ( .A(n908), .B(n677), .Y(mult_x_1_n739) );
  xo2d1_hd U896 ( .A(n922), .B(n747), .Y(mult_x_1_n793) );
  xo2d1_hd U897 ( .A(n929), .B(n782), .Y(mult_x_1_n820) );
  xo2d1_hd U898 ( .A(n915), .B(n712), .Y(mult_x_1_n766) );
  xo2d1_hd U899 ( .A(n902), .B(n643), .Y(mult_x_1_n713) );
  xo2d1_hd U900 ( .A(n944), .B(n851), .Y(mult_x_1_n875) );
  xo2d1_hd U901 ( .A(n923), .B(n748), .Y(mult_x_1_n794) );
  xo2d1_hd U902 ( .A(n896), .B(n608), .Y(mult_x_1_n686) );
  xo2d1_hd U903 ( .A(n930), .B(n783), .Y(mult_x_1_n821) );
  xo2d1_hd U904 ( .A(n937), .B(n818), .Y(mult_x_1_n848) );
  xo2d1_hd U905 ( .A(n916), .B(n713), .Y(mult_x_1_n767) );
  xo2d1_hd U906 ( .A(n909), .B(n678), .Y(mult_x_1_n740) );
  xo2d1_hd U907 ( .A(n916), .B(n714), .Y(mult_x_1_n768) );
  xo2d1_hd U908 ( .A(n909), .B(n679), .Y(mult_x_1_n741) );
  xo2d1_hd U909 ( .A(n894), .B(n609), .Y(mult_x_1_n687) );
  xo2d1_hd U910 ( .A(n944), .B(n852), .Y(mult_x_1_n876) );
  xo2d1_hd U911 ( .A(n930), .B(n784), .Y(mult_x_1_n822) );
  xo2d1_hd U912 ( .A(n937), .B(n819), .Y(mult_x_1_n849) );
  xo2d1_hd U913 ( .A(n902), .B(n644), .Y(mult_x_1_n714) );
  xo2d1_hd U914 ( .A(n923), .B(n749), .Y(mult_x_1_n795) );
  xo2d1_hd U915 ( .A(n944), .B(n854), .Y(mult_x_1_n877) );
  xo2d1_hd U916 ( .A(n896), .B(n610), .Y(mult_x_1_n688) );
  xo2d1_hd U917 ( .A(n896), .B(n614), .Y(mult_x_1_n689) );
  xo2d1_hd U918 ( .A(n924), .B(n754), .Y(mult_x_1_n797) );
  xo2d1_hd U919 ( .A(n903), .B(n649), .Y(mult_x_1_n716) );
  xo2d1_hd U920 ( .A(n944), .B(n858), .Y(mult_x_1_n878) );
  xo2d1_hd U921 ( .A(n931), .B(n789), .Y(mult_x_1_n824) );
  nid1_hd U922 ( .A(n751), .Y(n1094) );
  nid1_hd U923 ( .A(n788), .Y(n1103) );
  nid1_hd U924 ( .A(n1124), .Y(n1125) );
  ad2d1_hd U925 ( .A(n1171), .B(n1170), .Y(n1332) );
  nid1_hd U926 ( .A(n857), .Y(n1124) );
  nid1_hd U927 ( .A(n786), .Y(n1102) );
  nid1_hd U928 ( .A(n821), .Y(n1107) );
  nid1_hd U929 ( .A(n855), .Y(n1122) );
  xo2d1_hd U930 ( .A(a_s), .B(b_s), .Y(N35) );
  ivd1_hd U931 ( .A(b_m[23]), .Y(n946) );
  or2d1_hd U932 ( .A(n1415), .B(n528), .Y(n1419) );
  or2d1_hd U933 ( .A(n1430), .B(n530), .Y(n1434) );
  or2d1_hd U934 ( .A(n1445), .B(n528), .Y(n1449) );
  or2d1_hd U935 ( .A(n1461), .B(n529), .Y(n1465) );
  ad2d1_hd U936 ( .A(n571), .B(n407), .Y(n1472) );
  ad2d1_hd U937 ( .A(n1379), .B(n1378), .Y(n110) );
  nid1_hd U938 ( .A(n1484), .Y(n1154) );
  scg10d1_hd U939 ( .A(n1288), .B(n1287), .C(z[31]), .D(n1164), .Y(n229) );
  nid1_hd U940 ( .A(n1484), .Y(n1157) );
  scg2d1_hd U941 ( .A(n1131), .B(a[26]), .C(n517), .D(a_e[3]), .Y(C1_Z_3) );
  scg2d1_hd U942 ( .A(n1132), .B(a[25]), .C(n519), .D(a_e[2]), .Y(C1_Z_2) );
  scg2d1_hd U943 ( .A(n1139), .B(a[0]), .C(a_m[0]), .D(n1144), .Y(n349) );
  scg2d1_hd U944 ( .A(n1132), .B(a[27]), .C(n518), .D(a_e[4]), .Y(C1_Z_4) );
  or2d1_hd U945 ( .A(n1217), .B(n1148), .Y(n1363) );
  scg2d1_hd U946 ( .A(n1131), .B(a[28]), .C(n517), .D(a_e[5]), .Y(C1_Z_5) );
  or2d1_hd U947 ( .A(n1377), .B(n105), .Y(n1460) );
  scg2d1_hd U948 ( .A(n1140), .B(b[0]), .C(n1145), .D(b_m[0]), .Y(n308) );
  scg2d1_hd U949 ( .A(n1131), .B(a[24]), .C(n517), .D(a_e[1]), .Y(C1_Z_1) );
  scg2d1_hd U950 ( .A(n1131), .B(a[29]), .C(n518), .D(a_e[6]), .Y(C1_Z_6) );
  scg2d1_hd U951 ( .A(n1130), .B(b[28]), .C(n574), .D(b_e[5]), .Y(n1212) );
  scg2d1_hd U952 ( .A(n1130), .B(b[29]), .C(n575), .D(b_e[6]), .Y(n1213) );
  nid1_hd U953 ( .A(n1164), .Y(n1163) );
  xo2d1_hd U954 ( .A(n938), .B(n820), .Y(mult_x_1_n850) );
  xo2d1_hd U955 ( .A(n903), .B(n645), .Y(mult_x_1_n715) );
  xo2d1_hd U956 ( .A(n931), .B(n785), .Y(mult_x_1_n823) );
  xo2d1_hd U957 ( .A(n910), .B(n680), .Y(mult_x_1_n742) );
  xo2d1_hd U958 ( .A(n917), .B(n715), .Y(mult_x_1_n769) );
  xo2d1_hd U959 ( .A(n917), .B(n719), .Y(mult_x_1_n770) );
  xo2d1_hd U960 ( .A(n924), .B(n750), .Y(mult_x_1_n796) );
  xo2d1_hd U961 ( .A(n910), .B(n684), .Y(mult_x_1_n743) );
  xo2d1_hd U962 ( .A(n938), .B(n824), .Y(mult_x_1_n851) );
  nid1_hd U963 ( .A(n1215), .Y(n1140) );
  nid1_hd U964 ( .A(n1153), .Y(n1152) );
  nid1_hd U965 ( .A(n1111), .Y(n1112) );
  ad2d1_hd U966 ( .A(n519), .B(a_e[8]), .Y(n577) );
  nid1_hd U967 ( .A(n1098), .Y(n1096) );
  nid1_hd U968 ( .A(n1149), .Y(n1153) );
  nid1_hd U969 ( .A(n1104), .Y(n1105) );
  ad2d1_hd U970 ( .A(DP_OP_125J2_130_6300_n54), .B(n1205), .Y(
        DP_OP_125J2_130_6300_I5) );
  xo2d1_hd U971 ( .A(n903), .B(n651), .Y(mult_x_1_n717) );
  xo2d1_hd U972 ( .A(n924), .B(n756), .Y(mult_x_1_n798) );
  nid1_hd U973 ( .A(n716), .Y(n1085) );
  xo2d1_hd U974 ( .A(n917), .B(n721), .Y(mult_x_1_n771) );
  nid1_hd U975 ( .A(n1123), .Y(n1126) );
  xo2d1_hd U976 ( .A(n910), .B(n686), .Y(mult_x_1_n744) );
  nid1_hd U977 ( .A(n788), .Y(n1104) );
  nid1_hd U978 ( .A(n681), .Y(n1077) );
  xo2d1_hd U979 ( .A(n931), .B(n791), .Y(mult_x_1_n825) );
  nid1_hd U980 ( .A(n681), .Y(n1078) );
  xo2d1_hd U981 ( .A(n938), .B(n826), .Y(mult_x_1_n852) );
  nid1_hd U982 ( .A(n823), .Y(n1111) );
  nid1_hd U983 ( .A(n646), .Y(n1070) );
  xo2d1_hd U984 ( .A(n896), .B(n616), .Y(mult_x_1_n690) );
  nid1_hd U985 ( .A(n646), .Y(n1069) );
  nid1_hd U986 ( .A(n751), .Y(n1092) );
  nid1_hd U987 ( .A(n716), .Y(n1086) );
  nid1_hd U988 ( .A(n646), .Y(n1068) );
  nid1_hd U989 ( .A(n857), .Y(n1123) );
  or2d1_hd U990 ( .A(n798), .B(n825), .Y(n822) );
  nid1_hd U991 ( .A(n378), .Y(n1165) );
  ad2d1_hd U992 ( .A(n576), .B(b_e[8]), .Y(n578) );
  or2d1_hd U993 ( .A(n763), .B(n790), .Y(n787) );
  nid1_hd U994 ( .A(n855), .Y(n1120) );
  ad2d1_hd U995 ( .A(n1009), .B(n890), .Y(mult_x_1_n581) );
  ad2d1_hd U996 ( .A(n1047), .B(n890), .Y(mult_x_1_n588) );
  ad4d1_hd U997 ( .A(n1235), .B(n1234), .C(n1233), .D(n1232), .Y(n1236) );
  ad2d1_hd U998 ( .A(n1054), .B(n890), .Y(mult_x_1_n590) );
  ad2d1_hd U999 ( .A(n1037), .B(n890), .Y(mult_x_1_n586) );
  ad2d1_hd U1000 ( .A(n1042), .B(n890), .Y(mult_x_1_n587) );
  nid1_hd U1001 ( .A(n853), .Y(n1116) );
  or2d1_hd U1002 ( .A(n1289), .B(n1291), .Y(n1216) );
  ad2d1_hd U1003 ( .A(n977), .B(n889), .Y(mult_x_1_n574) );
  ad2d1_hd U1004 ( .A(b_m[8]), .B(n889), .Y(mult_x_1_n583) );
  ad2d1_hd U1005 ( .A(n982), .B(n889), .Y(mult_x_1_n575) );
  ad2d1_hd U1006 ( .A(n962), .B(a_m[23]), .Y(mult_x_1_n571) );
  ad2d1_hd U1007 ( .A(n1004), .B(n889), .Y(mult_x_1_n580) );
  ad2d1_hd U1008 ( .A(n1052), .B(n889), .Y(mult_x_1_n589) );
  or2d1_hd U1009 ( .A(state[2]), .B(n463), .Y(n1294) );
  ad2d1_hd U1010 ( .A(n992), .B(n889), .Y(mult_x_1_n577) );
  ad4d1_hd U1011 ( .A(n1227), .B(n1226), .C(n1225), .D(n1224), .Y(n1228) );
  nid1_hd U1012 ( .A(n962), .Y(n959) );
  nid1_hd U1013 ( .A(n1014), .Y(n1016) );
  nid1_hd U1014 ( .A(n1052), .Y(n1049) );
  nid1_hd U1015 ( .A(n1033), .Y(n1030) );
  nid1_hd U1016 ( .A(n1042), .Y(n1039) );
  nid1_hd U1017 ( .A(n1037), .Y(n1034) );
  nid1_hd U1018 ( .A(n1032), .Y(n1029) );
  nid1_hd U1019 ( .A(n1027), .Y(n1024) );
  nid1_hd U1020 ( .A(n1047), .Y(n1044) );
  nid1_hd U1021 ( .A(n1009), .Y(n1011) );
  nid1_hd U1022 ( .A(b_m[10]), .Y(n1012) );
  ad2d1_hd U1023 ( .A(i_Z_ACK), .B(o_Z_STB), .Y(n177) );
  nid1_hd U1024 ( .A(b_m[9]), .Y(n1017) );
  nid1_hd U1025 ( .A(b_m[1]), .Y(n1057) );
  nid1_hd U1026 ( .A(b_m[11]), .Y(n1007) );
  nid1_hd U1027 ( .A(b_m[9]), .Y(n1015) );
  nid1_hd U1028 ( .A(b_m[12]), .Y(n1002) );
  nid1_hd U1029 ( .A(b_m[10]), .Y(n1010) );
  or4d1_hd U1030 ( .A(product[20]), .B(product[9]), .C(product[7]), .D(
        product[23]), .Y(n1392) );
  nid1_hd U1031 ( .A(b_m[13]), .Y(n997) );
  nid1_hd U1032 ( .A(b_m[11]), .Y(n1005) );
  nid1_hd U1033 ( .A(b_m[12]), .Y(n1000) );
  nid1_hd U1034 ( .A(b_m[13]), .Y(n995) );
  nid1_hd U1035 ( .A(b_m[21]), .Y(n957) );
  nid1_hd U1036 ( .A(b_m[14]), .Y(n992) );
  nid1_hd U1037 ( .A(b_m[20]), .Y(n962) );
  nid1_hd U1038 ( .A(b_m[7]), .Y(n1027) );
  or4d1_hd U1039 ( .A(b_e[1]), .B(n14), .C(b_e[4]), .D(b_e[2]), .Y(n1231) );
  or4d1_hd U1040 ( .A(a_e[1]), .B(n10), .C(a_e[4]), .D(a_e[2]), .Y(n1223) );
  ivd1_hd U1041 ( .A(a_m[0]), .Y(n387) );
  ivd1_hd U1042 ( .A(n387), .Y(n388) );
  ivd1_hd U1043 ( .A(z_m[7]), .Y(n389) );
  ivd1_hd U1044 ( .A(n389), .Y(n390) );
  ivd1_hd U1045 ( .A(z_m[3]), .Y(n391) );
  ivd1_hd U1046 ( .A(n391), .Y(n392) );
  ivd1_hd U1047 ( .A(z_m[5]), .Y(n393) );
  ivd1_hd U1048 ( .A(n393), .Y(n394) );
  ivd1_hd U1049 ( .A(z_m[11]), .Y(n395) );
  ivd1_hd U1050 ( .A(n395), .Y(n396) );
  ivd1_hd U1051 ( .A(z_m[13]), .Y(n397) );
  ivd1_hd U1052 ( .A(n397), .Y(n398) );
  ivd1_hd U1053 ( .A(z_m[9]), .Y(n399) );
  ivd1_hd U1054 ( .A(n399), .Y(n400) );
  ivd1_hd U1055 ( .A(z_m[15]), .Y(n401) );
  ivd1_hd U1056 ( .A(n401), .Y(n402) );
  ivd1_hd U1057 ( .A(z_m[19]), .Y(n403) );
  ivd1_hd U1058 ( .A(n403), .Y(n404) );
  ivd1_hd U1059 ( .A(z_m[17]), .Y(n405) );
  ivd1_hd U1060 ( .A(n405), .Y(n406) );
  ivd1_hd U1061 ( .A(n461), .Y(n407) );
  ivd1_hd U1062 ( .A(mult_x_1_n662), .Y(n410) );
  ivd1_hd U1063 ( .A(n410), .Y(n411) );
  ivd1_hd U1064 ( .A(mult_x_1_n661), .Y(n412) );
  ivd1_hd U1065 ( .A(n412), .Y(n413) );
  ivd1_hd U1066 ( .A(mult_x_1_n660), .Y(n414) );
  ivd1_hd U1067 ( .A(n414), .Y(n415) );
  ivd1_hd U1068 ( .A(mult_x_1_n659), .Y(n416) );
  ivd1_hd U1069 ( .A(n416), .Y(n417) );
  ivd1_hd U1070 ( .A(mult_x_1_n658), .Y(n418) );
  ivd1_hd U1071 ( .A(n418), .Y(n419) );
  ivd1_hd U1072 ( .A(mult_x_1_n656), .Y(n420) );
  ivd1_hd U1073 ( .A(n420), .Y(n421) );
  ivd1_hd U1074 ( .A(mult_x_1_n657), .Y(n422) );
  ivd1_hd U1075 ( .A(n422), .Y(n423) );
  ivd1_hd U1076 ( .A(mult_x_1_n654), .Y(n424) );
  ivd1_hd U1077 ( .A(n424), .Y(n425) );
  ivd1_hd U1078 ( .A(mult_x_1_n655), .Y(n426) );
  ivd1_hd U1079 ( .A(n426), .Y(n427) );
  ivd1_hd U1080 ( .A(mult_x_1_n653), .Y(n428) );
  ivd1_hd U1081 ( .A(n428), .Y(n429) );
  ivd1_hd U1082 ( .A(mult_x_1_n652), .Y(n430) );
  ivd1_hd U1083 ( .A(n430), .Y(n431) );
  ivd1_hd U1084 ( .A(mult_x_1_n650), .Y(n432) );
  ivd1_hd U1085 ( .A(n432), .Y(n433) );
  ivd1_hd U1086 ( .A(mult_x_1_n651), .Y(n434) );
  ivd1_hd U1087 ( .A(n434), .Y(n435) );
  ivd1_hd U1088 ( .A(n436), .Y(n437) );
  ivd1_hd U1089 ( .A(n438), .Y(n439) );
  ivd1_hd U1090 ( .A(n440), .Y(n441) );
  ivd1_hd U1091 ( .A(mult_x_1_n663), .Y(n454) );
  ivd1_hd U1092 ( .A(n454), .Y(n455) );
  ivd1_hd U1093 ( .A(n1182), .Y(n456) );
  ivd1_hd U1094 ( .A(n456), .Y(n457) );
  ivd1_hd U1095 ( .A(n1199), .Y(n458) );
  ivd1_hd U1096 ( .A(n458), .Y(n459) );
  ivd1_hd U1097 ( .A(n1460), .Y(n460) );
  ivd1_hd U1098 ( .A(n1460), .Y(n461) );
  ivd1_hd U1099 ( .A(state[1]), .Y(n462) );
  ivd1_hd U1100 ( .A(n462), .Y(n463) );
  ivd1_hd U1101 ( .A(n579), .Y(n464) );
  ivd1_hd U1102 ( .A(n579), .Y(n465) );
  ivd1_hd U1103 ( .A(DP_OP_125J2_130_6300_I5), .Y(n466) );
  ivd1_hd U1104 ( .A(DP_OP_125J2_130_6300_I5), .Y(n467) );
  ivd1_hd U1105 ( .A(n110), .Y(n468) );
  ivd1_hd U1106 ( .A(n110), .Y(n469) );
  ivd1_hd U1107 ( .A(n472), .Y(n470) );
  ivd1_hd U1108 ( .A(n472), .Y(n471) );
  ivd1_hd U1109 ( .A(n1472), .Y(n472) );
  ivd1_hd U1110 ( .A(n1472), .Y(n473) );
  ivd1_hd U1111 ( .A(n1472), .Y(n474) );
  ivd1_hd U1112 ( .A(n1468), .Y(n475) );
  ivd1_hd U1113 ( .A(n1468), .Y(n476) );
  ivd1_hd U1114 ( .A(n1468), .Y(n477) );
  ivd1_hd U1115 ( .A(n1332), .Y(n478) );
  ivd1_hd U1116 ( .A(n1332), .Y(n479) );
  ivd1_hd U1117 ( .A(n1332), .Y(n480) );
  ivd1_hd U1118 ( .A(n1332), .Y(n481) );
  ivd1_hd U1119 ( .A(n579), .Y(n482) );
  ivd1_hd U1120 ( .A(n482), .Y(n483) );
  ivd1_hd U1121 ( .A(n482), .Y(n484) );
  ivd1_hd U1122 ( .A(n485), .Y(n487) );
  ivd1_hd U1123 ( .A(n485), .Y(n488) );
  ivd1_hd U1124 ( .A(n586), .Y(n489) );
  ivd1_hd U1125 ( .A(n586), .Y(n490) );
  ivd1_hd U1126 ( .A(n586), .Y(n491) );
  ivd1_hd U1127 ( .A(n586), .Y(n492) );
  ivd1_hd U1128 ( .A(n796), .Y(n493) );
  ivd1_hd U1129 ( .A(n796), .Y(n494) );
  ivd1_hd U1130 ( .A(n796), .Y(n495) );
  ivd1_hd U1131 ( .A(n796), .Y(n496) );
  ivd1_hd U1132 ( .A(n761), .Y(n497) );
  ivd1_hd U1133 ( .A(n761), .Y(n498) );
  ivd1_hd U1134 ( .A(n761), .Y(n499) );
  ivd1_hd U1135 ( .A(n761), .Y(n500) );
  ivd1_hd U1136 ( .A(n726), .Y(n501) );
  ivd1_hd U1137 ( .A(n726), .Y(n502) );
  ivd1_hd U1138 ( .A(n726), .Y(n503) );
  ivd1_hd U1139 ( .A(n726), .Y(n504) );
  ivd1_hd U1140 ( .A(n656), .Y(n505) );
  ivd1_hd U1141 ( .A(n656), .Y(n506) );
  ivd1_hd U1142 ( .A(n656), .Y(n507) );
  ivd1_hd U1143 ( .A(n656), .Y(n508) );
  ivd1_hd U1144 ( .A(n621), .Y(n509) );
  ivd1_hd U1145 ( .A(n621), .Y(n510) );
  ivd1_hd U1146 ( .A(n621), .Y(n511) );
  ivd1_hd U1147 ( .A(n621), .Y(n512) );
  ivd1_hd U1148 ( .A(n691), .Y(n513) );
  ivd1_hd U1149 ( .A(n691), .Y(n514) );
  ivd1_hd U1150 ( .A(n691), .Y(n515) );
  ivd1_hd U1151 ( .A(n691), .Y(n516) );
  ivd1_hd U1152 ( .A(n1216), .Y(n517) );
  ivd1_hd U1153 ( .A(n1216), .Y(n518) );
  ivd1_hd U1154 ( .A(n1216), .Y(n519) );
  ivd1_hd U1155 ( .A(n1363), .Y(n520) );
  ivd1_hd U1156 ( .A(n1363), .Y(n521) );
  ivd1_hd U1157 ( .A(n1363), .Y(n522) );
  ivd1_hd U1158 ( .A(n1363), .Y(n523) );
  nid1_hd U1159 ( .A(n1285), .Y(n524) );
  ivd1_hd U1160 ( .A(n1331), .Y(n526) );
  scg2d1_hd U1161 ( .A(C81_DATA2_6), .B(n459), .C(a_e[6]), .D(n526), .Y(n312)
         );
  scg2d1_hd U1162 ( .A(C81_DATA2_5), .B(n1199), .C(a_e[5]), .D(n1202), .Y(n313) );
  scg2d1_hd U1163 ( .A(C81_DATA2_4), .B(n459), .C(a_e[4]), .D(n1202), .Y(n314)
         );
  scg2d1_hd U1164 ( .A(C81_DATA2_3), .B(n459), .C(a_e[3]), .D(n1202), .Y(n315)
         );
  scg2d1_hd U1165 ( .A(C81_DATA2_2), .B(n459), .C(n526), .D(a_e[2]), .Y(n316)
         );
  ivd1_hd U1166 ( .A(n1297), .Y(n527) );
  scg2d1_hd U1167 ( .A(C82_DATA2_6), .B(n457), .C(b_e[6]), .D(n527), .Y(n321)
         );
  scg2d1_hd U1168 ( .A(C82_DATA2_5), .B(n1182), .C(b_e[5]), .D(n1186), .Y(n322) );
  scg2d1_hd U1169 ( .A(C82_DATA2_4), .B(n457), .C(b_e[4]), .D(n1186), .Y(n323)
         );
  scg2d1_hd U1170 ( .A(C82_DATA2_3), .B(n457), .C(b_e[3]), .D(n1186), .Y(n324)
         );
  scg2d1_hd U1171 ( .A(C82_DATA2_2), .B(n457), .C(n527), .D(b_e[2]), .Y(n325)
         );
  ivd1_hd U1172 ( .A(n475), .Y(n528) );
  ivd1_hd U1173 ( .A(n477), .Y(n529) );
  ivd1_hd U1174 ( .A(n476), .Y(n530) );
  ivd1_hd U1175 ( .A(n1252), .Y(n531) );
  ivd1_hd U1176 ( .A(n1252), .Y(n532) );
  ivd1_hd U1177 ( .A(n1252), .Y(n533) );
  ivd1_hd U1178 ( .A(n1252), .Y(n534) );
  scg2d1_hd U1179 ( .A(z_m[19]), .B(n532), .C(n1160), .D(z[19]), .Y(n241) );
  scg2d1_hd U1180 ( .A(z_m[18]), .B(n531), .C(n1158), .D(z[18]), .Y(n242) );
  scg2d1_hd U1181 ( .A(n406), .B(n534), .C(n1158), .D(z[17]), .Y(n243) );
  scg2d1_hd U1182 ( .A(z_m[16]), .B(n533), .C(n1158), .D(z[16]), .Y(n244) );
  scg2d1_hd U1183 ( .A(z_m[15]), .B(n532), .C(n1158), .D(z[15]), .Y(n245) );
  scg2d1_hd U1184 ( .A(z_m[14]), .B(n531), .C(n1158), .D(z[14]), .Y(n246) );
  scg2d1_hd U1185 ( .A(n398), .B(n534), .C(n1159), .D(z[13]), .Y(n247) );
  scg2d1_hd U1186 ( .A(z_m[12]), .B(n533), .C(n1159), .D(z[12]), .Y(n248) );
  scg2d1_hd U1187 ( .A(z_m[11]), .B(n532), .C(n1159), .D(z[11]), .Y(n249) );
  scg2d1_hd U1188 ( .A(z_m[10]), .B(n531), .C(n1159), .D(z[10]), .Y(n250) );
  scg2d1_hd U1189 ( .A(n400), .B(n534), .C(n1159), .D(z[9]), .Y(n251) );
  scg2d1_hd U1190 ( .A(z_m[8]), .B(n533), .C(n1159), .D(z[8]), .Y(n252) );
  scg2d1_hd U1191 ( .A(z_m[7]), .B(n532), .C(n1160), .D(z[7]), .Y(n253) );
  scg2d1_hd U1192 ( .A(z_m[6]), .B(n531), .C(n1160), .D(z[6]), .Y(n254) );
  scg2d1_hd U1193 ( .A(n394), .B(n534), .C(n1160), .D(z[5]), .Y(n255) );
  scg2d1_hd U1194 ( .A(z_m[4]), .B(n533), .C(n1160), .D(z[4]), .Y(n256) );
  scg2d1_hd U1195 ( .A(z_m[3]), .B(n532), .C(n1160), .D(z[3]), .Y(n257) );
  scg2d1_hd U1196 ( .A(z_m[2]), .B(n531), .C(n1161), .D(z[2]), .Y(n258) );
  scg2d1_hd U1197 ( .A(z_m[1]), .B(n534), .C(n1161), .D(z[1]), .Y(n259) );
  scg2d1_hd U1198 ( .A(z_m[0]), .B(n533), .C(n1161), .D(z[0]), .Y(n260) );
  scg2d1_hd U1199 ( .A(z_m[21]), .B(n532), .C(n1161), .D(z[21]), .Y(n239) );
  scg2d1_hd U1200 ( .A(z_m[20]), .B(n531), .C(n1158), .D(z[20]), .Y(n240) );
  or2d1_hd U1201 ( .A(n1216), .B(n1144), .Y(n1325) );
  ivd1_hd U1202 ( .A(n1325), .Y(n535) );
  ivd1_hd U1203 ( .A(n1325), .Y(n536) );
  ivd1_hd U1204 ( .A(n1325), .Y(n537) );
  ivd1_hd U1205 ( .A(n1325), .Y(n538) );
  ivd1_hd U1206 ( .A(n856), .Y(n539) );
  ivd1_hd U1207 ( .A(n856), .Y(n540) );
  ivd1_hd U1208 ( .A(n856), .Y(n541) );
  ivd1_hd U1209 ( .A(n856), .Y(n542) );
  ivd1_hd U1210 ( .A(n822), .Y(n543) );
  ivd1_hd U1211 ( .A(n822), .Y(n544) );
  ivd1_hd U1212 ( .A(n822), .Y(n545) );
  ivd1_hd U1213 ( .A(n822), .Y(n546) );
  ivd1_hd U1214 ( .A(n787), .Y(n547) );
  ivd1_hd U1215 ( .A(n787), .Y(n548) );
  ivd1_hd U1216 ( .A(n787), .Y(n549) );
  ivd1_hd U1217 ( .A(n787), .Y(n550) );
  ivd1_hd U1218 ( .A(n752), .Y(n551) );
  ivd1_hd U1219 ( .A(n752), .Y(n552) );
  ivd1_hd U1220 ( .A(n752), .Y(n553) );
  ivd1_hd U1221 ( .A(n752), .Y(n554) );
  ivd1_hd U1222 ( .A(n682), .Y(n555) );
  ivd1_hd U1223 ( .A(n682), .Y(n556) );
  ivd1_hd U1224 ( .A(n682), .Y(n557) );
  ivd1_hd U1225 ( .A(n682), .Y(n558) );
  ivd1_hd U1226 ( .A(n647), .Y(n559) );
  ivd1_hd U1227 ( .A(n647), .Y(n560) );
  ivd1_hd U1228 ( .A(n647), .Y(n561) );
  ivd1_hd U1229 ( .A(n647), .Y(n562) );
  ivd1_hd U1230 ( .A(n717), .Y(n563) );
  ivd1_hd U1231 ( .A(n717), .Y(n564) );
  ivd1_hd U1232 ( .A(n717), .Y(n565) );
  ivd1_hd U1233 ( .A(n717), .Y(n566) );
  ivd1_hd U1234 ( .A(n613), .Y(n567) );
  ivd1_hd U1235 ( .A(n613), .Y(n568) );
  ivd1_hd U1236 ( .A(n613), .Y(n569) );
  ivd1_hd U1237 ( .A(n613), .Y(n570) );
  or3d1_hd U1238 ( .A(n1291), .B(n1221), .C(n462), .Y(DP_OP_125J2_130_6300_n54) );
  ivd1_hd U1239 ( .A(DP_OP_125J2_130_6300_n54), .Y(n571) );
  ivd1_hd U1240 ( .A(DP_OP_125J2_130_6300_n54), .Y(n572) );
  ivd1_hd U1241 ( .A(DP_OP_125J2_130_6300_n54), .Y(n573) );
  scg2d1_hd U1242 ( .A(n572), .B(round_bit), .C(n29), .D(z_m[0]), .Y(n1383) );
  xo2d1_hd U1243 ( .A(DP_OP_125J2_130_6300_n33), .B(n571), .Y(
        DP_OP_125J2_130_6300_n1) );
  or2d1_hd U1244 ( .A(n1172), .B(state[1]), .Y(n1217) );
  ivd1_hd U1245 ( .A(n1217), .Y(n574) );
  ivd1_hd U1246 ( .A(n1217), .Y(n575) );
  ivd1_hd U1247 ( .A(n1217), .Y(n576) );
  scg2d1_hd U1248 ( .A(n1131), .B(b[24]), .C(n574), .D(b_e[1]), .Y(n1208) );
  scg2d1_hd U1249 ( .A(n1131), .B(b[25]), .C(n576), .D(b_e[2]), .Y(n1209) );
  scg2d1_hd U1250 ( .A(n1130), .B(b[26]), .C(n574), .D(b_e[3]), .Y(n1210) );
  scg2d1_hd U1251 ( .A(n1130), .B(b[27]), .C(n575), .D(b_e[4]), .Y(n1211) );
  nr2bd1_hd U1252 ( .AN(n685), .B(n653), .Y(n681) );
  nr2bd1_hd U1253 ( .AN(n658), .B(n685), .Y(n683) );
  nr2bd1_hd U1254 ( .AN(n650), .B(n618), .Y(n646) );
  nr2bd1_hd U1255 ( .AN(n623), .B(n650), .Y(n648) );
  nd2bd1_hd U1256 ( .AN(state[3]), .B(state[0]), .Y(n1291) );
  nr2bd1_hd U1257 ( .AN(n825), .B(n793), .Y(n821) );
  nr2bd1_hd U1258 ( .AN(n790), .B(n758), .Y(n786) );
  nr2bd1_hd U1259 ( .AN(n763), .B(n790), .Y(n788) );
  ivd1_hd U1260 ( .A(n932), .Y(n938) );
  nr2bd1_hd U1261 ( .AN(n755), .B(n723), .Y(n751) );
  nr2bd1_hd U1262 ( .AN(n728), .B(n755), .Y(n753) );
  nr2bd1_hd U1263 ( .AN(n720), .B(n688), .Y(n716) );
  scg4d1_hd U1264 ( .A(n612), .B(mult_x_1_n643), .C(n492), .D(b_m[19]), .E(
        n567), .F(n953), .G(b_m[20]), .H(n1060), .Y(n591) );
  ivd1_hd U1265 ( .A(n888), .Y(n893) );
  ivd1_hd U1266 ( .A(n888), .Y(n891) );
  ivd1_hd U1267 ( .A(n1489), .Y(n1164) );
  ivd1_hd U1268 ( .A(n1258), .Y(n1293) );
  ivd1_hd U1269 ( .A(n1398), .Y(n1483) );
  ivd1_hd U1270 ( .A(n1297), .Y(n1186) );
  scg14d1_hd U1271 ( .A(n1297), .B(n575), .C(n479), .Y(n1182) );
  ivd1_hd U1272 ( .A(n1333), .Y(n1361) );
  ivd1_hd U1273 ( .A(n1331), .Y(n1202) );
  scg14d1_hd U1274 ( .A(n1331), .B(n518), .C(n480), .Y(n1199) );
  ivd1_hd U1275 ( .A(n1301), .Y(n1327) );
  ivd1_hd U1276 ( .A(n478), .Y(n1215) );
  ivd1_hd U1277 ( .A(n1294), .Y(n1170) );
  ivd1_hd U1278 ( .A(n1291), .Y(n1171) );
  ivd1_hd U1279 ( .A(n939), .Y(n942) );
  ivd1_hd U1280 ( .A(n940), .Y(n943) );
  ivd1_hd U1281 ( .A(n939), .Y(n941) );
  nr2bd1_hd U1282 ( .AN(n798), .B(n825), .Y(n823) );
  ivd1_hd U1283 ( .A(n887), .Y(n894) );
  ivd1_hd U1284 ( .A(n947), .Y(n951) );
  ivd1_hd U1285 ( .A(n888), .Y(n890) );
  ivd1_hd U1286 ( .A(a_m[21]), .Y(n876) );
  ivd1_hd U1287 ( .A(n488), .Y(n862) );
  ivd1_hd U1288 ( .A(n888), .Y(n892) );
  ivd1_hd U1289 ( .A(n1164), .Y(n1158) );
  ivd1_hd U1290 ( .A(n1164), .Y(n1161) );
  scg20d1_hd U1291 ( .A(n1258), .B(n1257), .C(n1256), .Y(n1285) );
  ivd1_hd U1292 ( .A(n1163), .Y(n1159) );
  ivd1_hd U1293 ( .A(n1163), .Y(n1160) );
  ivd1_hd U1294 ( .A(n1330), .Y(n1338) );
  ivd1_hd U1295 ( .A(n940), .Y(n944) );
  ivd1_hd U1296 ( .A(n933), .Y(n936) );
  ivd1_hd U1297 ( .A(n933), .Y(n935) );
  ivd1_hd U1298 ( .A(n932), .Y(n934) );
  ivd1_hd U1299 ( .A(n926), .Y(n929) );
  ivd1_hd U1300 ( .A(n932), .Y(n937) );
  ivd1_hd U1301 ( .A(n926), .Y(n927) );
  ivd1_hd U1302 ( .A(n926), .Y(n930) );
  ivd1_hd U1303 ( .A(n919), .Y(n921) );
  ivd1_hd U1304 ( .A(n905), .Y(n908) );
  ivd1_hd U1305 ( .A(n912), .Y(n914) );
  nid2_hd U1306 ( .A(n1095), .Y(n1097) );
  ivd1_hd U1307 ( .A(n898), .Y(n901) );
  ivd1_hd U1308 ( .A(n905), .Y(n907) );
  ivd1_hd U1309 ( .A(n887), .Y(n895) );
  ivd1_hd U1310 ( .A(a_m[2]), .Y(n940) );
  ivd1_hd U1311 ( .A(n898), .Y(n900) );
  ivd1_hd U1312 ( .A(n947), .Y(n949) );
  ivd1_hd U1313 ( .A(n947), .Y(n950) );
  ivd1_hd U1314 ( .A(a_m[22]), .Y(n877) );
  ivd1_hd U1315 ( .A(n1164), .Y(n1162) );
  nd2bd1_hd U1316 ( .AN(n1294), .B(n1304), .Y(n155) );
  scg21d1_hd U1317 ( .A(n1296), .B(n1338), .C(n1293), .D(n1256), .Y(n1489) );
  nr2d1_hd U1318 ( .A(n1384), .B(n1394), .Y(n1484) );
  ivd1_hd U1319 ( .A(n105), .Y(n1384) );
  nr3d1_hd U1320 ( .A(n1291), .B(n463), .C(n1221), .Y(n1214) );
  ivd1_hd U1321 ( .A(z_m[23]), .Y(n1373) );
  nr2d1_hd U1322 ( .A(n1294), .B(n1220), .Y(n1219) );
  oa21d1_hd U1323 ( .A(n1334), .B(n1328), .C(n1148), .Y(n1297) );
  ivd1_hd U1324 ( .A(DP_OP_116J2_127_7148_n3), .Y(n1181) );
  oa21d1_hd U1325 ( .A(n1329), .B(n1328), .C(n1144), .Y(n1331) );
  nd3d1_hd U1326 ( .A(n1330), .B(n1296), .C(n1295), .Y(n1328) );
  ivd1_hd U1327 ( .A(DP_OP_113J2_124_6892_n3), .Y(n1193) );
  nd2bd1_hd U1328 ( .AN(state[2]), .B(n463), .Y(n1289) );
  ivd1_hd U1329 ( .A(a_m[1]), .Y(n863) );
  ivd1_hd U1330 ( .A(n925), .Y(n928) );
  ivd1_hd U1331 ( .A(n919), .Y(n922) );
  ivd1_hd U1332 ( .A(n912), .Y(n915) );
  nid2_hd U1333 ( .A(n1103), .Y(n1106) );
  ivd1_hd U1334 ( .A(n918), .Y(n920) );
  ivd1_hd U1335 ( .A(n918), .Y(n923) );
  ivd1_hd U1336 ( .A(n911), .Y(n913) );
  ivd1_hd U1337 ( .A(n911), .Y(n916) );
  ivd1_hd U1338 ( .A(n904), .Y(n906) );
  ivd1_hd U1339 ( .A(n904), .Y(n909) );
  ivd1_hd U1340 ( .A(n897), .Y(n899) );
  ivd1_hd U1341 ( .A(n886), .Y(n889) );
  scg14d1_hd U1342 ( .A(n957), .B(n521), .C(n1362), .Y(n287) );
  scg14d1_hd U1343 ( .A(n1027), .B(n520), .C(n1348), .Y(n300) );
  scg14d1_hd U1344 ( .A(n972), .B(n521), .C(n1359), .Y(n289) );
  ivd1_hd U1345 ( .A(n1275), .Y(n1282) );
  scg22d1_hd U1346 ( .A(z_e[1]), .B(n1255), .C(z_e[0]), .D(n1293), .Y(n1275)
         );
  oa21d1_hd U1347 ( .A(z_e[8]), .B(z_e[7]), .C(n1222), .Y(n1257) );
  ivd1_hd U1348 ( .A(z_e[9]), .Y(n1222) );
  scg14d1_hd U1349 ( .A(n1386), .B(n1484), .C(n1385), .Y(n284) );
  scg4d1_hd U1350 ( .A(n1406), .B(z_m[2]), .C(n1405), .D(z_m[1]), .E(n392), 
        .F(n1154), .G(n1152), .H(product[28]), .Y(n281) );
  ivd1_hd U1351 ( .A(z_m[21]), .Y(n1481) );
  ivd1_hd U1352 ( .A(net908), .Y(n1386) );
  scg17d1_hd U1353 ( .A(n470), .B(z_m[8]), .C(n1432), .D(n1431), .Y(n274) );
  scg17d1_hd U1354 ( .A(n471), .B(z_m[12]), .C(n1447), .D(n1446), .Y(n270) );
  scg17d1_hd U1355 ( .A(n470), .B(z_m[4]), .C(n1417), .D(n1416), .Y(n278) );
  scg17d1_hd U1356 ( .A(n471), .B(z_m[16]), .C(n1463), .D(n1462), .Y(n266) );
  scg4d1_hd U1357 ( .A(n1436), .B(z_m[10]), .C(n1435), .D(n400), .E(n396), .F(
        n1157), .G(n1152), .H(product[36]), .Y(n273) );
  scg4d1_hd U1358 ( .A(n1421), .B(z_m[6]), .C(n1420), .D(n394), .E(n390), .F(
        n1157), .G(n1151), .H(product[32]), .Y(n277) );
  scg4d1_hd U1359 ( .A(n1451), .B(z_m[14]), .C(n1450), .D(n398), .E(n402), .F(
        n1157), .G(n1152), .H(product[40]), .Y(n269) );
  scg4d1_hd U1360 ( .A(n1467), .B(z_m[18]), .C(n1466), .D(n406), .E(n404), .F(
        n1154), .G(n1153), .H(product[44]), .Y(n265) );
  scg4d1_hd U1361 ( .A(n1444), .B(z_m[12]), .C(n1443), .D(z_m[11]), .E(z_m[13]), .F(n1154), .G(n1152), .H(product[38]), .Y(n271) );
  scg4d1_hd U1362 ( .A(n1459), .B(z_m[16]), .C(n1458), .D(z_m[15]), .E(z_m[17]), .F(n1157), .G(n1149), .H(product[42]), .Y(n267) );
  scg4d1_hd U1363 ( .A(n1429), .B(z_m[8]), .C(n1428), .D(z_m[7]), .E(z_m[9]), 
        .F(n1157), .G(n1152), .H(product[34]), .Y(n275) );
  scg4d1_hd U1364 ( .A(n1414), .B(z_m[4]), .C(n1413), .D(z_m[3]), .E(z_m[5]), 
        .F(n1157), .G(n1152), .H(product[30]), .Y(n279) );
  scg12d1_hd U1365 ( .A(z_m[18]), .B(n406), .C(n1461), .Y(n1469) );
  scg12d1_hd U1366 ( .A(z_m[14]), .B(n398), .C(n1445), .Y(n1452) );
  scg12d1_hd U1367 ( .A(z_m[10]), .B(n400), .C(n1430), .Y(n1437) );
  scg12d1_hd U1368 ( .A(z_m[6]), .B(n394), .C(n1415), .Y(n1422) );
  ivd1_hd U1369 ( .A(z_m[22]), .Y(n1374) );
  ivd1_hd U1370 ( .A(state[2]), .Y(n1221) );
  nr2d1_hd U1371 ( .A(n1375), .B(n1151), .Y(n1393) );
  ivd1_hd U1372 ( .A(n1172), .Y(n1218) );
  ivd1_hd U1373 ( .A(state[0]), .Y(n34) );
  ivd1_hd U1374 ( .A(state[3]), .Y(n1220) );
  ivd1_hd U1375 ( .A(z_m[0]), .Y(n1380) );
  oa21d1_hd U1376 ( .A(n1217), .B(b_m[23]), .C(n481), .Y(n1333) );
  oa21d1_hd U1377 ( .A(n1216), .B(a_m[23]), .C(n478), .Y(n1301) );
  nr2d1_hd U1378 ( .A(n1245), .B(n1248), .Y(n1296) );
  nr2d1_hd U1379 ( .A(n1334), .B(n1244), .Y(n1248) );
  nd4d1_hd U1380 ( .A(n1241), .B(b_e[8]), .C(b_e[9]), .D(b_e[0]), .Y(n1334) );
  nr2d1_hd U1381 ( .A(n1329), .B(n1247), .Y(n1245) );
  nr2d1_hd U1382 ( .A(state[2]), .B(n1290), .Y(n1330) );
  nr2d1_hd U1383 ( .A(state[3]), .B(state[0]), .Y(n1304) );
  nd4d1_hd U1384 ( .A(n1239), .B(a_e[8]), .C(a_e[9]), .D(a_e[0]), .Y(n1329) );
  nr2d1_hd U1385 ( .A(n388), .B(n863), .Y(n855) );
  nr3d1_hd U1386 ( .A(a_m[1]), .B(a_m[0]), .C(n940), .Y(n853) );
  ivd1_hd U1387 ( .A(a_m[3]), .Y(n864) );
  ivd1_hd U1388 ( .A(a_m[4]), .Y(n865) );
  ao22d1_hd U1389 ( .A(n938), .B(n866), .C(a_m[6]), .D(n933), .Y(n790) );
  ivd1_hd U1390 ( .A(a_m[6]), .Y(n866) );
  ivd1_hd U1391 ( .A(a_m[7]), .Y(n867) );
  ivd1_hd U1392 ( .A(a_m[9]), .Y(n868) );
  ivd1_hd U1393 ( .A(a_m[12]), .Y(n870) );
  ivd1_hd U1394 ( .A(a_m[15]), .Y(n872) );
  ivd1_hd U1395 ( .A(n897), .Y(n902) );
  nr2d1_hd U1396 ( .A(n1338), .B(n1295), .Y(n1256) );
  nr3d1_hd U1397 ( .A(state[2]), .B(state[0]), .C(n1220), .Y(n1303) );
  ao22d1_hd U1398 ( .A(n945), .B(n864), .C(a_m[3]), .D(n940), .Y(n825) );
  ivd1_hd U1399 ( .A(a_e[0]), .Y(n1198) );
  ivd1_hd U1400 ( .A(b_e[0]), .Y(n1178) );
  ao22d1_hd U1401 ( .A(n1194), .B(n459), .C(a_e[7]), .D(n526), .Y(n141) );
  ao22d1_hd U1402 ( .A(n1183), .B(n457), .C(b_e[7]), .D(n527), .Y(n151) );
  oa21d1_hd U1403 ( .A(n480), .B(n1174), .C(n1173), .Y(n1207) );
  ivd1_hd U1404 ( .A(b[23]), .Y(n1174) );
  nr2d1_hd U1405 ( .A(n1246), .B(n1243), .Y(n1295) );
  nr4d1_hd U1406 ( .A(b_e[9]), .B(b_e[8]), .C(b_e[0]), .D(n1242), .Y(n1243) );
  nr4d1_hd U1407 ( .A(a_e[9]), .B(a_e[8]), .C(a_e[0]), .D(n1240), .Y(n1246) );
  oa21d1_hd U1408 ( .A(n479), .B(n1190), .C(n1189), .Y(n1206) );
  ivd1_hd U1409 ( .A(a[23]), .Y(n1190) );
  oa22d1_hd U1410 ( .A(n458), .B(n1206), .C(n1331), .D(n1198), .Y(n318) );
  scg15d1_hd U1411 ( .A(n1199), .B(C81_DATA2_1), .C(n1191), .D(n138), .Y(n317)
         );
  oa22d1_hd U1412 ( .A(n456), .B(n1207), .C(n1297), .D(n1178), .Y(n327) );
  scg15d1_hd U1413 ( .A(n1182), .B(C82_DATA2_1), .C(n1179), .D(n148), .Y(n326)
         );
  ivd1_hd U1414 ( .A(n1219), .Y(n1205) );
  oa21d1_hd U1415 ( .A(n1193), .B(n1192), .C(n1195), .Y(n1194) );
  oa21d1_hd U1416 ( .A(n1181), .B(n1180), .C(n1185), .Y(n1183) );
  oa211d1_hd U1417 ( .A(n1197), .B(n458), .C(n138), .D(n1196), .Y(n311) );
  ao21d1_hd U1418 ( .A(n577), .B(n1195), .C(n1200), .Y(n1197) );
  oa211d1_hd U1419 ( .A(n1188), .B(n456), .C(n148), .D(n1187), .Y(n320) );
  ao21d1_hd U1420 ( .A(n578), .B(n1185), .C(n1184), .Y(n1188) );
  oa211d1_hd U1421 ( .A(n1177), .B(n456), .C(n148), .D(n1176), .Y(n356) );
  nr2d1_hd U1422 ( .A(n1185), .B(n578), .Y(n1184) );
  ao22d1_hd U1423 ( .A(n1130), .B(b[30]), .C(n576), .D(b_e[7]), .Y(n1180) );
  oa211d1_hd U1424 ( .A(n1204), .B(n458), .C(n138), .D(n1203), .Y(n319) );
  nr2d1_hd U1425 ( .A(n1195), .B(n577), .Y(n1200) );
  ao22d1_hd U1426 ( .A(n1130), .B(a[30]), .C(n519), .D(a_e[7]), .Y(n1192) );
  ivd1_hd U1427 ( .A(n946), .Y(n948) );
  nr2d1_hd U1428 ( .A(n887), .B(n485), .Y(mult_x_1_n569) );
  nr2d1_hd U1429 ( .A(n887), .B(n465), .Y(mult_x_1_n591) );
  ao22d1_hd U1430 ( .A(n896), .B(a_m[22]), .C(n877), .D(n888), .Y(n588) );
  ao22d1_hd U1431 ( .A(a_m[22]), .B(n876), .C(a_m[21]), .D(n877), .Y(n583) );
  ao22d1_hd U1432 ( .A(n1066), .B(n525), .C(n952), .D(n491), .Y(n582) );
  oa211d1_hd U1433 ( .A(n485), .B(n586), .C(n585), .D(n584), .Y(n587) );
  scg4d1_hd U1434 ( .A(n612), .B(mult_x_1_n641), .C(n948), .D(n569), .E(n490), 
        .F(n953), .G(n1060), .H(n486), .Y(n589) );
  scg4d1_hd U1435 ( .A(n612), .B(mult_x_1_n642), .C(n1060), .D(n955), .E(n489), 
        .F(n962), .G(n568), .H(n488), .Y(n590) );
  scg4d1_hd U1436 ( .A(n1063), .B(mult_x_1_n644), .C(n491), .D(b_m[18]), .E(
        n962), .F(n570), .G(n965), .H(n1060), .Y(n592) );
  scg4d1_hd U1437 ( .A(n1065), .B(mult_x_1_n645), .C(n490), .D(b_m[17]), .E(
        n967), .F(n569), .G(n970), .H(n1059), .Y(n593) );
  scg4d1_hd U1438 ( .A(n1065), .B(mult_x_1_n646), .C(n489), .D(b_m[16]), .E(
        n972), .F(n568), .G(n975), .H(n1060), .Y(n594) );
  scg4d1_hd U1439 ( .A(n1065), .B(mult_x_1_n647), .C(n492), .D(b_m[15]), .E(
        n977), .F(n567), .G(n980), .H(n1062), .Y(n595) );
  scg4d1_hd U1440 ( .A(n1065), .B(mult_x_1_n648), .C(n491), .D(n989), .E(n982), 
        .F(n570), .G(n985), .H(n1062), .Y(n596) );
  scg4d1_hd U1441 ( .A(n1065), .B(mult_x_1_n649), .C(n490), .D(n996), .E(n987), 
        .F(n569), .G(n990), .H(n1062), .Y(n597) );
  scg4d1_hd U1442 ( .A(n1065), .B(mult_x_1_n650), .C(n489), .D(n1001), .E(n992), .F(n568), .G(n997), .H(n1062), .Y(n598) );
  scg4d1_hd U1443 ( .A(n1063), .B(mult_x_1_n651), .C(n492), .D(n1006), .E(n994), .F(n567), .G(n1002), .H(n1059), .Y(n599) );
  scg4d1_hd U1444 ( .A(n1063), .B(mult_x_1_n652), .C(n491), .D(n1011), .E(n999), .F(n570), .G(n1007), .H(n1061), .Y(n600) );
  scg4d1_hd U1445 ( .A(n1066), .B(mult_x_1_n653), .C(n490), .D(n1016), .E(
        n1004), .F(n569), .G(n1012), .H(n1061), .Y(n601) );
  scg4d1_hd U1446 ( .A(n1066), .B(mult_x_1_n654), .C(n489), .D(n1020), .E(
        n1009), .F(n568), .G(n1017), .H(n1061), .Y(n602) );
  scg4d1_hd U1447 ( .A(n1066), .B(mult_x_1_n655), .C(n492), .D(b_m[7]), .E(
        n1014), .F(n567), .G(n1021), .H(n1061), .Y(n603) );
  scg4d1_hd U1448 ( .A(n1063), .B(mult_x_1_n656), .C(n491), .D(n1033), .E(
        b_m[8]), .F(n570), .G(n1025), .H(n1061), .Y(n604) );
  scg4d1_hd U1449 ( .A(n1064), .B(mult_x_1_n657), .C(n490), .D(b_m[5]), .E(
        n1027), .F(n569), .G(n1030), .H(n1061), .Y(n605) );
  scg4d1_hd U1450 ( .A(n1064), .B(mult_x_1_n658), .C(n489), .D(b_m[4]), .E(
        n1032), .F(n568), .G(n1035), .H(n611), .Y(n606) );
  scg4d1_hd U1451 ( .A(n1063), .B(mult_x_1_n659), .C(n492), .D(n1048), .E(
        n1037), .F(n567), .G(n1040), .H(n611), .Y(n607) );
  scg4d1_hd U1452 ( .A(n1064), .B(mult_x_1_n660), .C(n491), .D(b_m[2]), .E(
        n1042), .F(n570), .G(n1045), .H(n1059), .Y(n608) );
  scg4d1_hd U1453 ( .A(n1064), .B(mult_x_1_n661), .C(n490), .D(b_m[1]), .E(
        n1047), .F(n569), .G(n1050), .H(n1059), .Y(n609) );
  scg4d1_hd U1454 ( .A(n1064), .B(mult_x_1_n662), .C(n489), .D(n483), .E(n1052), .F(n568), .G(b_m[1]), .H(n1062), .Y(n610) );
  scg5d1_hd U1455 ( .A(n567), .B(b_m[1]), .C(n1064), .D(mult_x_1_n663), .E(
        n579), .F(n1060), .Y(n614) );
  nr2d1_hd U1456 ( .A(n615), .B(n465), .Y(n616) );
  ao22d1_hd U1457 ( .A(n903), .B(a_m[19]), .C(n875), .D(n898), .Y(n623) );
  ao22d1_hd U1458 ( .A(n910), .B(n874), .C(a_m[18]), .D(n905), .Y(n650) );
  ao22d1_hd U1459 ( .A(a_m[19]), .B(n874), .C(a_m[18]), .D(n875), .Y(n618) );
  ao22d1_hd U1460 ( .A(n951), .B(n511), .C(n1073), .D(n525), .Y(n617) );
  oa211d1_hd U1461 ( .A(n862), .B(n621), .C(n620), .D(n619), .Y(n622) );
  scg4d1_hd U1462 ( .A(n487), .B(n1067), .C(n953), .D(n510), .E(n1073), .F(
        n409), .G(n949), .H(n561), .Y(n624) );
  scg4d1_hd U1463 ( .A(n486), .B(n560), .C(n959), .D(n509), .E(n648), .F(n449), 
        .G(n1067), .H(b_m[21]), .Y(n625) );
  scg4d1_hd U1464 ( .A(n955), .B(n559), .C(n964), .D(n512), .E(n1074), .F(n451), .G(n1067), .H(n961), .Y(n626) );
  scg4d1_hd U1465 ( .A(b_m[20]), .B(n562), .C(n969), .D(n511), .E(n1074), .F(
        n447), .G(n1067), .H(n965), .Y(n627) );
  scg4d1_hd U1466 ( .A(b_m[19]), .B(n561), .C(n974), .D(n510), .E(n648), .F(
        n445), .G(n646), .H(n970), .Y(n628) );
  scg4d1_hd U1467 ( .A(b_m[18]), .B(n560), .C(n979), .D(n509), .E(n648), .F(
        n443), .G(n1067), .H(n976), .Y(n629) );
  scg4d1_hd U1468 ( .A(b_m[17]), .B(n559), .C(n984), .D(n512), .E(n648), .F(
        n441), .G(n646), .H(n981), .Y(n630) );
  scg4d1_hd U1469 ( .A(b_m[16]), .B(n562), .C(b_m[14]), .D(n511), .E(n1071), 
        .F(n437), .G(n1070), .H(n985), .Y(n631) );
  scg4d1_hd U1470 ( .A(b_m[15]), .B(n561), .C(n995), .D(n510), .E(n1072), .F(
        n439), .G(n1070), .H(n991), .Y(n632) );
  scg4d1_hd U1471 ( .A(n989), .B(n560), .C(n1000), .D(n509), .E(n1072), .F(
        n433), .G(n1070), .H(n997), .Y(n633) );
  scg4d1_hd U1472 ( .A(n996), .B(n559), .C(n1005), .D(n512), .E(n1072), .F(
        n435), .G(n1070), .H(n1002), .Y(n634) );
  scg4d1_hd U1473 ( .A(n1001), .B(n562), .C(n1010), .D(n511), .E(n1072), .F(
        n431), .G(n1068), .H(n1008), .Y(n635) );
  scg4d1_hd U1474 ( .A(n1006), .B(n561), .C(n1015), .D(n510), .E(n1072), .F(
        n429), .G(n1068), .H(n1013), .Y(n636) );
  scg4d1_hd U1475 ( .A(n1011), .B(n560), .C(n1019), .D(n509), .E(n1071), .F(
        n425), .G(n1068), .H(n1017), .Y(n637) );
  scg4d1_hd U1476 ( .A(n1016), .B(n559), .C(n1024), .D(n512), .E(n1071), .F(
        n427), .G(n1068), .H(n1022), .Y(n638) );
  scg4d1_hd U1477 ( .A(n1020), .B(n562), .C(n1029), .D(n511), .E(n1071), .F(
        n421), .G(n1068), .H(n1025), .Y(n639) );
  scg4d1_hd U1478 ( .A(b_m[7]), .B(n561), .C(n1034), .D(n510), .E(n1072), .F(
        n423), .G(n1068), .H(n1030), .Y(n640) );
  scg4d1_hd U1479 ( .A(n1033), .B(n560), .C(n1039), .D(n509), .E(n1071), .F(
        n419), .G(n1069), .H(n1036), .Y(n641) );
  scg4d1_hd U1480 ( .A(b_m[5]), .B(n559), .C(n1044), .D(n512), .E(n1074), .F(
        n417), .G(n1069), .H(n1041), .Y(n642) );
  scg4d1_hd U1481 ( .A(b_m[4]), .B(n562), .C(n1049), .D(n511), .E(n1073), .F(
        n415), .G(n1069), .H(n1046), .Y(n643) );
  scg4d1_hd U1482 ( .A(n1048), .B(n561), .C(n1055), .D(n510), .E(n1074), .F(
        n413), .G(n1069), .H(n1051), .Y(n644) );
  scg4d1_hd U1483 ( .A(b_m[2]), .B(n560), .C(n579), .D(n509), .E(n1073), .F(
        n411), .G(n1069), .H(n1056), .Y(n645) );
  scg5d1_hd U1484 ( .A(n1073), .B(n455), .C(n1057), .D(n559), .E(n1067), .F(
        n484), .Y(n649) );
  nr2d1_hd U1485 ( .A(n465), .B(n650), .Y(n651) );
  ao22d1_hd U1486 ( .A(n910), .B(a_m[16]), .C(n873), .D(n905), .Y(n658) );
  ao22d1_hd U1487 ( .A(n917), .B(n872), .C(a_m[15]), .D(n912), .Y(n685) );
  ao22d1_hd U1488 ( .A(a_m[16]), .B(n872), .C(a_m[15]), .D(n873), .Y(n653) );
  ao22d1_hd U1489 ( .A(n951), .B(n507), .C(n1081), .D(n525), .Y(n652) );
  oa211d1_hd U1490 ( .A(n862), .B(n656), .C(n655), .D(n654), .Y(n657) );
  scg4d1_hd U1491 ( .A(b_m[22]), .B(n1075), .C(n954), .D(n506), .E(n1081), .F(
        mult_x_1_n641), .G(n949), .H(n557), .Y(n659) );
  scg4d1_hd U1492 ( .A(n488), .B(n556), .C(n959), .D(n505), .E(n683), .F(
        mult_x_1_n642), .G(n1075), .H(b_m[21]), .Y(n660) );
  scg4d1_hd U1493 ( .A(n955), .B(n555), .C(n964), .D(n508), .E(n1082), .F(
        mult_x_1_n643), .G(n1075), .H(n963), .Y(n661) );
  scg4d1_hd U1494 ( .A(n963), .B(n558), .C(n969), .D(n507), .E(n1082), .F(
        mult_x_1_n644), .G(n1075), .H(n965), .Y(n662) );
  scg4d1_hd U1495 ( .A(n968), .B(n557), .C(n974), .D(n506), .E(n683), .F(
        mult_x_1_n645), .G(n1076), .H(n970), .Y(n663) );
  scg4d1_hd U1496 ( .A(n973), .B(n556), .C(n979), .D(n505), .E(n683), .F(
        mult_x_1_n646), .G(n1075), .H(n975), .Y(n664) );
  scg4d1_hd U1497 ( .A(n975), .B(n555), .C(n984), .D(n508), .E(n683), .F(
        mult_x_1_n647), .G(n1076), .H(n980), .Y(n665) );
  scg4d1_hd U1498 ( .A(n980), .B(n558), .C(b_m[14]), .D(n507), .E(n1079), .F(
        mult_x_1_n648), .G(n1076), .H(n985), .Y(n666) );
  scg4d1_hd U1499 ( .A(n988), .B(n557), .C(n995), .D(n506), .E(n1080), .F(
        mult_x_1_n649), .G(n1076), .H(n990), .Y(n667) );
  scg4d1_hd U1500 ( .A(n990), .B(n556), .C(n1000), .D(n505), .E(n1080), .F(
        mult_x_1_n650), .G(n1076), .H(n997), .Y(n668) );
  scg4d1_hd U1501 ( .A(n996), .B(n555), .C(n1005), .D(n508), .E(n1080), .F(
        mult_x_1_n651), .G(n1076), .H(n1002), .Y(n669) );
  scg4d1_hd U1502 ( .A(n1001), .B(n558), .C(n1010), .D(n507), .E(n1080), .F(
        mult_x_1_n652), .G(n681), .H(n1007), .Y(n670) );
  scg4d1_hd U1503 ( .A(n1007), .B(n557), .C(n1015), .D(n506), .E(n1080), .F(
        mult_x_1_n653), .G(n681), .H(n1012), .Y(n671) );
  scg4d1_hd U1504 ( .A(n1012), .B(n556), .C(n1019), .D(n505), .E(n1079), .F(
        mult_x_1_n654), .G(n1078), .H(n1017), .Y(n672) );
  scg4d1_hd U1505 ( .A(n1016), .B(n555), .C(n1024), .D(n508), .E(n1079), .F(
        mult_x_1_n655), .G(n681), .H(n1021), .Y(n673) );
  scg4d1_hd U1506 ( .A(n1021), .B(n558), .C(n1029), .D(n507), .E(n1079), .F(
        mult_x_1_n656), .G(n1078), .H(n1025), .Y(n674) );
  scg4d1_hd U1507 ( .A(n1028), .B(n557), .C(n1034), .D(n506), .E(n1080), .F(
        mult_x_1_n657), .G(n1078), .H(n1030), .Y(n675) );
  scg4d1_hd U1508 ( .A(b_m[6]), .B(n556), .C(n1039), .D(n505), .E(n1079), .F(
        mult_x_1_n658), .G(n1077), .H(n1035), .Y(n676) );
  scg4d1_hd U1509 ( .A(n1035), .B(n555), .C(n1044), .D(n508), .E(n1082), .F(
        mult_x_1_n659), .G(n1077), .H(n1040), .Y(n677) );
  scg4d1_hd U1510 ( .A(n1040), .B(n558), .C(n1049), .D(n507), .E(n1081), .F(
        mult_x_1_n660), .G(n1077), .H(n1045), .Y(n678) );
  scg4d1_hd U1511 ( .A(n1045), .B(n557), .C(n1055), .D(n506), .E(n1082), .F(
        mult_x_1_n661), .G(n1077), .H(n1050), .Y(n679) );
  scg4d1_hd U1512 ( .A(n1050), .B(n556), .C(n483), .D(n505), .E(n1081), .F(
        mult_x_1_n662), .G(n1077), .H(n1056), .Y(n680) );
  scg5d1_hd U1513 ( .A(n1081), .B(mult_x_1_n663), .C(n1057), .D(n555), .E(
        n1075), .F(n579), .Y(n684) );
  nr2d1_hd U1514 ( .A(n465), .B(n685), .Y(n686) );
  ao22d1_hd U1515 ( .A(n917), .B(a_m[13]), .C(n871), .D(n912), .Y(n693) );
  ao22d1_hd U1516 ( .A(n924), .B(n870), .C(a_m[12]), .D(n919), .Y(n720) );
  ao22d1_hd U1517 ( .A(a_m[13]), .B(n870), .C(a_m[12]), .D(n871), .Y(n688) );
  ao22d1_hd U1518 ( .A(n951), .B(n515), .C(n1089), .D(mult_x_1_n639), .Y(n687)
         );
  oa211d1_hd U1519 ( .A(n862), .B(n691), .C(n690), .D(n689), .Y(n692) );
  scg4d1_hd U1520 ( .A(n487), .B(n1083), .C(n954), .D(n514), .E(n1089), .F(
        n409), .G(n949), .H(n565), .Y(n694) );
  scg4d1_hd U1521 ( .A(n486), .B(n564), .C(n959), .D(n513), .E(n718), .F(n449), 
        .G(n1083), .H(n958), .Y(n695) );
  scg4d1_hd U1522 ( .A(n955), .B(n563), .C(n964), .D(n516), .E(n1090), .F(n451), .G(n1083), .H(n963), .Y(n696) );
  scg4d1_hd U1523 ( .A(n960), .B(n566), .C(n969), .D(n515), .E(n1090), .F(n447), .G(n1083), .H(n965), .Y(n697) );
  scg4d1_hd U1524 ( .A(n968), .B(n565), .C(n974), .D(n514), .E(n718), .F(n445), 
        .G(n1084), .H(n970), .Y(n698) );
  scg4d1_hd U1525 ( .A(n973), .B(n564), .C(n979), .D(n513), .E(n718), .F(n443), 
        .G(n1083), .H(n975), .Y(n699) );
  scg4d1_hd U1526 ( .A(n978), .B(n563), .C(n984), .D(n516), .E(n718), .F(n441), 
        .G(n1084), .H(n980), .Y(n700) );
  scg4d1_hd U1527 ( .A(n983), .B(n566), .C(b_m[14]), .D(n515), .E(n1087), .F(
        n437), .G(n1084), .H(n985), .Y(n701) );
  scg4d1_hd U1528 ( .A(n988), .B(n565), .C(n995), .D(n514), .E(n1088), .F(n439), .G(n1084), .H(n990), .Y(n702) );
  scg4d1_hd U1529 ( .A(n989), .B(n564), .C(n1000), .D(n513), .E(n1088), .F(
        n433), .G(n1084), .H(n997), .Y(n703) );
  scg4d1_hd U1530 ( .A(n996), .B(n563), .C(n1005), .D(n516), .E(n1088), .F(
        n435), .G(n1084), .H(n1002), .Y(n704) );
  scg4d1_hd U1531 ( .A(n1001), .B(n566), .C(n1010), .D(n515), .E(n1088), .F(
        n431), .G(n716), .H(n1007), .Y(n705) );
  scg4d1_hd U1532 ( .A(n1006), .B(n565), .C(n1015), .D(n514), .E(n1088), .F(
        n429), .G(n716), .H(n1012), .Y(n706) );
  scg4d1_hd U1533 ( .A(n1011), .B(n564), .C(n1019), .D(n513), .E(n1087), .F(
        n425), .G(n1086), .H(n1017), .Y(n707) );
  scg4d1_hd U1534 ( .A(n1016), .B(n563), .C(n1024), .D(n516), .E(n1087), .F(
        n427), .G(n716), .H(n1021), .Y(n708) );
  scg4d1_hd U1535 ( .A(n1020), .B(n566), .C(n1029), .D(n515), .E(n1087), .F(
        n421), .G(n1086), .H(n1025), .Y(n709) );
  scg4d1_hd U1536 ( .A(n1028), .B(n565), .C(n1034), .D(n514), .E(n1088), .F(
        n423), .G(n1086), .H(n1030), .Y(n710) );
  scg4d1_hd U1537 ( .A(b_m[6]), .B(n564), .C(n1039), .D(n513), .E(n1087), .F(
        n419), .G(n1085), .H(n1035), .Y(n711) );
  scg4d1_hd U1538 ( .A(n1038), .B(n563), .C(n1044), .D(n516), .E(n1090), .F(
        n417), .G(n1085), .H(n1040), .Y(n712) );
  scg4d1_hd U1539 ( .A(n1043), .B(n566), .C(n1049), .D(n515), .E(n1089), .F(
        n415), .G(n1085), .H(n1045), .Y(n713) );
  scg4d1_hd U1540 ( .A(b_m[3]), .B(n565), .C(n1055), .D(n514), .E(n1090), .F(
        n413), .G(n1085), .H(n1050), .Y(n714) );
  scg4d1_hd U1541 ( .A(n1053), .B(n564), .C(b_m[0]), .D(n513), .E(n1089), .F(
        n411), .G(n1085), .H(n1058), .Y(n715) );
  scg5d1_hd U1542 ( .A(n1089), .B(n455), .C(n1054), .D(n563), .E(n1083), .F(
        n484), .Y(n719) );
  nr2d1_hd U1543 ( .A(n465), .B(n720), .Y(n721) );
  ao22d1_hd U1544 ( .A(n924), .B(a_m[10]), .C(n869), .D(n919), .Y(n728) );
  ao22d1_hd U1545 ( .A(n931), .B(n868), .C(a_m[9]), .D(n925), .Y(n755) );
  ao22d1_hd U1546 ( .A(a_m[10]), .B(n868), .C(a_m[9]), .D(n869), .Y(n723) );
  ao22d1_hd U1547 ( .A(n951), .B(n503), .C(n1097), .D(mult_x_1_n639), .Y(n722)
         );
  oa211d1_hd U1548 ( .A(n862), .B(n726), .C(n725), .D(n724), .Y(n727) );
  scg4d1_hd U1549 ( .A(b_m[22]), .B(n1091), .C(n954), .D(n502), .E(n1097), .F(
        mult_x_1_n641), .G(n948), .H(n553), .Y(n729) );
  scg4d1_hd U1550 ( .A(n488), .B(n552), .C(n960), .D(n501), .E(n753), .F(
        mult_x_1_n642), .G(n1091), .H(n958), .Y(n730) );
  scg4d1_hd U1551 ( .A(n955), .B(n551), .C(n964), .D(n504), .E(n1098), .F(
        mult_x_1_n643), .G(n1091), .H(n963), .Y(n731) );
  scg4d1_hd U1552 ( .A(n960), .B(n554), .C(n969), .D(n503), .E(n1098), .F(
        mult_x_1_n644), .G(n1091), .H(n965), .Y(n732) );
  scg4d1_hd U1553 ( .A(n968), .B(n553), .C(n974), .D(n502), .E(n753), .F(
        mult_x_1_n645), .G(n751), .H(n970), .Y(n733) );
  scg4d1_hd U1554 ( .A(n973), .B(n552), .C(n979), .D(n501), .E(n753), .F(
        mult_x_1_n646), .G(n1091), .H(n976), .Y(n734) );
  scg4d1_hd U1555 ( .A(n978), .B(n551), .C(n984), .D(n504), .E(n753), .F(
        mult_x_1_n647), .G(n751), .H(n981), .Y(n735) );
  scg4d1_hd U1556 ( .A(n983), .B(n554), .C(n992), .D(n503), .E(n1095), .F(
        mult_x_1_n648), .G(n1094), .H(n985), .Y(n736) );
  scg4d1_hd U1557 ( .A(n988), .B(n553), .C(n995), .D(n502), .E(n1096), .F(
        mult_x_1_n649), .G(n1094), .H(n991), .Y(n737) );
  scg4d1_hd U1558 ( .A(n989), .B(n552), .C(n1000), .D(n501), .E(n1096), .F(
        mult_x_1_n650), .G(n1094), .H(n997), .Y(n738) );
  scg4d1_hd U1559 ( .A(n996), .B(n551), .C(n1005), .D(n504), .E(n1096), .F(
        mult_x_1_n651), .G(n1094), .H(n1002), .Y(n739) );
  scg4d1_hd U1560 ( .A(n1001), .B(n554), .C(n1010), .D(n503), .E(n1096), .F(
        mult_x_1_n652), .G(n1092), .H(n1008), .Y(n740) );
  scg4d1_hd U1561 ( .A(n1006), .B(n553), .C(n1015), .D(n502), .E(n1096), .F(
        mult_x_1_n653), .G(n1092), .H(n1013), .Y(n741) );
  scg4d1_hd U1562 ( .A(n1011), .B(n552), .C(n1019), .D(n501), .E(n1095), .F(
        mult_x_1_n654), .G(n1092), .H(n1017), .Y(n742) );
  scg4d1_hd U1563 ( .A(n1016), .B(n551), .C(n1024), .D(n504), .E(n1095), .F(
        mult_x_1_n655), .G(n1092), .H(n1022), .Y(n743) );
  scg4d1_hd U1564 ( .A(n1020), .B(n554), .C(n1029), .D(n503), .E(n1095), .F(
        mult_x_1_n656), .G(n1092), .H(n1025), .Y(n744) );
  scg4d1_hd U1565 ( .A(n1028), .B(n553), .C(n1034), .D(n502), .E(n1096), .F(
        mult_x_1_n657), .G(n1092), .H(n1030), .Y(n745) );
  scg4d1_hd U1566 ( .A(b_m[6]), .B(n552), .C(n1039), .D(n501), .E(n1098), .F(
        mult_x_1_n658), .G(n1093), .H(n1036), .Y(n746) );
  scg4d1_hd U1567 ( .A(n1038), .B(n551), .C(n1044), .D(n504), .E(n1095), .F(
        mult_x_1_n659), .G(n1093), .H(n1041), .Y(n747) );
  scg4d1_hd U1568 ( .A(n1043), .B(n554), .C(n1049), .D(n503), .E(n1097), .F(
        mult_x_1_n660), .G(n1093), .H(n1046), .Y(n748) );
  scg4d1_hd U1569 ( .A(b_m[3]), .B(n553), .C(n1058), .D(n502), .E(n1098), .F(
        mult_x_1_n661), .G(n1093), .H(n1051), .Y(n749) );
  scg4d1_hd U1570 ( .A(n1053), .B(n552), .C(n483), .D(n501), .E(n1097), .F(
        mult_x_1_n662), .G(n1093), .H(n1058), .Y(n750) );
  scg5d1_hd U1571 ( .A(n1097), .B(mult_x_1_n663), .C(n1054), .D(n551), .E(
        n1091), .F(n484), .Y(n754) );
  nr2d1_hd U1572 ( .A(n465), .B(n755), .Y(n756) );
  ao22d1_hd U1573 ( .A(n931), .B(a_m[7]), .C(n867), .D(n925), .Y(n763) );
  ao22d1_hd U1574 ( .A(a_m[7]), .B(n866), .C(a_m[6]), .D(n867), .Y(n758) );
  ao22d1_hd U1575 ( .A(n952), .B(n499), .C(n1106), .D(mult_x_1_n639), .Y(n757)
         );
  oa211d1_hd U1576 ( .A(n862), .B(n761), .C(n760), .D(n759), .Y(n762) );
  scg4d1_hd U1577 ( .A(n487), .B(n1099), .C(n954), .D(n498), .E(n1106), .F(
        n409), .G(n949), .H(n549), .Y(n764) );
  scg4d1_hd U1578 ( .A(n486), .B(n548), .C(n959), .D(n497), .E(n1104), .F(n449), .G(n1099), .H(n958), .Y(n765) );
  scg4d1_hd U1579 ( .A(n954), .B(n547), .C(n967), .D(n500), .E(n788), .F(n451), 
        .G(n1099), .H(n961), .Y(n766) );
  scg4d1_hd U1580 ( .A(n960), .B(n550), .C(n972), .D(n499), .E(n788), .F(n447), 
        .G(n1099), .H(n966), .Y(n767) );
  scg4d1_hd U1581 ( .A(n968), .B(n549), .C(n974), .D(n498), .E(n1104), .F(n445), .G(n1100), .H(n971), .Y(n768) );
  scg4d1_hd U1582 ( .A(n973), .B(n548), .C(n979), .D(n497), .E(n1104), .F(n443), .G(n1099), .H(n975), .Y(n769) );
  scg4d1_hd U1583 ( .A(n978), .B(n547), .C(n987), .D(n500), .E(n1104), .F(n441), .G(n1100), .H(n980), .Y(n770) );
  scg4d1_hd U1584 ( .A(n983), .B(n550), .C(n992), .D(n499), .E(n1104), .F(n437), .G(n1100), .H(n986), .Y(n771) );
  scg4d1_hd U1585 ( .A(n988), .B(n549), .C(n994), .D(n498), .E(n1105), .F(n439), .G(n1100), .H(n990), .Y(n772) );
  scg4d1_hd U1586 ( .A(n989), .B(n548), .C(n999), .D(n497), .E(n1105), .F(n433), .G(n1100), .H(n998), .Y(n773) );
  scg4d1_hd U1587 ( .A(n996), .B(n547), .C(n1005), .D(n500), .E(n1105), .F(
        n435), .G(n1100), .H(n1003), .Y(n774) );
  scg4d1_hd U1588 ( .A(n1001), .B(n550), .C(n1010), .D(n499), .E(n1105), .F(
        n431), .G(n786), .H(n1007), .Y(n775) );
  scg4d1_hd U1589 ( .A(n1006), .B(n549), .C(n1014), .D(n498), .E(n1105), .F(
        n429), .G(n786), .H(n1012), .Y(n776) );
  scg4d1_hd U1590 ( .A(n1011), .B(n548), .C(n1019), .D(n497), .E(n1103), .F(
        n425), .G(n1102), .H(n1018), .Y(n777) );
  scg4d1_hd U1591 ( .A(n1016), .B(n547), .C(n1027), .D(n500), .E(n1103), .F(
        n427), .G(n786), .H(n1021), .Y(n778) );
  scg4d1_hd U1592 ( .A(n1020), .B(n550), .C(n1032), .D(n499), .E(n1103), .F(
        n421), .G(n1102), .H(n1026), .Y(n779) );
  scg4d1_hd U1593 ( .A(n1028), .B(n549), .C(n1034), .D(n498), .E(n1105), .F(
        n423), .G(n1102), .H(n1031), .Y(n780) );
  scg4d1_hd U1594 ( .A(n1033), .B(n548), .C(n1039), .D(n497), .E(n788), .F(
        n419), .G(n1101), .H(n1035), .Y(n781) );
  scg4d1_hd U1595 ( .A(n1038), .B(n547), .C(n1044), .D(n500), .E(n1103), .F(
        n417), .G(n1101), .H(n1040), .Y(n782) );
  scg4d1_hd U1596 ( .A(n1043), .B(n550), .C(n1049), .D(n499), .E(n1106), .F(
        n415), .G(n1101), .H(n1045), .Y(n783) );
  scg4d1_hd U1597 ( .A(b_m[3]), .B(n549), .C(n1055), .D(n498), .E(n788), .F(
        n413), .G(n1101), .H(n1050), .Y(n784) );
  scg4d1_hd U1598 ( .A(n1053), .B(n548), .C(b_m[0]), .D(n497), .E(n1106), .F(
        n411), .G(n1101), .H(n1058), .Y(n785) );
  scg5d1_hd U1599 ( .A(n1106), .B(n455), .C(n1054), .D(n547), .E(n1099), .F(
        n484), .Y(n789) );
  nr2d1_hd U1600 ( .A(n464), .B(n790), .Y(n791) );
  ao22d1_hd U1601 ( .A(n938), .B(a_m[4]), .C(n865), .D(n933), .Y(n798) );
  ao22d1_hd U1602 ( .A(a_m[4]), .B(n864), .C(a_m[3]), .D(n865), .Y(n793) );
  ao22d1_hd U1603 ( .A(n952), .B(n495), .C(n1114), .D(mult_x_1_n639), .Y(n792)
         );
  oa211d1_hd U1604 ( .A(n862), .B(n796), .C(n795), .D(n794), .Y(n797) );
  scg4d1_hd U1605 ( .A(b_m[22]), .B(n1108), .C(n953), .D(n494), .E(n1114), .F(
        n409), .G(n949), .H(n545), .Y(n799) );
  scg4d1_hd U1606 ( .A(n486), .B(n544), .C(n959), .D(n493), .E(n1111), .F(n449), .G(n1108), .H(n958), .Y(n800) );
  scg4d1_hd U1607 ( .A(n954), .B(n543), .C(n967), .D(n496), .E(n823), .F(n451), 
        .G(n1108), .H(n961), .Y(n801) );
  scg4d1_hd U1608 ( .A(n960), .B(n546), .C(n972), .D(n495), .E(n823), .F(n447), 
        .G(n1108), .H(n966), .Y(n802) );
  scg4d1_hd U1609 ( .A(n964), .B(n545), .C(n977), .D(n494), .E(n1111), .F(n445), .G(n821), .H(n971), .Y(n803) );
  scg4d1_hd U1610 ( .A(n969), .B(n544), .C(n982), .D(n493), .E(n1111), .F(n443), .G(n1108), .H(n976), .Y(n804) );
  scg4d1_hd U1611 ( .A(n978), .B(n543), .C(n987), .D(n496), .E(n1111), .F(n441), .G(n821), .H(n981), .Y(n805) );
  scg4d1_hd U1612 ( .A(n983), .B(n546), .C(n992), .D(n495), .E(n1111), .F(n437), .G(n821), .H(n986), .Y(n806) );
  scg4d1_hd U1613 ( .A(n984), .B(n545), .C(n994), .D(n494), .E(n1112), .F(n439), .G(n1107), .H(n991), .Y(n807) );
  scg4d1_hd U1614 ( .A(n989), .B(n544), .C(n999), .D(n493), .E(n1112), .F(n433), .G(n1107), .H(n998), .Y(n808) );
  scg4d1_hd U1615 ( .A(n995), .B(n543), .C(n1004), .D(n496), .E(n1112), .F(
        n435), .G(n1107), .H(n1003), .Y(n809) );
  scg4d1_hd U1616 ( .A(n1000), .B(n546), .C(n1009), .D(n495), .E(n1112), .F(
        n431), .G(n1109), .H(n1008), .Y(n810) );
  scg4d1_hd U1617 ( .A(n1006), .B(n545), .C(n1014), .D(n494), .E(n1112), .F(
        n429), .G(n1109), .H(n1013), .Y(n811) );
  scg4d1_hd U1618 ( .A(n1011), .B(n544), .C(n1023), .D(n493), .E(n1113), .F(
        n425), .G(n1109), .H(n1018), .Y(n812) );
  scg4d1_hd U1619 ( .A(n1015), .B(n543), .C(n1027), .D(n496), .E(n1113), .F(
        n427), .G(n1109), .H(n1022), .Y(n813) );
  scg4d1_hd U1620 ( .A(n1020), .B(n546), .C(n1032), .D(n495), .E(n1113), .F(
        n421), .G(n1109), .H(n1026), .Y(n814) );
  scg4d1_hd U1621 ( .A(n1024), .B(n545), .C(n1037), .D(n494), .E(n1112), .F(
        n423), .G(n1109), .H(n1031), .Y(n815) );
  scg4d1_hd U1622 ( .A(n1029), .B(n544), .C(n1042), .D(n493), .E(n1113), .F(
        n419), .G(n1110), .H(n1036), .Y(n816) );
  scg4d1_hd U1623 ( .A(n1038), .B(n543), .C(n1047), .D(n496), .E(n1113), .F(
        n417), .G(n1110), .H(n1041), .Y(n817) );
  scg4d1_hd U1624 ( .A(n1043), .B(n546), .C(n1052), .D(n495), .E(n1114), .F(
        n415), .G(n1110), .H(n1046), .Y(n818) );
  scg4d1_hd U1625 ( .A(n1048), .B(n545), .C(n1055), .D(n494), .E(n1113), .F(
        n413), .G(n1110), .H(n1051), .Y(n819) );
  scg4d1_hd U1626 ( .A(n1053), .B(n544), .C(n483), .D(n493), .E(n1114), .F(
        n411), .G(n1110), .H(n1056), .Y(n820) );
  scg5d1_hd U1627 ( .A(n1114), .B(n455), .C(n1054), .D(n543), .E(n1108), .F(
        b_m[0]), .Y(n824) );
  nr2d1_hd U1628 ( .A(n464), .B(n825), .Y(n826) );
  ao22d1_hd U1629 ( .A(n952), .B(n1117), .C(mult_x_1_n639), .D(n857), .Y(n827)
         );
  scg15d1_hd U1630 ( .A(n487), .B(n853), .C(n829), .D(n828), .Y(n830) );
  scg4d1_hd U1631 ( .A(b_m[22]), .B(n1119), .C(n953), .D(n1118), .E(n1123), 
        .F(n409), .G(n949), .H(n541), .Y(n832) );
  scg4d1_hd U1632 ( .A(n488), .B(n540), .C(n959), .D(n1118), .E(n1123), .F(
        n449), .G(n1119), .H(n956), .Y(n833) );
  scg4d1_hd U1633 ( .A(n955), .B(n539), .C(n964), .D(n1118), .E(n1123), .F(
        n451), .G(n1119), .H(n961), .Y(n834) );
  scg4d1_hd U1634 ( .A(n960), .B(n542), .C(n969), .D(n1118), .E(n1123), .F(
        n447), .G(n1119), .H(n966), .Y(n835) );
  scg4d1_hd U1635 ( .A(n965), .B(n541), .C(n974), .D(n853), .E(n1126), .F(n445), .G(n855), .H(n971), .Y(n836) );
  scg4d1_hd U1636 ( .A(n970), .B(n540), .C(n979), .D(n1115), .E(n1126), .F(
        n443), .G(n1119), .H(n976), .Y(n837) );
  scg4d1_hd U1637 ( .A(n975), .B(n539), .C(n984), .D(n1115), .E(n1126), .F(
        n441), .G(n855), .H(n981), .Y(n838) );
  scg4d1_hd U1638 ( .A(n980), .B(n542), .C(n992), .D(n1115), .E(n1126), .F(
        n437), .G(n1122), .H(n986), .Y(n839) );
  scg4d1_hd U1639 ( .A(n985), .B(n541), .C(n995), .D(n1115), .E(n1126), .F(
        n439), .G(n1122), .H(n991), .Y(n840) );
  scg4d1_hd U1640 ( .A(n990), .B(n540), .C(n1000), .D(n1115), .E(n1126), .F(
        n433), .G(n1122), .H(n998), .Y(n841) );
  scg4d1_hd U1641 ( .A(n997), .B(n539), .C(n1005), .D(n1116), .E(n1125), .F(
        n435), .G(n1122), .H(n1003), .Y(n842) );
  scg4d1_hd U1642 ( .A(n1002), .B(n542), .C(n1010), .D(n1116), .E(n1125), .F(
        n431), .G(n1120), .H(n1008), .Y(n843) );
  scg4d1_hd U1643 ( .A(n1007), .B(n541), .C(n1015), .D(n1116), .E(n1124), .F(
        n429), .G(n1120), .H(n1013), .Y(n844) );
  scg4d1_hd U1644 ( .A(n1012), .B(n540), .C(n1019), .D(n1116), .E(n1124), .F(
        n425), .G(n1120), .H(n1018), .Y(n845) );
  scg4d1_hd U1645 ( .A(n1017), .B(n539), .C(n1024), .D(n1116), .E(n1124), .F(
        n427), .G(n1120), .H(n1022), .Y(n846) );
  scg4d1_hd U1646 ( .A(n1021), .B(n542), .C(n1029), .D(n1116), .E(n1124), .F(
        n421), .G(n1120), .H(n1026), .Y(n847) );
  scg4d1_hd U1647 ( .A(n1025), .B(n541), .C(n1034), .D(n1117), .E(n1125), .F(
        n423), .G(n1120), .H(n1031), .Y(n848) );
  scg4d1_hd U1648 ( .A(n1030), .B(n540), .C(n1039), .D(n1117), .E(n857), .F(
        n419), .G(n1121), .H(n1036), .Y(n849) );
  scg4d1_hd U1649 ( .A(n1035), .B(n539), .C(n1044), .D(n1117), .E(n857), .F(
        n417), .G(n1121), .H(n1041), .Y(n850) );
  scg4d1_hd U1650 ( .A(n1040), .B(n542), .C(n1049), .D(n1117), .E(n857), .F(
        n415), .G(n1121), .H(n1046), .Y(n851) );
  scg4d1_hd U1651 ( .A(n1045), .B(n541), .C(n1055), .D(n1117), .E(n1124), .F(
        n413), .G(n1121), .H(n1051), .Y(n852) );
  scg4d1_hd U1652 ( .A(n1050), .B(n540), .C(b_m[0]), .D(n1115), .E(n1125), .F(
        n411), .G(n1121), .H(n1056), .Y(n854) );
  scg5d1_hd U1653 ( .A(n455), .B(n1125), .C(n1054), .D(n539), .E(n1119), .F(
        n484), .Y(n858) );
  nr2d1_hd U1654 ( .A(n464), .B(n387), .Y(n859) );
  oa211d1_hd U1655 ( .A(n946), .B(n956), .C(n892), .D(n860), .Y(n861) );
  ivd1_hd U1656 ( .A(a_m[10]), .Y(n869) );
  ivd1_hd U1657 ( .A(a_m[13]), .Y(n871) );
  ivd1_hd U1658 ( .A(a_m[16]), .Y(n873) );
  ivd1_hd U1659 ( .A(a_m[18]), .Y(n874) );
  ivd1_hd U1660 ( .A(a_m[19]), .Y(n875) );
  ivd1_hd U1661 ( .A(mult_x_1_n315), .Y(n878) );
  ivd1_hd U1662 ( .A(mult_x_1_n302), .Y(n879) );
  ivd1_hd U1663 ( .A(mult_x_1_n277), .Y(n880) );
  ivd1_hd U1664 ( .A(mult_x_1_n245), .Y(n881) );
  ivd1_hd U1665 ( .A(mult_x_1_n236), .Y(n882) );
  ivd1_hd U1666 ( .A(mult_x_1_n219), .Y(n883) );
  ivd1_hd U1667 ( .A(mult_x_1_n199), .Y(n884) );
  ivd1_hd U1668 ( .A(mult_x_1_n194), .Y(n885) );
  nr4d1_hd U1669 ( .A(a_e[3]), .B(a_e[5]), .C(a_e[6]), .D(n1223), .Y(n1239) );
  nr4d1_hd U1670 ( .A(a_m[6]), .B(a_m[10]), .C(a_m[14]), .D(n388), .Y(n1230)
         );
  nr4d1_hd U1671 ( .A(a_m[13]), .B(a_m[17]), .C(a_m[12]), .D(a_m[16]), .Y(
        n1229) );
  nr4d1_hd U1672 ( .A(a_m[2]), .B(a_m[15]), .C(a_m[4]), .D(a_m[1]), .Y(n1227)
         );
  nr4d1_hd U1673 ( .A(a_m[20]), .B(a_m[21]), .C(a_m[22]), .D(a_m[19]), .Y(
        n1226) );
  nr4d1_hd U1674 ( .A(a_m[23]), .B(a_m[3]), .C(a_m[5]), .D(a_m[11]), .Y(n1225)
         );
  nr4d1_hd U1675 ( .A(a_m[18]), .B(a_m[7]), .C(a_m[8]), .D(a_m[9]), .Y(n1224)
         );
  nd3d1_hd U1676 ( .A(n1230), .B(n1229), .C(n1228), .Y(n1247) );
  nr4d1_hd U1677 ( .A(b_e[3]), .B(b_e[5]), .C(b_e[6]), .D(n1231), .Y(n1241) );
  nr4d1_hd U1678 ( .A(b_m[11]), .B(b_m[10]), .C(b_m[14]), .D(n484), .Y(n1238)
         );
  nr4d1_hd U1679 ( .A(b_m[13]), .B(b_m[17]), .C(b_m[12]), .D(b_m[16]), .Y(
        n1237) );
  nr4d1_hd U1680 ( .A(b_m[2]), .B(b_m[15]), .C(b_m[4]), .D(b_m[1]), .Y(n1235)
         );
  nr4d1_hd U1681 ( .A(b_m[20]), .B(b_m[21]), .C(b_m[22]), .D(b_m[19]), .Y(
        n1234) );
  nr4d1_hd U1682 ( .A(b_m[23]), .B(b_m[6]), .C(b_m[3]), .D(b_m[5]), .Y(n1233)
         );
  nr4d1_hd U1683 ( .A(b_m[18]), .B(b_m[7]), .C(b_m[8]), .D(b_m[9]), .Y(n1232)
         );
  nd3d1_hd U1684 ( .A(n1238), .B(n1237), .C(n1236), .Y(n1244) );
  ivd1_hd U1685 ( .A(n1239), .Y(n1240) );
  ivd1_hd U1686 ( .A(n1241), .Y(n1242) );
  oa21d1_hd U1687 ( .A(n1245), .B(n1244), .C(n1243), .Y(n1250) );
  oa21d1_hd U1688 ( .A(n1248), .B(n1247), .C(n1246), .Y(n1249) );
  ao21d1_hd U1689 ( .A(n1250), .B(n1249), .C(n1338), .Y(n1288) );
  ao21d1_hd U1690 ( .A(n1161), .B(z[22]), .C(n1288), .Y(n1251) );
  oa21d1_hd U1691 ( .A(n1374), .B(n1252), .C(n1251), .Y(n238) );
  nr2d1_hd U1692 ( .A(z_e[4]), .B(z_e[3]), .Y(n1254) );
  nr2d1_hd U1693 ( .A(z_e[6]), .B(z_e[5]), .Y(n1253) );
  nr4d1_hd U1694 ( .A(z_m[23]), .B(z_e[2]), .C(n1364), .D(n1365), .Y(n1255) );
  oa211d1_hd U1695 ( .A(z_e[0]), .B(n1275), .C(n1285), .D(n1259), .Y(n237) );
  nr2d1_hd U1696 ( .A(z_e[1]), .B(z_e[0]), .Y(n1263) );
  ao21d1_hd U1697 ( .A(z_e[0]), .B(z_e[1]), .C(n1263), .Y(n1261) );
  oa211d1_hd U1698 ( .A(n1261), .B(n1275), .C(n1285), .D(n1260), .Y(n236) );
  ivd1_hd U1699 ( .A(z_e[2]), .Y(n1262) );
  oa21d1_hd U1700 ( .A(n1263), .B(n1262), .C(n1266), .Y(n1264) );
  ao22d1_hd U1701 ( .A(n1162), .B(z[25]), .C(n1282), .D(n1264), .Y(n1265) );
  nr2d1_hd U1702 ( .A(z_e[3]), .B(n1266), .Y(n1270) );
  ao21d1_hd U1703 ( .A(z_e[3]), .B(n1266), .C(n1270), .Y(n1268) );
  oa211d1_hd U1704 ( .A(n1268), .B(n1275), .C(n524), .D(n1267), .Y(n234) );
  ivd1_hd U1705 ( .A(z_e[4]), .Y(n1269) );
  oa21d1_hd U1706 ( .A(n1270), .B(n1269), .C(n1273), .Y(n1271) );
  ao22d1_hd U1707 ( .A(n1162), .B(z[27]), .C(n1282), .D(n1271), .Y(n1272) );
  nr2d1_hd U1708 ( .A(z_e[5]), .B(n1273), .Y(n1278) );
  ao21d1_hd U1709 ( .A(z_e[5]), .B(n1273), .C(n1278), .Y(n1276) );
  oa211d1_hd U1710 ( .A(n1276), .B(n1275), .C(n524), .D(n1274), .Y(n232) );
  ivd1_hd U1711 ( .A(z_e[6]), .Y(n1277) );
  oa21d1_hd U1712 ( .A(n1278), .B(n1277), .C(n1283), .Y(n1279) );
  ao22d1_hd U1713 ( .A(n1161), .B(z[29]), .C(n1282), .D(n1279), .Y(n1280) );
  oa211d1_hd U1714 ( .A(z_e[7]), .B(n1283), .C(n1282), .D(n1281), .Y(n1284) );
  scg15d1_hd U1715 ( .A(n1489), .B(z[30]), .C(n524), .D(n1284), .Y(n230) );
  ao22d1_hd U1716 ( .A(n1330), .B(N35), .C(n1293), .D(z_s), .Y(n1286) );
  nr2d1_hd U1717 ( .A(n1165), .B(o_Z_STB), .Y(n179) );
  nr3d1_hd U1718 ( .A(n573), .B(n1219), .C(n1164), .Y(n171) );
  oa211d1_hd U1719 ( .A(state[1]), .B(n1291), .C(n1290), .D(n1368), .Y(n1292)
         );
  nr2d1_hd U1720 ( .A(n1293), .B(n1292), .Y(n160) );
  ao22d1_hd U1721 ( .A(n572), .B(z_m[23]), .C(n1165), .D(n177), .Y(n172) );
  ao22d1_hd U1722 ( .A(b_m[23]), .B(n574), .C(a_m[23]), .D(n517), .Y(n173) );
  ivd1_hd U1723 ( .A(n1328), .Y(n1335) );
  ao21d1_hd U1724 ( .A(n1335), .B(n1329), .C(n1301), .Y(n1300) );
  oa211d1_hd U1725 ( .A(n1300), .B(n1338), .C(n1299), .D(n1298), .Y(n355) );
  ao22d1_hd U1726 ( .A(n1135), .B(a[22]), .C(a_m[22]), .D(n1141), .Y(n1302) );
  scg14d1_hd U1727 ( .A(a_m[21]), .B(n536), .C(n1302), .Y(n354) );
  nr2d1_hd U1728 ( .A(n1304), .B(n1303), .Y(n161) );
  nr3d1_hd U1729 ( .A(n1218), .B(n518), .C(n1127), .Y(n156) );
  ao22d1_hd U1730 ( .A(n1132), .B(a[1]), .C(a_m[1]), .D(n1141), .Y(n1305) );
  scg14d1_hd U1731 ( .A(n388), .B(n535), .C(n1305), .Y(n348) );
  ao22d1_hd U1732 ( .A(n1133), .B(a[2]), .C(a_m[2]), .D(n1141), .Y(n1306) );
  scg14d1_hd U1733 ( .A(a_m[1]), .B(n535), .C(n1306), .Y(n347) );
  ao22d1_hd U1734 ( .A(n1133), .B(a[3]), .C(a_m[3]), .D(n1141), .Y(n1307) );
  scg14d1_hd U1735 ( .A(a_m[2]), .B(n537), .C(n1307), .Y(n346) );
  ao22d1_hd U1736 ( .A(n1133), .B(a[4]), .C(a_m[4]), .D(n1142), .Y(n1308) );
  scg14d1_hd U1737 ( .A(a_m[3]), .B(n535), .C(n1308), .Y(n345) );
  ao22d1_hd U1738 ( .A(n1133), .B(a[5]), .C(a_m[5]), .D(n1141), .Y(n1309) );
  scg14d1_hd U1739 ( .A(a_m[4]), .B(n538), .C(n1309), .Y(n344) );
  ao22d1_hd U1740 ( .A(n1133), .B(a[6]), .C(a_m[6]), .D(n1141), .Y(n1310) );
  scg14d1_hd U1741 ( .A(a_m[5]), .B(n536), .C(n1310), .Y(n343) );
  ao22d1_hd U1742 ( .A(n1133), .B(a[7]), .C(a_m[7]), .D(n1142), .Y(n1311) );
  scg14d1_hd U1743 ( .A(a_m[6]), .B(n536), .C(n1311), .Y(n342) );
  ao22d1_hd U1744 ( .A(n1134), .B(a[8]), .C(a_m[8]), .D(n1142), .Y(n1312) );
  scg14d1_hd U1745 ( .A(a_m[7]), .B(n535), .C(n1312), .Y(n341) );
  ao22d1_hd U1746 ( .A(n1134), .B(a[9]), .C(a_m[9]), .D(n1142), .Y(n1313) );
  scg14d1_hd U1747 ( .A(a_m[8]), .B(n538), .C(n1313), .Y(n340) );
  ao22d1_hd U1748 ( .A(n1134), .B(a[10]), .C(a_m[10]), .D(n1142), .Y(n1314) );
  scg14d1_hd U1749 ( .A(a_m[9]), .B(n536), .C(n1314), .Y(n339) );
  ao22d1_hd U1750 ( .A(n1134), .B(a[11]), .C(a_m[11]), .D(n1142), .Y(n1315) );
  scg14d1_hd U1751 ( .A(a_m[10]), .B(n536), .C(n1315), .Y(n338) );
  ao22d1_hd U1752 ( .A(n1134), .B(a[12]), .C(a_m[12]), .D(n1143), .Y(n1316) );
  scg14d1_hd U1753 ( .A(a_m[11]), .B(n537), .C(n1316), .Y(n337) );
  ao22d1_hd U1754 ( .A(n1134), .B(a[13]), .C(a_m[13]), .D(n1143), .Y(n1317) );
  scg14d1_hd U1755 ( .A(a_m[12]), .B(n537), .C(n1317), .Y(n336) );
  ao22d1_hd U1756 ( .A(n1215), .B(a[14]), .C(a_m[14]), .D(n1143), .Y(n1318) );
  scg14d1_hd U1757 ( .A(a_m[13]), .B(n536), .C(n1318), .Y(n335) );
  ao22d1_hd U1758 ( .A(n1215), .B(a[15]), .C(a_m[15]), .D(n1143), .Y(n1319) );
  scg14d1_hd U1759 ( .A(a_m[14]), .B(n535), .C(n1319), .Y(n334) );
  ao22d1_hd U1760 ( .A(n1140), .B(a[16]), .C(a_m[16]), .D(n1143), .Y(n1320) );
  scg14d1_hd U1761 ( .A(a_m[15]), .B(n537), .C(n1320), .Y(n333) );
  ao22d1_hd U1762 ( .A(n1140), .B(a[17]), .C(a_m[17]), .D(n1143), .Y(n1321) );
  scg14d1_hd U1763 ( .A(a_m[16]), .B(n537), .C(n1321), .Y(n332) );
  ao22d1_hd U1764 ( .A(n1215), .B(a[18]), .C(a_m[18]), .D(n1144), .Y(n1322) );
  scg14d1_hd U1765 ( .A(a_m[17]), .B(n538), .C(n1322), .Y(n331) );
  ao22d1_hd U1766 ( .A(n1215), .B(a[19]), .C(a_m[19]), .D(n1144), .Y(n1323) );
  scg14d1_hd U1767 ( .A(a_m[18]), .B(n538), .C(n1323), .Y(n330) );
  ao22d1_hd U1768 ( .A(n1135), .B(a[20]), .C(a_m[20]), .D(n1144), .Y(n1324) );
  scg14d1_hd U1769 ( .A(a_m[19]), .B(n538), .C(n1324), .Y(n329) );
  ao22d1_hd U1770 ( .A(n1135), .B(a[21]), .C(a_m[20]), .D(n535), .Y(n1326) );
  scg14d1_hd U1771 ( .A(a_m[21]), .B(n1327), .C(n1326), .Y(n328) );
  ao21d1_hd U1772 ( .A(n1335), .B(n1334), .C(n1333), .Y(n1339) );
  oa211d1_hd U1773 ( .A(n1339), .B(n1338), .C(n1337), .D(n1336), .Y(n310) );
  ao22d1_hd U1774 ( .A(n1135), .B(b[21]), .C(n1145), .D(n953), .Y(n1340) );
  scg14d1_hd U1775 ( .A(n962), .B(n523), .C(n1340), .Y(n309) );
  ao22d1_hd U1776 ( .A(n1135), .B(b[1]), .C(n1145), .D(n1057), .Y(n1341) );
  scg14d1_hd U1777 ( .A(n483), .B(n520), .C(n1341), .Y(n307) );
  ao22d1_hd U1778 ( .A(n1135), .B(b[2]), .C(n1145), .D(n1052), .Y(n1342) );
  scg14d1_hd U1779 ( .A(n1057), .B(n523), .C(n1342), .Y(n306) );
  ao22d1_hd U1780 ( .A(n1136), .B(b[3]), .C(n1146), .D(n1047), .Y(n1343) );
  scg14d1_hd U1781 ( .A(n1052), .B(n522), .C(n1343), .Y(n305) );
  ao22d1_hd U1782 ( .A(n1136), .B(b[4]), .C(n1145), .D(n1042), .Y(n1344) );
  scg14d1_hd U1783 ( .A(n1047), .B(n520), .C(n1344), .Y(n304) );
  ao22d1_hd U1784 ( .A(n1136), .B(b[5]), .C(n1146), .D(n1037), .Y(n1345) );
  scg14d1_hd U1785 ( .A(n1042), .B(n520), .C(n1345), .Y(n303) );
  ao22d1_hd U1786 ( .A(n1136), .B(b[6]), .C(n1146), .D(n1032), .Y(n1346) );
  scg14d1_hd U1787 ( .A(n1037), .B(n521), .C(n1346), .Y(n302) );
  ao22d1_hd U1788 ( .A(n1136), .B(b[7]), .C(n1146), .D(n1027), .Y(n1347) );
  scg14d1_hd U1789 ( .A(n1032), .B(n521), .C(n1347), .Y(n301) );
  ao22d1_hd U1790 ( .A(n1136), .B(b[8]), .C(n1146), .D(b_m[8]), .Y(n1348) );
  ao22d1_hd U1791 ( .A(n1137), .B(b[9]), .C(n1146), .D(n1014), .Y(n1349) );
  scg14d1_hd U1792 ( .A(b_m[8]), .B(n523), .C(n1349), .Y(n299) );
  ao22d1_hd U1793 ( .A(n1137), .B(b[10]), .C(n1147), .D(n1009), .Y(n1350) );
  scg14d1_hd U1794 ( .A(n1014), .B(n521), .C(n1350), .Y(n298) );
  ao22d1_hd U1795 ( .A(n1137), .B(b[11]), .C(n1147), .D(n1004), .Y(n1351) );
  scg14d1_hd U1796 ( .A(n1009), .B(n521), .C(n1351), .Y(n297) );
  ao22d1_hd U1797 ( .A(n1137), .B(b[12]), .C(n1147), .D(n999), .Y(n1352) );
  scg14d1_hd U1798 ( .A(n1004), .B(n522), .C(n1352), .Y(n296) );
  ao22d1_hd U1799 ( .A(n1137), .B(b[13]), .C(n1147), .D(n994), .Y(n1353) );
  scg14d1_hd U1800 ( .A(n999), .B(n522), .C(n1353), .Y(n295) );
  ao22d1_hd U1801 ( .A(n1137), .B(b[14]), .C(n1147), .D(n993), .Y(n1354) );
  scg14d1_hd U1802 ( .A(n994), .B(n522), .C(n1354), .Y(n294) );
  ao22d1_hd U1803 ( .A(n1138), .B(b[15]), .C(n1147), .D(n987), .Y(n1355) );
  scg14d1_hd U1804 ( .A(n993), .B(n520), .C(n1355), .Y(n293) );
  ao22d1_hd U1805 ( .A(n1138), .B(b[16]), .C(n1148), .D(n982), .Y(n1356) );
  scg14d1_hd U1806 ( .A(n987), .B(n522), .C(n1356), .Y(n292) );
  ao22d1_hd U1807 ( .A(n1138), .B(b[17]), .C(n1148), .D(n977), .Y(n1357) );
  scg14d1_hd U1808 ( .A(n982), .B(n523), .C(n1357), .Y(n291) );
  ao22d1_hd U1809 ( .A(n1138), .B(b[18]), .C(n1148), .D(n972), .Y(n1358) );
  scg14d1_hd U1810 ( .A(n977), .B(n523), .C(n1358), .Y(n290) );
  ao22d1_hd U1811 ( .A(n1138), .B(b[19]), .C(n1148), .D(n967), .Y(n1359) );
  ao22d1_hd U1812 ( .A(n1138), .B(b[20]), .C(n967), .D(n520), .Y(n1360) );
  scg14d1_hd U1813 ( .A(n1361), .B(n962), .C(n1360), .Y(n288) );
  ao22d1_hd U1814 ( .A(n1132), .B(b[22]), .C(n1145), .D(n487), .Y(n1362) );
  nr3d1_hd U1815 ( .A(z_e[2]), .B(z_e[1]), .C(n1364), .Y(n1366) );
  oa21d1_hd U1816 ( .A(n1366), .B(n1365), .C(z_e[9]), .Y(n36) );
  nr2d1_hd U1817 ( .A(n36), .B(n1394), .Y(n1375) );
  nr2d1_hd U1818 ( .A(round_bit), .B(sticky), .Y(n1367) );
  ao211d1_hd U1819 ( .A(n1367), .B(n1380), .C(net908), .D(n1368), .Y(n1377) );
  scg12d1_hd U1820 ( .A(z_m[1]), .B(z_m[2]), .C(n1380), .Y(n1407) );
  nd3d1_hd U1821 ( .A(z_m[4]), .B(n392), .C(n1407), .Y(n1415) );
  nd3d1_hd U1822 ( .A(z_m[8]), .B(n390), .C(n1422), .Y(n1430) );
  nd3d1_hd U1823 ( .A(z_m[12]), .B(n396), .C(n1437), .Y(n1445) );
  nd3d1_hd U1824 ( .A(z_m[16]), .B(n402), .C(n1452), .Y(n1461) );
  nd3d1_hd U1825 ( .A(n404), .B(n1469), .C(z_m[20]), .Y(n1372) );
  ao21d1_hd U1826 ( .A(n476), .B(n1372), .C(n460), .Y(n1482) );
  oa21d1_hd U1827 ( .A(z_m[21]), .B(n530), .C(n1482), .Y(n1485) );
  ao21d1_hd U1828 ( .A(n477), .B(n1374), .C(n1485), .Y(n1371) );
  nr2d1_hd U1829 ( .A(n528), .B(n1372), .Y(n1478) );
  oa21d1_hd U1830 ( .A(z_m[23]), .B(n1488), .C(n472), .Y(n1369) );
  ao22d1_hd U1831 ( .A(z_m[22]), .B(n1369), .C(n1150), .D(product[49]), .Y(
        n1370) );
  oa21d1_hd U1832 ( .A(n1371), .B(n1373), .C(n1370), .Y(n286) );
  nr4d1_hd U1833 ( .A(n1374), .B(n1373), .C(n1481), .D(n1372), .Y(n1376) );
  ao211d1_hd U1834 ( .A(n1377), .B(n1376), .C(n1375), .D(n1127), .Y(n1379) );
  ao22d1_hd U1835 ( .A(n1151), .B(product[26]), .C(z_m[0]), .D(n461), .Y(n1382) );
  ao22d1_hd U1836 ( .A(n1156), .B(z_m[1]), .C(n471), .D(n1386), .Y(n1381) );
  nd3d1_hd U1837 ( .A(n1382), .B(n1381), .C(n1400), .Y(n285) );
  ivd1_hd U1838 ( .A(n1394), .Y(n29) );
  ao21d1_hd U1839 ( .A(n1150), .B(product[25]), .C(n1383), .Y(n104) );
  ao22d1_hd U1840 ( .A(n1151), .B(product[24]), .C(n1384), .D(round_bit), .Y(
        n1385) );
  nr4d1_hd U1841 ( .A(product[12]), .B(product[13]), .C(product[14]), .D(
        product[15]), .Y(n1390) );
  nr4d1_hd U1842 ( .A(product[16]), .B(product[6]), .C(product[18]), .D(
        product[5]), .Y(n1389) );
  nr4d1_hd U1843 ( .A(product[17]), .B(product[22]), .C(product[10]), .D(
        product[11]), .Y(n1388) );
  nr4d1_hd U1844 ( .A(product[2]), .B(product[3]), .C(product[21]), .D(
        product[19]), .Y(n1387) );
  nd4d1_hd U1845 ( .A(n1390), .B(n1389), .C(n1388), .D(n1387), .Y(n1391) );
  nr4d1_hd U1846 ( .A(product[4]), .B(product[8]), .C(n1392), .D(n1391), .Y(
        n1399) );
  nr2d1_hd U1847 ( .A(n1393), .B(n1394), .Y(n1396) );
  ao22d1_hd U1848 ( .A(round_bit), .B(n1396), .C(sticky), .D(n1395), .Y(n1397)
         );
  oa21d1_hd U1849 ( .A(n1399), .B(n1398), .C(n1397), .Y(n283) );
  nd2bd1_hd U1850 ( .AN(z_m[1]), .B(n475), .Y(n1402) );
  scg4d1_hd U1851 ( .A(n1401), .B(z_m[0]), .C(n1403), .D(z_m[1]), .E(z_m[2]), 
        .F(n1484), .G(n1149), .H(product[27]), .Y(n282) );
  nd2bd1_hd U1852 ( .AN(n1403), .B(n1402), .Y(n1406) );
  nd3bd1_hd U1853 ( .AN(z_m[2]), .B(z_m[0]), .C(n476), .Y(n1404) );
  ao22d1_hd U1854 ( .A(n1151), .B(product[29]), .C(z_m[4]), .D(n1155), .Y(
        n1409) );
  oa21d1_hd U1855 ( .A(n529), .B(n1407), .C(n407), .Y(n1410) );
  ao22d1_hd U1856 ( .A(n470), .B(z_m[2]), .C(n392), .D(n1410), .Y(n1408) );
  oa211d1_hd U1857 ( .A(n392), .B(n1412), .C(n1409), .D(n1408), .Y(n280) );
  ivd1_hd U1858 ( .A(n1410), .Y(n1411) );
  oa21d1_hd U1859 ( .A(n392), .B(n1468), .C(n1411), .Y(n1414) );
  oa21d1_hd U1860 ( .A(z_m[4]), .B(n1412), .C(n473), .Y(n1413) );
  ao21d1_hd U1861 ( .A(n477), .B(n1415), .C(n461), .Y(n1418) );
  ao22d1_hd U1862 ( .A(n394), .B(n1418), .C(n1419), .D(n393), .Y(n1417) );
  ao22d1_hd U1863 ( .A(n1483), .B(product[31]), .C(z_m[6]), .D(n1155), .Y(
        n1416) );
  oa21d1_hd U1864 ( .A(n394), .B(n1468), .C(n1418), .Y(n1421) );
  oa21d1_hd U1865 ( .A(z_m[6]), .B(n1419), .C(n474), .Y(n1420) );
  ao22d1_hd U1866 ( .A(n1153), .B(product[33]), .C(z_m[8]), .D(n1156), .Y(
        n1424) );
  oa21d1_hd U1867 ( .A(n528), .B(n1422), .C(n407), .Y(n1425) );
  ao22d1_hd U1868 ( .A(n471), .B(z_m[6]), .C(n390), .D(n1425), .Y(n1423) );
  oa211d1_hd U1869 ( .A(n390), .B(n1427), .C(n1424), .D(n1423), .Y(n276) );
  ivd1_hd U1870 ( .A(n1425), .Y(n1426) );
  oa21d1_hd U1871 ( .A(n390), .B(n530), .C(n1426), .Y(n1429) );
  oa21d1_hd U1872 ( .A(z_m[8]), .B(n1427), .C(n474), .Y(n1428) );
  ao21d1_hd U1873 ( .A(n475), .B(n1430), .C(n460), .Y(n1433) );
  ao22d1_hd U1874 ( .A(n400), .B(n1433), .C(n1434), .D(n399), .Y(n1432) );
  ao22d1_hd U1875 ( .A(n1483), .B(product[35]), .C(z_m[10]), .D(n1156), .Y(
        n1431) );
  oa21d1_hd U1876 ( .A(n400), .B(n530), .C(n1433), .Y(n1436) );
  oa21d1_hd U1877 ( .A(z_m[10]), .B(n1434), .C(n472), .Y(n1435) );
  ao22d1_hd U1878 ( .A(n1149), .B(product[37]), .C(z_m[12]), .D(n1156), .Y(
        n1439) );
  oa21d1_hd U1879 ( .A(n530), .B(n1437), .C(n407), .Y(n1440) );
  ao22d1_hd U1880 ( .A(n470), .B(z_m[10]), .C(n396), .D(n1440), .Y(n1438) );
  oa211d1_hd U1881 ( .A(n396), .B(n1442), .C(n1439), .D(n1438), .Y(n272) );
  ivd1_hd U1882 ( .A(n1440), .Y(n1441) );
  oa21d1_hd U1883 ( .A(n396), .B(n529), .C(n1441), .Y(n1444) );
  oa21d1_hd U1884 ( .A(z_m[12]), .B(n1442), .C(n472), .Y(n1443) );
  ao21d1_hd U1885 ( .A(n476), .B(n1445), .C(n461), .Y(n1448) );
  ao22d1_hd U1886 ( .A(n398), .B(n1448), .C(n1449), .D(n397), .Y(n1447) );
  ao22d1_hd U1887 ( .A(n1483), .B(product[39]), .C(z_m[14]), .D(n1155), .Y(
        n1446) );
  oa21d1_hd U1888 ( .A(n398), .B(n529), .C(n1448), .Y(n1451) );
  oa21d1_hd U1889 ( .A(z_m[14]), .B(n1449), .C(n473), .Y(n1450) );
  ao22d1_hd U1890 ( .A(n1483), .B(product[41]), .C(z_m[16]), .D(n1155), .Y(
        n1454) );
  oa21d1_hd U1891 ( .A(n530), .B(n1452), .C(n1460), .Y(n1455) );
  ao22d1_hd U1892 ( .A(n471), .B(z_m[14]), .C(n402), .D(n1455), .Y(n1453) );
  oa211d1_hd U1893 ( .A(n402), .B(n1457), .C(n1454), .D(n1453), .Y(n268) );
  ivd1_hd U1894 ( .A(n1455), .Y(n1456) );
  oa21d1_hd U1895 ( .A(n402), .B(n528), .C(n1456), .Y(n1459) );
  oa21d1_hd U1896 ( .A(z_m[16]), .B(n1457), .C(n473), .Y(n1458) );
  ao21d1_hd U1897 ( .A(n477), .B(n1461), .C(n460), .Y(n1464) );
  ao22d1_hd U1898 ( .A(n406), .B(n1464), .C(n1465), .D(n405), .Y(n1463) );
  ao22d1_hd U1899 ( .A(n1150), .B(product[43]), .C(z_m[18]), .D(n1155), .Y(
        n1462) );
  oa21d1_hd U1900 ( .A(n406), .B(n528), .C(n1464), .Y(n1467) );
  oa21d1_hd U1901 ( .A(z_m[18]), .B(n1465), .C(n474), .Y(n1466) );
  ao22d1_hd U1902 ( .A(n1150), .B(product[45]), .C(z_m[20]), .D(n1155), .Y(
        n1471) );
  oa21d1_hd U1903 ( .A(n529), .B(n1469), .C(n407), .Y(n1474) );
  ao22d1_hd U1904 ( .A(n470), .B(z_m[18]), .C(n404), .D(n1474), .Y(n1470) );
  oa211d1_hd U1905 ( .A(n404), .B(n1473), .C(n1471), .D(n1470), .Y(n264) );
  oa21d1_hd U1906 ( .A(z_m[20]), .B(n1473), .C(n473), .Y(n1477) );
  ivd1_hd U1907 ( .A(n1474), .Y(n1475) );
  oa21d1_hd U1908 ( .A(n404), .B(n1468), .C(n1475), .Y(n1476) );
  scg4d1_hd U1909 ( .A(n1477), .B(z_m[19]), .C(n1476), .D(z_m[20]), .E(z_m[21]), .F(n1154), .G(n1149), .H(product[46]), .Y(n263) );
  ao22d1_hd U1910 ( .A(z_m[22]), .B(n1156), .C(n1150), .D(product[47]), .Y(
        n1480) );
  ao22d1_hd U1911 ( .A(n471), .B(z_m[20]), .C(n1478), .D(n1481), .Y(n1479) );
  oa211d1_hd U1912 ( .A(n1482), .B(n1481), .C(n1480), .D(n1479), .Y(n262) );
  ao22d1_hd U1913 ( .A(z_m[23]), .B(n1156), .C(n1150), .D(product[48]), .Y(
        n1487) );
  ao22d1_hd U1914 ( .A(z_m[22]), .B(n1485), .C(n470), .D(z_m[21]), .Y(n1486)
         );
  oa211d1_hd U1915 ( .A(z_m[22]), .B(n1488), .C(n1487), .D(n1486), .Y(n261) );
  ivd1_hd U1916 ( .A(o_AB_ACK), .Y(n20) );
endmodule

