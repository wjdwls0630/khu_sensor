
module float_adder ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3, C91_DATA2_4,
         C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8, n1, n2, n27, n265,
         n266, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n509, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23,
         C2_Z_22, C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16,
         C2_Z_15, C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_43J2_124_6938_n58, DP_OP_43J2_124_6938_n57,
         DP_OP_43J2_124_6938_n56, DP_OP_43J2_124_6938_n55,
         DP_OP_43J2_124_6938_n54, DP_OP_43J2_124_6938_n53,
         DP_OP_43J2_124_6938_n52, DP_OP_43J2_124_6938_n51,
         DP_OP_43J2_124_6938_n50, DP_OP_43J2_124_6938_n49,
         DP_OP_43J2_124_6938_n48, DP_OP_43J2_124_6938_n47,
         DP_OP_43J2_124_6938_n46, DP_OP_43J2_124_6938_n45,
         DP_OP_43J2_124_6938_n44, DP_OP_43J2_124_6938_n43,
         DP_OP_43J2_124_6938_n42, DP_OP_43J2_124_6938_n41,
         DP_OP_43J2_124_6938_n40, DP_OP_43J2_124_6938_n39,
         DP_OP_43J2_124_6938_n38, DP_OP_43J2_124_6938_n37,
         DP_OP_43J2_124_6938_n36, DP_OP_43J2_124_6938_n35,
         DP_OP_43J2_124_6938_n34, DP_OP_43J2_124_6938_n33,
         DP_OP_43J2_124_6938_n32, DP_OP_43J2_124_6938_n27,
         DP_OP_43J2_124_6938_n26, DP_OP_43J2_124_6938_n25,
         DP_OP_43J2_124_6938_n24, DP_OP_43J2_124_6938_n23,
         DP_OP_43J2_124_6938_n22, DP_OP_43J2_124_6938_n21,
         DP_OP_43J2_124_6938_n20, DP_OP_43J2_124_6938_n19,
         DP_OP_43J2_124_6938_n18, DP_OP_43J2_124_6938_n17,
         DP_OP_43J2_124_6938_n16, DP_OP_43J2_124_6938_n15,
         DP_OP_43J2_124_6938_n14, DP_OP_43J2_124_6938_n13,
         DP_OP_43J2_124_6938_n12, DP_OP_43J2_124_6938_n11,
         DP_OP_43J2_124_6938_n10, DP_OP_43J2_124_6938_n9,
         DP_OP_43J2_124_6938_n8, DP_OP_43J2_124_6938_n7,
         DP_OP_43J2_124_6938_n6, DP_OP_43J2_124_6938_n5,
         DP_OP_43J2_124_6938_n4, DP_OP_43J2_124_6938_n3,
         DP_OP_43J2_124_6938_n2, DP_OP_43J2_124_6938_n1,
         DP_OP_154J2_137_6175_n9, DP_OP_154J2_137_6175_n8,
         DP_OP_154J2_137_6175_n7, DP_OP_154J2_137_6175_n6,
         DP_OP_154J2_137_6175_n5, DP_OP_154J2_137_6175_n4,
         DP_OP_154J2_137_6175_n3, DP_OP_154J2_137_6175_n2, n1907, n1274, n1303,
         n1885, n1886, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J2_137_6175_U10 ( .A(n1907), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J2_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J2_137_6175_U9 ( .A(n1907), .B(z_e[2]), .CI(
        DP_OP_154J2_137_6175_n9), .CO(DP_OP_154J2_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J2_137_6175_U8 ( .A(n1907), .B(z_e[3]), .CI(
        DP_OP_154J2_137_6175_n8), .CO(DP_OP_154J2_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J2_137_6175_U7 ( .A(n1907), .B(z_e[4]), .CI(
        DP_OP_154J2_137_6175_n7), .CO(DP_OP_154J2_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J2_137_6175_U6 ( .A(n1907), .B(z_e[5]), .CI(
        DP_OP_154J2_137_6175_n6), .CO(DP_OP_154J2_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J2_137_6175_U5 ( .A(n1907), .B(z_e[6]), .CI(
        DP_OP_154J2_137_6175_n5), .CO(DP_OP_154J2_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J2_137_6175_U4 ( .A(n1907), .B(z_e[7]), .CI(
        DP_OP_154J2_137_6175_n4), .CO(DP_OP_154J2_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J2_137_6175_U3 ( .A(n1907), .B(z_e[8]), .CI(
        DP_OP_154J2_137_6175_n3), .CO(DP_OP_154J2_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n509), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n509), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n509), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n509), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n509), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n509), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n509), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n509), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n509), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n509), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n509), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n509), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n509), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n509), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n509), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n509), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n509), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n509), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n509), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n509), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n509), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n509), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n509), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n509), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n509), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n509), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n509), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n509), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n509), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n509), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n509), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n875), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n875), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n875), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n875), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n1274), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n1274), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n875), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n875), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n875), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n875), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n875), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n875), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n875), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n875), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n875), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n875), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n875), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n875), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n875), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n875), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n875), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n875), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n875), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n875), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n875), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n875), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n875), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n875), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n875), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n875), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n875), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n875), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n875), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n875), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n875), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n875), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n875), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n875), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n875), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n875), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n875), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n875), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n875), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n875), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n875), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n875), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n875), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n875), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n875), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n875), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n875), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n875), .CK(i_CLK), .Q(b[22]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n1274), .CK(i_CLK), .Q(sum[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n1274), .CK(i_CLK), .Q(sum[2]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n1274), .CK(i_CLK), .Q(sum[26]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n1274), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n1274), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n1274), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n1274), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n1274), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n1274), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n1274), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n1274), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n1274), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n1274), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n1274), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n1274), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n1274), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n1274), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n1274), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n1274), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n1274), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n1274), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n1274), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n1274), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n1274), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n1274), .CK(i_CLK), .Q(sum[25]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n1274), .CK(i_CLK), .Q(sum[1]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n875), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n875), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n875), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n875), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n1274), .CK(i_CLK), .Q(sum[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n875), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n875), .CK(i_CLK), .Q(b[28]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n875), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n875), .CK(i_CLK), .Q(b[25]) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n875), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n875), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n875), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n875), .CK(i_CLK), .Q(b[26]) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n875), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n875), .CK(i_CLK), .Q(b[23]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n265), .CK(i_CLK), .Q(guard) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1885), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1885), .CK(i_CLK), .Q(a_s) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n1886), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n1886), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J2_124_6938_U28 ( .A(C2_Z_0), .B(n1303), .CI(
        DP_OP_43J2_124_6938_n58), .CO(DP_OP_43J2_124_6938_n27), .S(N310) );
  fd1d1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK), .QN(n871) );
  fad1_hd DP_OP_43J2_124_6938_U27 ( .A(DP_OP_43J2_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J2_124_6938_n27), .CO(DP_OP_43J2_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J2_124_6938_U26 ( .A(DP_OP_43J2_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J2_124_6938_n26), .CO(DP_OP_43J2_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J2_124_6938_U25 ( .A(DP_OP_43J2_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J2_124_6938_n25), .CO(DP_OP_43J2_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J2_124_6938_U24 ( .A(DP_OP_43J2_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J2_124_6938_n24), .CO(DP_OP_43J2_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J2_124_6938_U23 ( .A(DP_OP_43J2_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J2_124_6938_n23), .CO(DP_OP_43J2_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J2_124_6938_U2 ( .A(DP_OP_43J2_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J2_124_6938_n2), .CO(DP_OP_43J2_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J2_124_6938_U3 ( .A(DP_OP_43J2_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J2_124_6938_n3), .CO(DP_OP_43J2_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J2_124_6938_U4 ( .A(DP_OP_43J2_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J2_124_6938_n4), .CO(DP_OP_43J2_124_6938_n3), .S(N334) );
  fad1_hd DP_OP_43J2_124_6938_U13 ( .A(DP_OP_43J2_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J2_124_6938_n13), .CO(DP_OP_43J2_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J2_124_6938_U14 ( .A(DP_OP_43J2_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J2_124_6938_n14), .CO(DP_OP_43J2_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J2_124_6938_U15 ( .A(DP_OP_43J2_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J2_124_6938_n15), .CO(DP_OP_43J2_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J2_124_6938_U16 ( .A(DP_OP_43J2_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J2_124_6938_n16), .CO(DP_OP_43J2_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J2_124_6938_U17 ( .A(DP_OP_43J2_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J2_124_6938_n17), .CO(DP_OP_43J2_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J2_124_6938_U18 ( .A(DP_OP_43J2_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J2_124_6938_n18), .CO(DP_OP_43J2_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J2_124_6938_U19 ( .A(DP_OP_43J2_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J2_124_6938_n19), .CO(DP_OP_43J2_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J2_124_6938_U20 ( .A(DP_OP_43J2_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J2_124_6938_n20), .CO(DP_OP_43J2_124_6938_n19), .S(N318)
         );
  fad1_hd DP_OP_43J2_124_6938_U21 ( .A(DP_OP_43J2_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J2_124_6938_n21), .CO(DP_OP_43J2_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J2_124_6938_U22 ( .A(DP_OP_43J2_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J2_124_6938_n22), .CO(DP_OP_43J2_124_6938_n21), .S(N316)
         );
  fad1_hd DP_OP_43J2_124_6938_U12 ( .A(DP_OP_43J2_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J2_124_6938_n12), .CO(DP_OP_43J2_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J2_124_6938_U11 ( .A(DP_OP_43J2_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J2_124_6938_n11), .CO(DP_OP_43J2_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J2_124_6938_U10 ( .A(DP_OP_43J2_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J2_124_6938_n10), .CO(DP_OP_43J2_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J2_124_6938_U9 ( .A(DP_OP_43J2_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J2_124_6938_n9), .CO(DP_OP_43J2_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J2_124_6938_U8 ( .A(DP_OP_43J2_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J2_124_6938_n8), .CO(DP_OP_43J2_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J2_124_6938_U7 ( .A(DP_OP_43J2_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J2_124_6938_n7), .CO(DP_OP_43J2_124_6938_n6), .S(N331) );
  fad1_hd DP_OP_43J2_124_6938_U6 ( .A(DP_OP_43J2_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J2_124_6938_n6), .CO(DP_OP_43J2_124_6938_n5), .S(N332) );
  fad1_hd DP_OP_43J2_124_6938_U5 ( .A(DP_OP_43J2_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J2_124_6938_n5), .CO(DP_OP_43J2_124_6938_n4), .S(N333) );
  clknd2d1_hd U523 ( .A(b_m[11]), .B(n1368), .Y(n891) );
  clknd2d1_hd U524 ( .A(b_m[10]), .B(n889), .Y(n890) );
  clknd2d1_hd U525 ( .A(n908), .B(n907), .Y(n909) );
  clknd2d1_hd U526 ( .A(a_m[23]), .B(n1293), .Y(n916) );
  clknd2d1_hd U527 ( .A(b_m[23]), .B(n1344), .Y(n914) );
  clknd2d1_hd U528 ( .A(b_m[9]), .B(n1372), .Y(n888) );
  clknd2d1_hd U529 ( .A(b_m[14]), .B(n1362), .Y(n896) );
  clknd2d1_hd U530 ( .A(a_e[4]), .B(n1487), .Y(n980) );
  clknd2d1_hd U531 ( .A(z_e[7]), .B(z_e[8]), .Y(n999) );
  clknd2d1_hd U532 ( .A(a_m[21]), .B(n1297), .Y(n912) );
  clknd2d1_hd U533 ( .A(n1510), .B(n1487), .Y(n964) );
  clknd2d1_hd U534 ( .A(n1013), .B(n1004), .Y(n1456) );
  clknd2d1_hd U535 ( .A(n996), .B(n995), .Y(n1528) );
  clknd2d1_hd U536 ( .A(b_e[1]), .B(n1391), .Y(n989) );
  clknd2d1_hd U537 ( .A(n1260), .B(n1520), .Y(n1526) );
  clknd2d1_hd U538 ( .A(n1521), .B(n1261), .Y(n1535) );
  clknd2d1_hd U539 ( .A(n1537), .B(n1261), .Y(n1530) );
  clknd2d1_hd U540 ( .A(n1012), .B(n1005), .Y(n1029) );
  clknd2d1_hd U541 ( .A(n977), .B(n976), .Y(n1005) );
  clknd2d1_hd U542 ( .A(n1524), .B(n1520), .Y(n1523) );
  clknd2d1_hd U543 ( .A(n1552), .B(n1483), .Y(n1336) );
  clknd2d1_hd U544 ( .A(n1521), .B(n1002), .Y(n1522) );
  clknd2d1_hd U545 ( .A(n1482), .B(n1461), .Y(n1468) );
  clknd2d1_hd U546 ( .A(n1450), .B(n1445), .Y(n1446) );
  clknd2d1_hd U547 ( .A(n1501), .B(n1510), .Y(n1508) );
  clknd2d1_hd U548 ( .A(b_e[2]), .B(n1498), .Y(n1492) );
  clknd2d1_hd U549 ( .A(a_e[2]), .B(n1392), .Y(n1426) );
  clknd2d1_hd U550 ( .A(n1450), .B(n1427), .Y(n1425) );
  clknd2d1_hd U551 ( .A(a_e[4]), .B(n1416), .Y(n1410) );
  clknd2d1_hd U552 ( .A(n1450), .B(n1411), .Y(n1409) );
  clknd2d1_hd U553 ( .A(a_e[6]), .B(n1402), .Y(n1395) );
  clknd2d1_hd U554 ( .A(n1405), .B(n1394), .Y(n1451) );
  clknd2d1_hd U555 ( .A(b_e[5]), .B(n1477), .Y(n1476) );
  clknd2d1_hd U556 ( .A(n1484), .B(b[28]), .Y(n1478) );
  clknd2d1_hd U557 ( .A(n1458), .B(n1483), .Y(n1555) );
  clknd2d1_hd U558 ( .A(n1002), .B(n1537), .Y(n1541) );
  clknd2d1_hd U559 ( .A(state[2]), .B(n1563), .Y(n1545) );
  clknd2d1_hd U560 ( .A(N41), .B(n1562), .Y(n1564) );
  clknd2d1_hd U561 ( .A(n1253), .B(n1243), .Y(n1234) );
  clknd2d1_hd U562 ( .A(n1253), .B(n1213), .Y(n1220) );
  clknd2d1_hd U563 ( .A(n1239), .B(n1234), .Y(n1230) );
  clknd2d1_hd U564 ( .A(n1268), .B(sum[27]), .Y(n1266) );
  clknd2d1_hd U565 ( .A(n1253), .B(n1189), .Y(n1196) );
  clknd2d1_hd U566 ( .A(n1253), .B(n1165), .Y(n1172) );
  clknd2d1_hd U567 ( .A(n1253), .B(n1141), .Y(n1148) );
  clknd2d1_hd U568 ( .A(n1253), .B(n1262), .Y(n1123) );
  clknd2d1_hd U569 ( .A(n1524), .B(n1261), .Y(n1098) );
  clknd2d1_hd U570 ( .A(n1264), .B(n1110), .Y(n1255) );
  clknd2d1_hd U571 ( .A(n1111), .B(n1110), .Y(n1113) );
  clknd2d1_hd U572 ( .A(z_m[19]), .B(z_m[20]), .Y(n1114) );
  clknd2d1_hd U573 ( .A(n1434), .B(n1502), .Y(n1066) );
  clknd2d1_hd U574 ( .A(n1420), .B(n1487), .Y(n1053) );
  clknd2d1_hd U575 ( .A(n1273), .B(n1462), .Y(n1039) );
  clknd2d1_hd U576 ( .A(a_e[0]), .B(b_e[0]), .Y(n1080) );
  clknd2d1_hd U577 ( .A(n1073), .B(n1068), .Y(n1067) );
  clknd2d1_hd U578 ( .A(n1059), .B(n1055), .Y(n1054) );
  clknd2d1_hd U579 ( .A(a_e[7]), .B(b_e[7]), .Y(n1034) );
  clknd2d1_hd U580 ( .A(n1045), .B(n1041), .Y(n1040) );
  clknd2d1_hd U581 ( .A(n1031), .B(n1030), .Y(n1083) );
  clknd2d1_hd U582 ( .A(n1559), .B(n1886), .Y(n1075) );
  clknd2d1_hd U583 ( .A(n953), .B(n1303), .Y(n940) );
  ivd1_hd U584 ( .A(a_m[26]), .Y(n1389) );
  clknd2d1_hd U585 ( .A(a_s), .B(n1005), .Y(n1011) );
  ivd2_hd U586 ( .A(n940), .Y(n950) );
  ivd2_hd U587 ( .A(n951), .Y(n1303) );
  clknd2d1_hd U588 ( .A(n1261), .B(n1260), .Y(n1525) );
  ivd4_hd U589 ( .A(n953), .Y(n869) );
  oa21d1_hd U590 ( .A(n920), .B(n919), .C(n918), .Y(n921) );
  clknd2d1_hd U591 ( .A(n1002), .B(n1260), .Y(n1519) );
  clknd2d1_hd U592 ( .A(n1444), .B(n1446), .Y(n1440) );
  clknd2d1_hd U593 ( .A(n1443), .B(a[25]), .Y(n1435) );
  clknd2d1_hd U594 ( .A(n1430), .B(a[26]), .Y(n1429) );
  clknd2d1_hd U595 ( .A(b[23]), .B(b[24]), .Y(n1512) );
  clknd2d1_hd U596 ( .A(n1417), .B(a[28]), .Y(n1413) );
  clknd2d1_hd U597 ( .A(n1412), .B(n1409), .Y(n1406) );
  clknd2d1_hd U598 ( .A(n1886), .B(n1444), .Y(n1452) );
  clknd2d1_hd U599 ( .A(b_e[4]), .B(n1501), .Y(n1491) );
  clknd2d1_hd U600 ( .A(n1499), .B(b[26]), .Y(n1495) );
  clknd2d1_hd U601 ( .A(n1002), .B(n1524), .Y(n1518) );
  clknd2d1_hd U602 ( .A(b[30]), .B(n1465), .Y(n1470) );
  clknd2d1_hd U603 ( .A(n1447), .B(n1446), .Y(n488) );
  clknd2d1_hd U604 ( .A(n1497), .B(n1496), .Y(n495) );
  clknd2d1_hd U605 ( .A(n1478), .B(n1471), .Y(n1472) );
  clknd2d1_hd U606 ( .A(n1254), .B(n1234), .Y(n1236) );
  clknd2d1_hd U607 ( .A(n1289), .B(n1288), .Y(n428) );
  clknd2d1_hd U608 ( .A(DP_OP_154J2_137_6175_n2), .B(n1287), .Y(n1285) );
  clknd2d1_hd U609 ( .A(n1267), .B(n1098), .Y(n265) );
  clknd2d1_hd U610 ( .A(n1561), .B(n1531), .Y(n1101) );
  clknd2d1_hd U611 ( .A(n1241), .B(sum[1]), .Y(n1099) );
  clknd2d1_hd U612 ( .A(n1082), .B(n1037), .Y(n362) );
  clknd2d1_hd U613 ( .A(n1088), .B(n1087), .Y(n1089) );
  clknd2d1_hd U614 ( .A(n1022), .B(n1021), .Y(n1025) );
  clknd2d1_hd U615 ( .A(n1450), .B(n1416), .Y(n1424) );
  clknd2d1_hd U616 ( .A(n1501), .B(n1498), .Y(n1507) );
  clknd2d1_hd U617 ( .A(n1450), .B(n1402), .Y(n1408) );
  clknd2d1_hd U618 ( .A(n1413), .B(n1403), .Y(n1404) );
  oa22d2_hd U619 ( .A(n954), .B(n1028), .C(a_s), .D(b_s), .Y(n951) );
  xo2d1_hd U620 ( .A(n1303), .B(DP_OP_43J2_124_6938_n1), .Y(N337) );
  oa211d8_hd U621 ( .A(b_m[26]), .B(n1389), .C(n1303), .D(n921), .Y(n953) );
  scg6d1_hd U622 ( .A(a_m[22]), .B(n915), .C(n1295), .Y(n913) );
  ivd3_hd U623 ( .A(n1525), .Y(n1274) );
  ivd4_hd U624 ( .A(n1518), .Y(n1885) );
  ivd1_hd U625 ( .A(a_m[24]), .Y(n1342) );
  scg6d1_hd U626 ( .A(n897), .B(a_m[13]), .C(n1314), .Y(n895) );
  scg10d1_hd U627 ( .A(n1445), .B(n1444), .C(n1518), .D(a[23]), .Y(n1447) );
  ad4d1_hd U628 ( .A(z_m[23]), .B(z_m[22]), .C(guard), .D(n1262), .Y(n1263) );
  nd2d2_hd U629 ( .A(n1483), .B(n870), .Y(n1388) );
  ivd2_hd U630 ( .A(n1455), .Y(n1552) );
  ivd2_hd U631 ( .A(n1559), .Y(n1096) );
  ivd2_hd U632 ( .A(n1266), .Y(n1241) );
  ad2d4_hd U633 ( .A(n1521), .B(n1520), .Y(n509) );
  ad2d1_hd U634 ( .A(a[23]), .B(a[24]), .Y(n1443) );
  ivd1_hd U635 ( .A(b_m[0]), .Y(n1338) );
  ivd1_hd U636 ( .A(b_m[1]), .Y(n1337) );
  ivd1_hd U637 ( .A(b_m[2]), .Y(n1335) );
  nr2d2_hd U638 ( .A(n1084), .B(n1523), .Y(n1094) );
  nid6_hd U639 ( .A(n27), .Y(n875) );
  clknd2d2_hd U640 ( .A(n1249), .B(n1560), .Y(n1228) );
  nr2ad1_hd U641 ( .A(n1269), .B(n1283), .Y(n1286) );
  ivd2_hd U642 ( .A(n1093), .Y(n1097) );
  nr2ad1_hd U643 ( .A(n1530), .B(n1229), .Y(n1235) );
  nr2ad1_hd U644 ( .A(n1106), .B(n265), .Y(n1229) );
  ivd1_hd U645 ( .A(b_m[3]), .Y(n1334) );
  ivd1_hd U646 ( .A(b_m[4]), .Y(n1332) );
  ivd1_hd U647 ( .A(n1281), .Y(n1283) );
  ivd1_hd U648 ( .A(b_m[5]), .Y(n1330) );
  ivd1_hd U649 ( .A(b_m[6]), .Y(n1328) );
  ivd1_hd U650 ( .A(b_m[7]), .Y(n1326) );
  ivd1_hd U651 ( .A(n1535), .Y(n1907) );
  scg6d1_hd U652 ( .A(n1527), .B(n1528), .C(n1885), .Y(n870) );
  ivd1_hd U653 ( .A(b_m[8]), .Y(n1324) );
  ivd1_hd U654 ( .A(b_m[9]), .Y(n1322) );
  nid2_hd U655 ( .A(n1095), .Y(n872) );
  ivd1_hd U656 ( .A(n1555), .Y(n1501) );
  nid2_hd U657 ( .A(n1240), .Y(n873) );
  ivd1_hd U658 ( .A(n1235), .Y(n1242) );
  ivd1_hd U659 ( .A(n1228), .Y(n1253) );
  ivd1_hd U660 ( .A(n1526), .Y(n1560) );
  ivd1_hd U661 ( .A(n1098), .Y(n1268) );
  ivd1_hd U662 ( .A(n1545), .Y(n1261) );
  ivd1_hd U663 ( .A(n1541), .Y(n1483) );
  nr2d1_hd U664 ( .A(n1541), .B(n1419), .Y(n1450) );
  ivd1_hd U665 ( .A(n1444), .Y(n1419) );
  ivd2_hd U666 ( .A(n870), .Y(n874) );
  ivd1_hd U667 ( .A(b_m[23]), .Y(n1293) );
  ivd1_hd U668 ( .A(b_m[16]), .Y(n1308) );
  ivd1_hd U669 ( .A(a_m[9]), .Y(n1372) );
  ivd1_hd U670 ( .A(b_m[12]), .Y(n1316) );
  ivd1_hd U671 ( .A(b_m[11]), .Y(n1318) );
  ivd1_hd U672 ( .A(b_m[15]), .Y(n1310) );
  ivd1_hd U673 ( .A(b_m[19]), .Y(n1301) );
  ivd1_hd U674 ( .A(b_m[20]), .Y(n1299) );
  ivd1_hd U675 ( .A(b_m[21]), .Y(n1297) );
  nr3d1_hd U676 ( .A(n1085), .B(n1046), .C(n1522), .Y(n1095) );
  ivd1_hd U677 ( .A(n1003), .Y(n1046) );
  ivd1_hd U678 ( .A(n1005), .Y(n1085) );
  nr2bd1_hd U679 ( .AN(n1488), .B(n1491), .Y(n1477) );
  ivd1_hd U680 ( .A(n1458), .Y(n1516) );
  ivd2_hd U681 ( .A(n1336), .Y(n1550) );
  ao21d1_hd U682 ( .A(n1483), .B(n997), .C(n1885), .Y(n1455) );
  ivd2_hd U683 ( .A(n1226), .Y(n1254) );
  nr2d1_hd U684 ( .A(n1535), .B(n1229), .Y(n1226) );
  ivd1_hd U685 ( .A(n1229), .Y(n1249) );
  ivd1_hd U686 ( .A(z_m[0]), .Y(n1250) );
  ivd1_hd U687 ( .A(n1530), .Y(n1561) );
  nr2bd1_hd U688 ( .AN(z_e[1]), .B(n999), .Y(n1023) );
  ivd1_hd U689 ( .A(n1522), .Y(n1886) );
  ivd1_hd U690 ( .A(n1450), .Y(n1433) );
  oa21d1_hd U691 ( .A(n1390), .B(n1456), .C(n874), .Y(n1444) );
  oa22ad1_hd U692 ( .A(n988), .B(n987), .C(n1453), .D(b_e[9]), .Y(n997) );
  ivd1_hd U693 ( .A(a_e[7]), .Y(n1400) );
  ivd1_hd U694 ( .A(a_e[0]), .Y(n1445) );
  ivd1_hd U695 ( .A(a_e[9]), .Y(n1453) );
  ivd1_hd U696 ( .A(b_e[4]), .Y(n1487) );
  ivd1_hd U697 ( .A(a_e[5]), .Y(n1411) );
  ivd1_hd U698 ( .A(a_e[3]), .Y(n1427) );
  nr2d1_hd U699 ( .A(n1548), .B(n1543), .Y(n1537) );
  ivd1_hd U700 ( .A(state[0]), .Y(n1548) );
  nr2d1_hd U701 ( .A(state[2]), .B(state[3]), .Y(n1002) );
  ivd1_hd U702 ( .A(a_m[25]), .Y(n1340) );
  ivd1_hd U703 ( .A(b_m[22]), .Y(n1295) );
  ivd1_hd U704 ( .A(a_m[21]), .Y(n1348) );
  ivd1_hd U705 ( .A(a_s), .Y(n1028) );
  ivd1_hd U706 ( .A(round_bit), .Y(n1104) );
  nd3d1_hd U707 ( .A(n1008), .B(n1004), .C(n1046), .Y(n1093) );
  oa21d1_hd U708 ( .A(n1536), .B(n1535), .C(n1534), .Y(n1562) );
  scg12d1_hd U709 ( .A(o_AB_ACK), .B(i_AB_STB), .C(n1519), .Y(n27) );
  oa21d1_hd U710 ( .A(n1522), .B(n1014), .C(n1523), .Y(n1559) );
  ao22d1_hd U711 ( .A(n1886), .B(n1029), .C(n1031), .D(n1084), .Y(n1082) );
  scg20d1_hd U712 ( .A(z_e[7]), .B(z_e[8]), .C(z_e[9]), .Y(n1084) );
  ivd1_hd U713 ( .A(n1523), .Y(n1031) );
  ivd1_hd U714 ( .A(n1557), .Y(n1505) );
  nr2d1_hd U715 ( .A(n1522), .B(n1516), .Y(n1557) );
  scg6d1_hd U716 ( .A(n1457), .B(n1547), .C(n1552), .Y(n2) );
  ivd1_hd U717 ( .A(n1456), .Y(n1547) );
  ivd1_hd U718 ( .A(z_m[20]), .Y(n1128) );
  ivd1_hd U719 ( .A(z_m[23]), .Y(n1258) );
  ivd1_hd U720 ( .A(z_m[22]), .Y(n1252) );
  ao211d1_hd U721 ( .A(n1105), .B(n1250), .C(n1244), .D(n1526), .Y(n1106) );
  ivd1_hd U722 ( .A(guard), .Y(n1244) );
  scg14d1_hd U723 ( .A(z_e[8]), .B(n1283), .C(n1270), .Y(n419) );
  ivd1_hd U724 ( .A(z_e[0]), .Y(n1282) );
  ivd1_hd U725 ( .A(z_m[17]), .Y(n1146) );
  ivd1_hd U726 ( .A(z_m[18]), .Y(n1134) );
  ivd1_hd U727 ( .A(z_m[14]), .Y(n1158) );
  ivd1_hd U728 ( .A(z_m[13]), .Y(n1170) );
  ivd1_hd U729 ( .A(z_m[10]), .Y(n1182) );
  ivd1_hd U730 ( .A(z_m[9]), .Y(n1194) );
  ivd1_hd U731 ( .A(z_m[6]), .Y(n1206) );
  ivd1_hd U732 ( .A(z_m[5]), .Y(n1218) );
  ivd1_hd U733 ( .A(z_m[2]), .Y(n1225) );
  ivd1_hd U734 ( .A(z_m[1]), .Y(n1243) );
  ivd1_hd U735 ( .A(z_m[21]), .Y(n1111) );
  ivd1_hd U736 ( .A(state[3]), .Y(n1563) );
  ivd1_hd U737 ( .A(a[30]), .Y(n1394) );
  nr2d1_hd U738 ( .A(n1548), .B(state[1]), .Y(n1524) );
  nr2d1_hd U739 ( .A(n997), .B(n1541), .Y(n1527) );
  ivd1_hd U740 ( .A(a_e[2]), .Y(n1434) );
  ivd1_hd U741 ( .A(a_e[1]), .Y(n1391) );
  ivd1_hd U742 ( .A(a_e[6]), .Y(n1273) );
  ivd1_hd U743 ( .A(b_e[8]), .Y(n1464) );
  ivd1_hd U744 ( .A(a_e[8]), .Y(n1449) );
  nr2d1_hd U745 ( .A(n1457), .B(n1007), .Y(n1008) );
  nr2d1_hd U746 ( .A(n965), .B(n964), .Y(n977) );
  ivd1_hd U747 ( .A(b_e[1]), .Y(n1510) );
  ivd1_hd U748 ( .A(b_e[3]), .Y(n1459) );
  ivd1_hd U749 ( .A(b_e[6]), .Y(n1462) );
  ivd1_hd U750 ( .A(b_e[5]), .Y(n1481) );
  ivd1_hd U751 ( .A(b_e[7]), .Y(n1466) );
  ivd1_hd U752 ( .A(b_e[0]), .Y(n1509) );
  nr2d1_hd U753 ( .A(n1390), .B(n1006), .Y(n1003) );
  ivd1_hd U754 ( .A(a_e[4]), .Y(n1420) );
  ivd1_hd U755 ( .A(state[1]), .Y(n1543) );
  ivd1_hd U756 ( .A(a_m[0]), .Y(n1386) );
  ivd1_hd U757 ( .A(a_m[1]), .Y(n1385) );
  ivd1_hd U758 ( .A(a_m[2]), .Y(n1384) );
  ivd1_hd U759 ( .A(a_m[4]), .Y(n1382) );
  ivd1_hd U760 ( .A(a_m[7]), .Y(n1376) );
  ivd1_hd U761 ( .A(b_m[10]), .Y(n1320) );
  ivd1_hd U762 ( .A(a_m[10]), .Y(n1370) );
  ivd1_hd U763 ( .A(a_m[13]), .Y(n1364) );
  ivd1_hd U764 ( .A(a_m[15]), .Y(n1360) );
  ivd1_hd U765 ( .A(a_m[20]), .Y(n1350) );
  ivd1_hd U766 ( .A(a_m[22]), .Y(n1346) );
  ivd1_hd U767 ( .A(b_m[25]), .Y(n1553) );
  ivd1_hd U768 ( .A(a_m[23]), .Y(n1344) );
  ivd1_hd U769 ( .A(b_m[18]), .Y(n1304) );
  ivd1_hd U770 ( .A(b_m[17]), .Y(n1306) );
  ivd1_hd U771 ( .A(b_m[13]), .Y(n1314) );
  ivd1_hd U772 ( .A(a_m[14]), .Y(n1362) );
  ivd1_hd U773 ( .A(a_m[11]), .Y(n1368) );
  ivd1_hd U774 ( .A(a_m[6]), .Y(n1378) );
  ivd1_hd U775 ( .A(a_m[5]), .Y(n1380) );
  ivd1_hd U776 ( .A(a_m[3]), .Y(n1383) );
  ivd1_hd U777 ( .A(a_m[8]), .Y(n1374) );
  ivd1_hd U778 ( .A(a_m[12]), .Y(n1366) );
  ivd1_hd U779 ( .A(b_m[14]), .Y(n1312) );
  ivd1_hd U780 ( .A(a_m[16]), .Y(n1358) );
  ivd1_hd U781 ( .A(a_m[17]), .Y(n1356) );
  ivd1_hd U782 ( .A(a_m[18]), .Y(n1354) );
  ivd1_hd U783 ( .A(a_m[19]), .Y(n1352) );
  ivd1_hd U784 ( .A(b_s), .Y(n954) );
  nd2bd1_hd U785 ( .AN(b[30]), .B(n1473), .Y(n1556) );
  nr2d1_hd U786 ( .A(n1563), .B(state[2]), .Y(n1520) );
  nr2d1_hd U787 ( .A(state[0]), .B(state[1]), .Y(n1260) );
  nr2d1_hd U788 ( .A(b_e[9]), .B(n1453), .Y(n988) );
  nr2d1_hd U789 ( .A(n1543), .B(state[0]), .Y(n1521) );
  ivd1_hd U790 ( .A(b_m[24]), .Y(n1291) );
  nr2d1_hd U791 ( .A(sum[27]), .B(n1098), .Y(n1240) );
  nr2d1_hd U792 ( .A(n1522), .B(n1029), .Y(n1004) );
  ao211d1_hd U793 ( .A(b_m[19]), .B(n1352), .C(b_m[18]), .D(n1354), .Y(n910)
         );
  ao22d1_hd U794 ( .A(a_m[20]), .B(n1299), .C(a_m[19]), .D(n1301), .Y(n908) );
  oa22d1_hd U795 ( .A(b_m[17]), .B(n1356), .C(b_m[16]), .D(n1358), .Y(n906) );
  ao22d1_hd U796 ( .A(a_m[14]), .B(n1312), .C(a_m[15]), .D(n1310), .Y(n901) );
  ao22d1_hd U797 ( .A(a_m[11]), .B(n1318), .C(a_m[12]), .D(n1316), .Y(n894) );
  ao211d1_hd U798 ( .A(a_m[1]), .B(n1337), .C(a_m[0]), .D(n1338), .Y(n877) );
  oa22d1_hd U799 ( .A(a_m[2]), .B(n1335), .C(a_m[1]), .D(n1337), .Y(n876) );
  oa22d1_hd U800 ( .A(n877), .B(n876), .C(b_m[3]), .D(n1383), .Y(n878) );
  ao21d1_hd U801 ( .A(a_m[2]), .B(n1335), .C(n878), .Y(n880) );
  oa22d1_hd U802 ( .A(a_m[4]), .B(n1332), .C(a_m[3]), .D(n1334), .Y(n879) );
  oa22d1_hd U803 ( .A(n880), .B(n879), .C(b_m[5]), .D(n1380), .Y(n881) );
  ao21d1_hd U804 ( .A(a_m[4]), .B(n1332), .C(n881), .Y(n883) );
  oa22d1_hd U805 ( .A(a_m[6]), .B(n1328), .C(a_m[5]), .D(n1330), .Y(n882) );
  oa22d1_hd U806 ( .A(n883), .B(n882), .C(b_m[6]), .D(n1378), .Y(n884) );
  ao21d1_hd U807 ( .A(a_m[7]), .B(n1326), .C(n884), .Y(n886) );
  oa22d1_hd U808 ( .A(a_m[7]), .B(n1326), .C(a_m[8]), .D(n1324), .Y(n885) );
  oa22d1_hd U809 ( .A(b_m[8]), .B(n1374), .C(n886), .D(n885), .Y(n887) );
  ao22d1_hd U810 ( .A(a_m[9]), .B(n1322), .C(n888), .D(n887), .Y(n889) );
  nr2d1_hd U811 ( .A(b_m[10]), .B(n889), .Y(n892) );
  oa211d1_hd U812 ( .A(a_m[10]), .B(n892), .C(n891), .D(n890), .Y(n893) );
  ao22d1_hd U813 ( .A(b_m[12]), .B(n1366), .C(n894), .D(n893), .Y(n897) );
  oa211d1_hd U814 ( .A(n897), .B(a_m[13]), .C(n896), .D(n895), .Y(n900) );
  nr2d1_hd U815 ( .A(a_m[15]), .B(n1310), .Y(n899) );
  nr2d1_hd U816 ( .A(a_m[16]), .B(n1308), .Y(n898) );
  ao211d1_hd U817 ( .A(n901), .B(n900), .C(n899), .D(n898), .Y(n905) );
  nr2d1_hd U818 ( .A(a_m[19]), .B(n1301), .Y(n903) );
  oa22d1_hd U819 ( .A(a_m[17]), .B(n1306), .C(a_m[18]), .D(n1304), .Y(n902) );
  nr2d1_hd U820 ( .A(n903), .B(n902), .Y(n904) );
  oa21d1_hd U821 ( .A(n906), .B(n905), .C(n904), .Y(n907) );
  oa22d1_hd U822 ( .A(n910), .B(n909), .C(a_m[20]), .D(n1299), .Y(n911) );
  ao22d1_hd U823 ( .A(b_m[21]), .B(n1348), .C(n912), .D(n911), .Y(n915) );
  oa211d1_hd U824 ( .A(a_m[22]), .B(n915), .C(n914), .D(n913), .Y(n917) );
  ao22d1_hd U825 ( .A(b_m[24]), .B(n1342), .C(n917), .D(n916), .Y(n920) );
  oa22d1_hd U826 ( .A(b_m[25]), .B(n1340), .C(b_m[24]), .D(n1342), .Y(n919) );
  ao22d1_hd U827 ( .A(b_m[25]), .B(n1340), .C(b_m[26]), .D(n1389), .Y(n918) );
  ao22d1_hd U828 ( .A(n869), .B(n1338), .C(n1386), .D(n953), .Y(C2_Z_0) );
  ao22d1_hd U829 ( .A(n869), .B(n1337), .C(n1385), .D(n953), .Y(C2_Z_1) );
  ao22d1_hd U830 ( .A(n869), .B(n1320), .C(n1370), .D(n953), .Y(C2_Z_10) );
  ao22d1_hd U831 ( .A(n869), .B(n1318), .C(n1368), .D(n953), .Y(C2_Z_11) );
  ao22d1_hd U832 ( .A(n869), .B(n1316), .C(n1366), .D(n953), .Y(C2_Z_12) );
  ao22d1_hd U833 ( .A(n869), .B(n1314), .C(n1364), .D(n953), .Y(C2_Z_13) );
  ao22d1_hd U834 ( .A(n869), .B(n1312), .C(n1362), .D(n953), .Y(C2_Z_14) );
  ao22d1_hd U835 ( .A(n869), .B(n1310), .C(n1360), .D(n953), .Y(C2_Z_15) );
  ao22d1_hd U836 ( .A(n869), .B(n1308), .C(n1358), .D(n953), .Y(C2_Z_16) );
  ao22d1_hd U837 ( .A(n869), .B(n1306), .C(n1356), .D(n953), .Y(C2_Z_17) );
  ao22d1_hd U838 ( .A(n869), .B(n1304), .C(n1354), .D(n953), .Y(C2_Z_18) );
  ao22d1_hd U839 ( .A(n869), .B(n1301), .C(n1352), .D(n953), .Y(C2_Z_19) );
  ao22d1_hd U840 ( .A(n869), .B(n1335), .C(n1384), .D(n953), .Y(C2_Z_2) );
  ao22d1_hd U841 ( .A(n869), .B(n1299), .C(n1350), .D(n953), .Y(C2_Z_20) );
  ao22d1_hd U842 ( .A(n869), .B(n1297), .C(n1348), .D(n953), .Y(C2_Z_21) );
  ao22d1_hd U843 ( .A(n869), .B(n1295), .C(n1346), .D(n953), .Y(C2_Z_22) );
  ao22d1_hd U844 ( .A(n869), .B(n1293), .C(n1344), .D(n953), .Y(C2_Z_23) );
  ao22d1_hd U845 ( .A(n869), .B(n1291), .C(n1342), .D(n953), .Y(C2_Z_24) );
  ao22d1_hd U846 ( .A(n869), .B(n1553), .C(n1340), .D(n953), .Y(C2_Z_25) );
  ivd1_hd U847 ( .A(b_m[26]), .Y(n922) );
  oa21d1_hd U848 ( .A(n951), .B(n922), .C(n1389), .Y(C2_Z_26) );
  ao22d1_hd U849 ( .A(n869), .B(n1334), .C(n1383), .D(n953), .Y(C2_Z_3) );
  ao22d1_hd U850 ( .A(n869), .B(n1332), .C(n1382), .D(n953), .Y(C2_Z_4) );
  ao22d1_hd U851 ( .A(n869), .B(n1330), .C(n1380), .D(n953), .Y(C2_Z_5) );
  ao22d1_hd U852 ( .A(n869), .B(n1328), .C(n1378), .D(n953), .Y(C2_Z_6) );
  ao22d1_hd U853 ( .A(n869), .B(n1326), .C(n1376), .D(n953), .Y(C2_Z_7) );
  ao22d1_hd U854 ( .A(n869), .B(n1324), .C(n1374), .D(n953), .Y(C2_Z_8) );
  ao22d1_hd U855 ( .A(n869), .B(n1322), .C(n1372), .D(n953), .Y(C2_Z_9) );
  nr2d1_hd U856 ( .A(n1389), .B(n922), .Y(n923) );
  ao22d1_hd U857 ( .A(n1303), .B(n923), .C(n922), .D(n951), .Y(
        DP_OP_43J2_124_6938_n32) );
  ao22d1_hd U858 ( .A(b_m[25]), .B(n951), .C(n950), .D(n1553), .Y(n924) );
  oa21d1_hd U859 ( .A(a_m[25]), .B(n953), .C(n924), .Y(DP_OP_43J2_124_6938_n33) );
  ao22d1_hd U860 ( .A(n869), .B(n1342), .C(b_m[24]), .D(n951), .Y(n925) );
  oa21d1_hd U861 ( .A(b_m[24]), .B(n940), .C(n925), .Y(DP_OP_43J2_124_6938_n34) );
  ao22d1_hd U862 ( .A(n950), .B(n1293), .C(n869), .D(n1344), .Y(n926) );
  oa21d1_hd U863 ( .A(n1303), .B(n1293), .C(n926), .Y(DP_OP_43J2_124_6938_n35)
         );
  ao22d1_hd U864 ( .A(b_m[22]), .B(n951), .C(n950), .D(n1295), .Y(n927) );
  oa21d1_hd U865 ( .A(a_m[22]), .B(n953), .C(n927), .Y(DP_OP_43J2_124_6938_n36) );
  ao22d1_hd U866 ( .A(n950), .B(n1297), .C(n869), .D(n1348), .Y(n928) );
  oa21d1_hd U867 ( .A(n1303), .B(n1297), .C(n928), .Y(DP_OP_43J2_124_6938_n37)
         );
  ao22d1_hd U868 ( .A(b_m[20]), .B(n951), .C(n950), .D(n1299), .Y(n929) );
  oa21d1_hd U869 ( .A(a_m[20]), .B(n953), .C(n929), .Y(DP_OP_43J2_124_6938_n38) );
  ao22d1_hd U870 ( .A(n950), .B(n1301), .C(n869), .D(n1352), .Y(n930) );
  oa21d1_hd U871 ( .A(n1303), .B(n1301), .C(n930), .Y(DP_OP_43J2_124_6938_n39)
         );
  ao22d1_hd U872 ( .A(n950), .B(n1304), .C(n869), .D(n1354), .Y(n931) );
  oa21d1_hd U873 ( .A(n1303), .B(n1304), .C(n931), .Y(DP_OP_43J2_124_6938_n40)
         );
  ao22d1_hd U874 ( .A(n950), .B(n1306), .C(n869), .D(n1356), .Y(n932) );
  oa21d1_hd U875 ( .A(n1303), .B(n1306), .C(n932), .Y(DP_OP_43J2_124_6938_n41)
         );
  ao22d1_hd U876 ( .A(n950), .B(n1308), .C(n869), .D(n1358), .Y(n933) );
  oa21d1_hd U877 ( .A(n1303), .B(n1308), .C(n933), .Y(DP_OP_43J2_124_6938_n42)
         );
  ao22d1_hd U878 ( .A(b_m[15]), .B(n951), .C(n950), .D(n1310), .Y(n934) );
  oa21d1_hd U879 ( .A(a_m[15]), .B(n953), .C(n934), .Y(DP_OP_43J2_124_6938_n43) );
  ao22d1_hd U880 ( .A(n950), .B(n1312), .C(n869), .D(n1362), .Y(n935) );
  oa21d1_hd U881 ( .A(n1303), .B(n1312), .C(n935), .Y(DP_OP_43J2_124_6938_n44)
         );
  ao22d1_hd U882 ( .A(b_m[13]), .B(n951), .C(n950), .D(n1314), .Y(n936) );
  oa21d1_hd U883 ( .A(a_m[13]), .B(n953), .C(n936), .Y(DP_OP_43J2_124_6938_n45) );
  ao22d1_hd U884 ( .A(n950), .B(n1316), .C(n869), .D(n1366), .Y(n937) );
  oa21d1_hd U885 ( .A(n1303), .B(n1316), .C(n937), .Y(DP_OP_43J2_124_6938_n46)
         );
  ao22d1_hd U886 ( .A(n950), .B(n1318), .C(n869), .D(n1368), .Y(n938) );
  oa21d1_hd U887 ( .A(n1303), .B(n1318), .C(n938), .Y(DP_OP_43J2_124_6938_n47)
         );
  ao22d1_hd U888 ( .A(n869), .B(n1370), .C(b_m[10]), .D(n951), .Y(n939) );
  oa21d1_hd U889 ( .A(b_m[10]), .B(n940), .C(n939), .Y(DP_OP_43J2_124_6938_n48) );
  ao22d1_hd U890 ( .A(n950), .B(n1322), .C(n869), .D(n1372), .Y(n941) );
  oa21d1_hd U891 ( .A(n1303), .B(n1322), .C(n941), .Y(DP_OP_43J2_124_6938_n49)
         );
  ao22d1_hd U892 ( .A(n950), .B(n1324), .C(n869), .D(n1374), .Y(n942) );
  oa21d1_hd U893 ( .A(n1303), .B(n1324), .C(n942), .Y(DP_OP_43J2_124_6938_n50)
         );
  ao22d1_hd U894 ( .A(b_m[7]), .B(n951), .C(n950), .D(n1326), .Y(n943) );
  oa21d1_hd U895 ( .A(a_m[7]), .B(n953), .C(n943), .Y(DP_OP_43J2_124_6938_n51)
         );
  ao22d1_hd U896 ( .A(n950), .B(n1328), .C(n869), .D(n1378), .Y(n944) );
  oa21d1_hd U897 ( .A(n1303), .B(n1328), .C(n944), .Y(DP_OP_43J2_124_6938_n52)
         );
  ao22d1_hd U898 ( .A(n950), .B(n1330), .C(n869), .D(n1380), .Y(n945) );
  oa21d1_hd U899 ( .A(n1303), .B(n1330), .C(n945), .Y(DP_OP_43J2_124_6938_n53)
         );
  ao22d1_hd U900 ( .A(b_m[4]), .B(n951), .C(n950), .D(n1332), .Y(n946) );
  oa21d1_hd U901 ( .A(a_m[4]), .B(n953), .C(n946), .Y(DP_OP_43J2_124_6938_n54)
         );
  ao22d1_hd U902 ( .A(n950), .B(n1334), .C(n869), .D(n1383), .Y(n947) );
  oa21d1_hd U903 ( .A(n1303), .B(n1334), .C(n947), .Y(DP_OP_43J2_124_6938_n55)
         );
  ao22d1_hd U904 ( .A(b_m[2]), .B(n951), .C(n950), .D(n1335), .Y(n948) );
  oa21d1_hd U905 ( .A(a_m[2]), .B(n953), .C(n948), .Y(DP_OP_43J2_124_6938_n56)
         );
  ao22d1_hd U906 ( .A(b_m[1]), .B(n951), .C(n950), .D(n1337), .Y(n949) );
  oa21d1_hd U907 ( .A(a_m[1]), .B(n953), .C(n949), .Y(DP_OP_43J2_124_6938_n57)
         );
  ao22d1_hd U908 ( .A(b_m[0]), .B(n951), .C(n950), .D(n1338), .Y(n952) );
  oa21d1_hd U909 ( .A(a_m[0]), .B(n953), .C(n952), .Y(DP_OP_43J2_124_6938_n58)
         );
  ao22d1_hd U910 ( .A(n869), .B(n954), .C(n1028), .D(n953), .Y(N338) );
  nd4d1_hd U911 ( .A(a_e[7]), .B(n1427), .C(n1420), .D(n1411), .Y(n955) );
  nr4d1_hd U912 ( .A(a_e[6]), .B(a_e[1]), .C(a_e[2]), .D(n955), .Y(n975) );
  nd4d1_hd U913 ( .A(n975), .B(a_e[0]), .C(a_e[9]), .D(a_e[8]), .Y(n1390) );
  nr4d1_hd U914 ( .A(a_m[22]), .B(a_m[18]), .C(a_m[17]), .D(a_m[24]), .Y(n963)
         );
  nd4d1_hd U915 ( .A(n1350), .B(n1362), .C(n1364), .D(n1389), .Y(n956) );
  nr4d1_hd U916 ( .A(a_m[23]), .B(a_m[16]), .C(a_m[25]), .D(n956), .Y(n962) );
  nd4d1_hd U917 ( .A(n1372), .B(n1374), .C(n1378), .D(n1376), .Y(n960) );
  nd4d1_hd U918 ( .A(n1348), .B(n1370), .C(n1368), .D(n1366), .Y(n959) );
  nd4d1_hd U919 ( .A(n1360), .B(n1382), .C(n1380), .D(n1352), .Y(n958) );
  nd4d1_hd U920 ( .A(n1386), .B(n1385), .C(n1384), .D(n1383), .Y(n957) );
  nr4d1_hd U921 ( .A(n960), .B(n959), .C(n958), .D(n957), .Y(n961) );
  nd3d1_hd U922 ( .A(n963), .B(n962), .C(n961), .Y(n1006) );
  nr2d1_hd U923 ( .A(n1509), .B(n1466), .Y(n966) );
  ivd1_hd U924 ( .A(b_e[2]), .Y(n1502) );
  nd4d1_hd U925 ( .A(n1481), .B(n1462), .C(n1502), .D(n1459), .Y(n965) );
  nd4d1_hd U926 ( .A(n966), .B(b_e[8]), .C(b_e[9]), .D(n977), .Y(n1457) );
  nr4d1_hd U927 ( .A(b_m[25]), .B(b_m[23]), .C(b_m[15]), .D(b_m[26]), .Y(n974)
         );
  nr4d1_hd U928 ( .A(b_m[22]), .B(b_m[6]), .C(b_m[18]), .D(b_m[24]), .Y(n973)
         );
  nd4d1_hd U929 ( .A(n1297), .B(n1312), .C(n1301), .D(n1308), .Y(n971) );
  nr4d1_hd U930 ( .A(b_m[0]), .B(b_m[1]), .C(b_m[2]), .D(b_m[3]), .Y(n967) );
  nd4d1_hd U931 ( .A(n967), .B(n1299), .C(n1320), .D(n1330), .Y(n970) );
  nd4d1_hd U932 ( .A(n1324), .B(n1318), .C(n1316), .D(n1306), .Y(n969) );
  nd4d1_hd U933 ( .A(n1314), .B(n1322), .C(n1332), .D(n1326), .Y(n968) );
  nr4d1_hd U934 ( .A(n971), .B(n970), .C(n969), .D(n968), .Y(n972) );
  nd3d1_hd U935 ( .A(n974), .B(n973), .C(n972), .Y(n1007) );
  nr2d1_hd U936 ( .A(n1003), .B(n1008), .Y(n1013) );
  nd4d1_hd U937 ( .A(n975), .B(n1453), .C(n1445), .D(n1449), .Y(n1012) );
  nr4d1_hd U938 ( .A(b_e[0]), .B(b_e[8]), .C(b_e[9]), .D(n1466), .Y(n976) );
  ao22d1_hd U939 ( .A(b_e[8]), .B(n1449), .C(b_e[7]), .D(n1400), .Y(n996) );
  ao22d1_hd U940 ( .A(n1411), .B(b_e[5]), .C(n1273), .D(b_e[6]), .Y(n991) );
  ao211d1_hd U941 ( .A(b_e[1]), .B(n1391), .C(b_e[0]), .D(n1445), .Y(n979) );
  oa22d1_hd U942 ( .A(b_e[2]), .B(n1434), .C(b_e[1]), .D(n1391), .Y(n978) );
  ao22d1_hd U943 ( .A(b_e[3]), .B(n1427), .C(b_e[2]), .D(n1434), .Y(n992) );
  oa21d1_hd U944 ( .A(n979), .B(n978), .C(n992), .Y(n981) );
  oa211d1_hd U945 ( .A(b_e[3]), .B(n1427), .C(n981), .D(n980), .Y(n983) );
  nr2d1_hd U946 ( .A(n1487), .B(a_e[4]), .Y(n994) );
  ivd1_hd U947 ( .A(n994), .Y(n982) );
  ao22d1_hd U948 ( .A(a_e[5]), .B(n1481), .C(n983), .D(n982), .Y(n985) );
  ao22d1_hd U949 ( .A(a_e[6]), .B(n1462), .C(a_e[7]), .D(n1466), .Y(n984) );
  scg16d1_hd U950 ( .A(n991), .B(n985), .C(n984), .Y(n986) );
  ao22d1_hd U951 ( .A(a_e[8]), .B(n1464), .C(n996), .D(n986), .Y(n987) );
  ivd1_hd U952 ( .A(n988), .Y(n990) );
  nd4d1_hd U953 ( .A(n992), .B(n991), .C(n990), .D(n989), .Y(n993) );
  ao211d1_hd U954 ( .A(b_e[0]), .B(n1445), .C(n994), .D(n993), .Y(n995) );
  scg6d1_hd U955 ( .A(n1390), .B(n1547), .C(n870), .Y(n1) );
  ivd1_hd U956 ( .A(z_e[4]), .Y(n1055) );
  nd3bd1_hd U957 ( .AN(z_e[3]), .B(z_e[9]), .C(n1055), .Y(n998) );
  nr4d1_hd U958 ( .A(z_e[5]), .B(z_e[6]), .C(z_e[2]), .D(n998), .Y(n1024) );
  ao21d1_hd U959 ( .A(z_e[9]), .B(n999), .C(n1024), .Y(n1001) );
  ao21d1_hd U960 ( .A(z_e[0]), .B(n1023), .C(n1001), .Y(n1000) );
  nr2d1_hd U961 ( .A(z_m[23]), .B(n1000), .Y(n1536) );
  nr2d1_hd U962 ( .A(n1001), .B(n1023), .Y(n1531) );
  ao22d1_hd U963 ( .A(n1536), .B(n1907), .C(n1561), .D(n1531), .Y(n1267) );
  scg4d1_hd U964 ( .A(n1907), .B(round_bit), .C(n1241), .D(sum[3]), .E(n1561), 
        .F(z_m[0]), .G(n873), .H(sum[2]), .Y(n266) );
  ivd1_hd U965 ( .A(n1012), .Y(n1086) );
  ao22d1_hd U966 ( .A(n1085), .B(n1007), .C(n1086), .D(n1006), .Y(n1087) );
  ao21d1_hd U967 ( .A(n1008), .B(n1028), .C(n1046), .Y(n1009) );
  oa21d1_hd U968 ( .A(n1085), .B(n1009), .C(b_s), .Y(n1010) );
  oa211d1_hd U969 ( .A(n1012), .B(n1011), .C(n1087), .D(n1010), .Y(n1015) );
  nr2bd1_hd U970 ( .AN(n1013), .B(n1029), .Y(n1014) );
  ao22d1_hd U971 ( .A(n1886), .B(n1015), .C(n1096), .D(z[31]), .Y(n1027) );
  ivd1_hd U972 ( .A(z_m[4]), .Y(n1212) );
  ivd1_hd U973 ( .A(z_m[3]), .Y(n1219) );
  nd4d1_hd U974 ( .A(n1225), .B(n1212), .C(n1219), .D(n1218), .Y(n1016) );
  nr4d1_hd U975 ( .A(z_m[22]), .B(z_m[0]), .C(z_m[1]), .D(n1016), .Y(n1022) );
  ivd1_hd U976 ( .A(z_m[12]), .Y(n1164) );
  ivd1_hd U977 ( .A(z_m[11]), .Y(n1171) );
  nd4d1_hd U978 ( .A(n1182), .B(n1164), .C(n1171), .D(n1170), .Y(n1020) );
  ivd1_hd U979 ( .A(z_m[8]), .Y(n1188) );
  ivd1_hd U980 ( .A(z_m[7]), .Y(n1195) );
  nd4d1_hd U981 ( .A(n1206), .B(n1188), .C(n1195), .D(n1194), .Y(n1019) );
  ivd1_hd U982 ( .A(z_m[19]), .Y(n1118) );
  nd4d1_hd U983 ( .A(n1111), .B(n1118), .C(n1128), .D(n1146), .Y(n1018) );
  ivd1_hd U984 ( .A(z_m[16]), .Y(n1135) );
  ivd1_hd U985 ( .A(z_m[15]), .Y(n1147) );
  nd4d1_hd U986 ( .A(n1158), .B(n1135), .C(n1147), .D(n1134), .Y(n1017) );
  nr4d1_hd U987 ( .A(n1020), .B(n1019), .C(n1018), .D(n1017), .Y(n1021) );
  nd4d1_hd U988 ( .A(n1024), .B(n1023), .C(n1258), .D(n1282), .Y(n1030) );
  oa211d1_hd U989 ( .A(n1025), .B(n1030), .C(n1031), .D(z_s), .Y(n1026) );
  oa211d1_hd U990 ( .A(n1028), .B(n1093), .C(n1027), .D(n1026), .Y(n361) );
  nr2d1_hd U991 ( .A(z_e[1]), .B(z_e[0]), .Y(n1073) );
  ivd1_hd U992 ( .A(z_e[2]), .Y(n1068) );
  nr2d1_hd U993 ( .A(z_e[3]), .B(n1067), .Y(n1059) );
  nr2d1_hd U994 ( .A(z_e[5]), .B(n1054), .Y(n1045) );
  ivd1_hd U995 ( .A(z_e[6]), .Y(n1041) );
  nr2d1_hd U996 ( .A(z_e[7]), .B(n1040), .Y(n1032) );
  ao211d1_hd U997 ( .A(z_e[7]), .B(n1040), .C(n1083), .D(n1032), .Y(n1036) );
  nd3d1_hd U998 ( .A(n1391), .B(n1510), .C(n1080), .Y(n1074) );
  nr2d1_hd U999 ( .A(n1074), .B(n1066), .Y(n1065) );
  nd3d1_hd U1000 ( .A(n1065), .B(n1427), .C(n1459), .Y(n1060) );
  nr2d1_hd U1001 ( .A(n1060), .B(n1053), .Y(n1052) );
  nd3d1_hd U1002 ( .A(n1052), .B(n1411), .C(n1481), .Y(n1047) );
  nr2d1_hd U1003 ( .A(n1047), .B(n1039), .Y(n1038) );
  nr2d1_hd U1004 ( .A(n1038), .B(n1034), .Y(n1033) );
  ao211d1_hd U1005 ( .A(n1038), .B(n1034), .C(n1075), .D(n1033), .Y(n1035) );
  ao211d1_hd U1006 ( .A(n1096), .B(z[30]), .C(n1036), .D(n1035), .Y(n1037) );
  ao21d1_hd U1007 ( .A(n1047), .B(n1039), .C(n1038), .Y(n1044) );
  ivd1_hd U1008 ( .A(n1083), .Y(n1070) );
  oa21d1_hd U1009 ( .A(n1045), .B(n1041), .C(n1040), .Y(n1042) );
  ao22d1_hd U1010 ( .A(n1096), .B(z[29]), .C(n1070), .D(n1042), .Y(n1043) );
  oa211d1_hd U1011 ( .A(n1044), .B(n1075), .C(n1082), .D(n1043), .Y(n363) );
  ao21d1_hd U1012 ( .A(z_e[5]), .B(n1054), .C(n1045), .Y(n1051) );
  ivd1_hd U1013 ( .A(n1075), .Y(n1090) );
  ao22d1_hd U1014 ( .A(a_e[5]), .B(n1090), .C(b_e[5]), .D(n1095), .Y(n1048) );
  oa22d1_hd U1015 ( .A(n1052), .B(n1048), .C(n1075), .D(n1047), .Y(n1049) );
  ao21d1_hd U1016 ( .A(n1096), .B(z[28]), .C(n1049), .Y(n1050) );
  oa211d1_hd U1017 ( .A(n1051), .B(n1083), .C(n1082), .D(n1050), .Y(n364) );
  ao21d1_hd U1018 ( .A(n1060), .B(n1053), .C(n1052), .Y(n1058) );
  oa21d1_hd U1019 ( .A(n1059), .B(n1055), .C(n1054), .Y(n1056) );
  ao22d1_hd U1020 ( .A(n1096), .B(z[27]), .C(n1070), .D(n1056), .Y(n1057) );
  oa211d1_hd U1021 ( .A(n1058), .B(n1075), .C(n1082), .D(n1057), .Y(n365) );
  ao21d1_hd U1022 ( .A(z_e[3]), .B(n1067), .C(n1059), .Y(n1064) );
  ao22d1_hd U1023 ( .A(a_e[3]), .B(n1090), .C(b_e[3]), .D(n1095), .Y(n1061) );
  oa22d1_hd U1024 ( .A(n1065), .B(n1061), .C(n1075), .D(n1060), .Y(n1062) );
  ao21d1_hd U1025 ( .A(n1096), .B(z[26]), .C(n1062), .Y(n1063) );
  oa211d1_hd U1026 ( .A(n1064), .B(n1083), .C(n1082), .D(n1063), .Y(n366) );
  ao21d1_hd U1027 ( .A(n1074), .B(n1066), .C(n1065), .Y(n1072) );
  oa21d1_hd U1028 ( .A(n1073), .B(n1068), .C(n1067), .Y(n1069) );
  ao22d1_hd U1029 ( .A(n1096), .B(z[25]), .C(n1070), .D(n1069), .Y(n1071) );
  oa211d1_hd U1030 ( .A(n1072), .B(n1075), .C(n1082), .D(n1071), .Y(n367) );
  ao21d1_hd U1031 ( .A(z_e[0]), .B(z_e[1]), .C(n1073), .Y(n1079) );
  ao22d1_hd U1032 ( .A(a_e[1]), .B(n1090), .C(b_e[1]), .D(n1095), .Y(n1076) );
  oa22d1_hd U1033 ( .A(n1076), .B(n1080), .C(n1075), .D(n1074), .Y(n1077) );
  ao21d1_hd U1034 ( .A(n1096), .B(z[24]), .C(n1077), .Y(n1078) );
  oa211d1_hd U1035 ( .A(n1079), .B(n1083), .C(n1082), .D(n1078), .Y(n368) );
  ao22d1_hd U1036 ( .A(n1096), .B(z[23]), .C(n1090), .D(n1080), .Y(n1081) );
  oa211d1_hd U1037 ( .A(z_e[0]), .B(n1083), .C(n1082), .D(n1081), .Y(n369) );
  ao22d1_hd U1038 ( .A(b_m[25]), .B(n872), .C(z_m[22]), .D(n1094), .Y(n1092)
         );
  nd3d1_hd U1039 ( .A(n1086), .B(n1085), .C(n1303), .Y(n1088) );
  ao22d1_hd U1040 ( .A(n1096), .B(z[22]), .C(n1090), .D(n1089), .Y(n1091) );
  oa211d1_hd U1041 ( .A(n1340), .B(n1093), .C(n1092), .D(n1091), .Y(n370) );
  scg4d1_hd U1042 ( .A(a_m[24]), .B(n1097), .C(n1096), .D(z[21]), .E(n872), 
        .F(b_m[24]), .G(n1094), .H(z_m[21]), .Y(n371) );
  scg4d1_hd U1043 ( .A(a_m[23]), .B(n1097), .C(n1096), .D(z[20]), .E(n1095), 
        .F(b_m[23]), .G(n1094), .H(z_m[20]), .Y(n372) );
  scg4d1_hd U1044 ( .A(a_m[22]), .B(n1097), .C(n1096), .D(z[19]), .E(n872), 
        .F(b_m[22]), .G(n1094), .H(z_m[19]), .Y(n373) );
  scg4d1_hd U1045 ( .A(a_m[21]), .B(n1097), .C(n1096), .D(z[18]), .E(n872), 
        .F(b_m[21]), .G(n1094), .H(z_m[18]), .Y(n374) );
  scg4d1_hd U1046 ( .A(a_m[20]), .B(n1097), .C(n1096), .D(z[17]), .E(n872), 
        .F(b_m[20]), .G(n1094), .H(z_m[17]), .Y(n375) );
  scg4d1_hd U1047 ( .A(a_m[19]), .B(n1097), .C(n1096), .D(z[16]), .E(n872), 
        .F(b_m[19]), .G(n1094), .H(z_m[16]), .Y(n376) );
  scg4d1_hd U1048 ( .A(a_m[18]), .B(n1097), .C(n1096), .D(z[15]), .E(n872), 
        .F(b_m[18]), .G(n1094), .H(z_m[15]), .Y(n377) );
  scg4d1_hd U1049 ( .A(a_m[17]), .B(n1097), .C(n1096), .D(z[14]), .E(n872), 
        .F(b_m[17]), .G(n1094), .H(z_m[14]), .Y(n378) );
  scg4d1_hd U1050 ( .A(a_m[16]), .B(n1097), .C(n1096), .D(z[13]), .E(n872), 
        .F(b_m[16]), .G(n1094), .H(z_m[13]), .Y(n379) );
  scg4d1_hd U1051 ( .A(a_m[15]), .B(n1097), .C(n1096), .D(z[12]), .E(n872), 
        .F(b_m[15]), .G(n1094), .H(z_m[12]), .Y(n380) );
  scg4d1_hd U1052 ( .A(a_m[14]), .B(n1097), .C(n1096), .D(z[11]), .E(n872), 
        .F(b_m[14]), .G(n1094), .H(z_m[11]), .Y(n381) );
  scg4d1_hd U1053 ( .A(b_m[13]), .B(n1095), .C(n1096), .D(z[10]), .E(a_m[13]), 
        .F(n1097), .G(n1094), .H(z_m[10]), .Y(n382) );
  scg4d1_hd U1054 ( .A(a_m[12]), .B(n1097), .C(n1096), .D(z[9]), .E(n872), .F(
        b_m[12]), .G(n1094), .H(z_m[9]), .Y(n383) );
  scg4d1_hd U1055 ( .A(a_m[11]), .B(n1097), .C(n1096), .D(z[8]), .E(n872), .F(
        b_m[11]), .G(n1094), .H(z_m[8]), .Y(n384) );
  scg4d1_hd U1056 ( .A(b_m[10]), .B(n1095), .C(n1096), .D(z[7]), .E(a_m[10]), 
        .F(n1097), .G(n1094), .H(z_m[7]), .Y(n385) );
  scg4d1_hd U1057 ( .A(a_m[9]), .B(n1097), .C(n1096), .D(z[6]), .E(n872), .F(
        b_m[9]), .G(n1094), .H(z_m[6]), .Y(n386) );
  scg4d1_hd U1058 ( .A(a_m[8]), .B(n1097), .C(n1096), .D(z[5]), .E(n872), .F(
        b_m[8]), .G(n1094), .H(z_m[5]), .Y(n387) );
  scg4d1_hd U1059 ( .A(a_m[7]), .B(n1097), .C(n1096), .D(z[4]), .E(n872), .F(
        b_m[7]), .G(n1094), .H(z_m[4]), .Y(n388) );
  scg4d1_hd U1060 ( .A(a_m[6]), .B(n1097), .C(n1096), .D(z[3]), .E(n872), .F(
        b_m[6]), .G(n1094), .H(z_m[3]), .Y(n389) );
  scg4d1_hd U1061 ( .A(a_m[5]), .B(n1097), .C(n1096), .D(z[2]), .E(n872), .F(
        b_m[5]), .G(n1094), .H(z_m[2]), .Y(n390) );
  scg4d1_hd U1062 ( .A(a_m[4]), .B(n1097), .C(n1096), .D(z[1]), .E(n872), .F(
        b_m[4]), .G(n1094), .H(z_m[1]), .Y(n391) );
  scg4d1_hd U1063 ( .A(a_m[3]), .B(n1097), .C(n1096), .D(z[0]), .E(n872), .F(
        b_m[3]), .G(n1094), .H(z_m[0]), .Y(n392) );
  ao22d1_hd U1064 ( .A(n1268), .B(sum[0]), .C(sticky), .D(n1098), .Y(n1100) );
  oa211d1_hd U1065 ( .A(n1104), .B(n1101), .C(n1100), .D(n1099), .Y(n393) );
  ao22d1_hd U1066 ( .A(n1241), .B(sum[2]), .C(n873), .D(sum[1]), .Y(n1103) );
  nd3d1_hd U1067 ( .A(n1561), .B(guard), .C(n265), .Y(n1102) );
  oa211d1_hd U1068 ( .A(n1104), .B(n265), .C(n1103), .D(n1102), .Y(n394) );
  nr2d1_hd U1069 ( .A(sticky), .B(round_bit), .Y(n1105) );
  ao22d1_hd U1070 ( .A(n1241), .B(sum[26]), .C(n873), .D(sum[25]), .Y(n1109)
         );
  nr3d1_hd U1071 ( .A(n1250), .B(n1243), .C(n1225), .Y(n1213) );
  nd3d1_hd U1072 ( .A(n1213), .B(z_m[4]), .C(z_m[3]), .Y(n1201) );
  nr3d1_hd U1073 ( .A(n1201), .B(n1218), .C(n1206), .Y(n1189) );
  nd3d1_hd U1074 ( .A(n1189), .B(z_m[8]), .C(z_m[7]), .Y(n1177) );
  nr3d1_hd U1075 ( .A(n1177), .B(n1194), .C(n1182), .Y(n1165) );
  nd3d1_hd U1076 ( .A(n1165), .B(z_m[12]), .C(z_m[11]), .Y(n1153) );
  nr3d1_hd U1077 ( .A(n1153), .B(n1170), .C(n1158), .Y(n1141) );
  nd3d1_hd U1078 ( .A(n1141), .B(z_m[16]), .C(z_m[15]), .Y(n1129) );
  nr3d1_hd U1079 ( .A(n1129), .B(n1134), .C(n1146), .Y(n1262) );
  oa21d1_hd U1080 ( .A(n1262), .B(n1526), .C(n1249), .Y(n1125) );
  ao21d1_hd U1081 ( .A(n1560), .B(n1114), .C(n1125), .Y(n1112) );
  oa21d1_hd U1082 ( .A(z_m[21]), .B(n1228), .C(n1112), .Y(n1251) );
  nr2d1_hd U1083 ( .A(n1111), .B(n1114), .Y(n1264) );
  ivd1_hd U1084 ( .A(n1123), .Y(n1110) );
  oa22d1_hd U1085 ( .A(z_m[22]), .B(n1255), .C(n1254), .D(n1111), .Y(n1107) );
  ao21d1_hd U1086 ( .A(z_m[22]), .B(n1251), .C(n1107), .Y(n1108) );
  oa211d1_hd U1087 ( .A(n1258), .B(n1242), .C(n1109), .D(n1108), .Y(n395) );
  ao22d1_hd U1088 ( .A(n1241), .B(sum[25]), .C(n873), .D(sum[24]), .Y(n1117)
         );
  oa22d1_hd U1089 ( .A(n1114), .B(n1113), .C(n1112), .D(n1111), .Y(n1115) );
  ao21d1_hd U1090 ( .A(z_m[20]), .B(n1226), .C(n1115), .Y(n1116) );
  oa211d1_hd U1091 ( .A(n1252), .B(n1242), .C(n1117), .D(n1116), .Y(n396) );
  ao21d1_hd U1092 ( .A(n1253), .B(n1118), .C(n1125), .Y(n1122) );
  ao22d1_hd U1093 ( .A(n1241), .B(sum[24]), .C(n873), .D(sum[23]), .Y(n1121)
         );
  oa21d1_hd U1094 ( .A(z_m[20]), .B(n1123), .C(n1254), .Y(n1119) );
  ao22d1_hd U1095 ( .A(z_m[21]), .B(n1235), .C(z_m[19]), .D(n1119), .Y(n1120)
         );
  oa211d1_hd U1096 ( .A(n1122), .B(n1128), .C(n1121), .D(n1120), .Y(n397) );
  ao22d1_hd U1097 ( .A(n1241), .B(sum[23]), .C(n873), .D(sum[22]), .Y(n1127)
         );
  oa22d1_hd U1098 ( .A(z_m[19]), .B(n1123), .C(n1254), .D(n1134), .Y(n1124) );
  ao21d1_hd U1099 ( .A(z_m[19]), .B(n1125), .C(n1124), .Y(n1126) );
  oa211d1_hd U1100 ( .A(n1128), .B(n1242), .C(n1127), .D(n1126), .Y(n398) );
  nr2d1_hd U1101 ( .A(n1228), .B(n1129), .Y(n1137) );
  ao21d1_hd U1102 ( .A(n1137), .B(n1134), .C(n1226), .Y(n1133) );
  ao22d1_hd U1103 ( .A(n1241), .B(sum[22]), .C(n873), .D(sum[21]), .Y(n1132)
         );
  ao21d1_hd U1104 ( .A(n1560), .B(n1129), .C(n1229), .Y(n1140) );
  oa21d1_hd U1105 ( .A(z_m[17]), .B(n1228), .C(n1140), .Y(n1130) );
  ao22d1_hd U1106 ( .A(z_m[19]), .B(n1235), .C(z_m[18]), .D(n1130), .Y(n1131)
         );
  oa211d1_hd U1107 ( .A(n1133), .B(n1146), .C(n1132), .D(n1131), .Y(n399) );
  ao22d1_hd U1108 ( .A(n1241), .B(sum[21]), .C(n873), .D(sum[20]), .Y(n1139)
         );
  oa22d1_hd U1109 ( .A(n1135), .B(n1254), .C(n1134), .D(n1242), .Y(n1136) );
  ao21d1_hd U1110 ( .A(n1137), .B(n1146), .C(n1136), .Y(n1138) );
  oa211d1_hd U1111 ( .A(n1140), .B(n1146), .C(n1139), .D(n1138), .Y(n400) );
  ao22d1_hd U1112 ( .A(n1241), .B(sum[20]), .C(n873), .D(sum[19]), .Y(n1145)
         );
  scg20d1_hd U1113 ( .A(n1526), .B(n1141), .C(n1229), .Y(n1149) );
  oa21d1_hd U1114 ( .A(z_m[15]), .B(n1228), .C(n1149), .Y(n1143) );
  oa21d1_hd U1115 ( .A(z_m[16]), .B(n1148), .C(n1254), .Y(n1142) );
  ao22d1_hd U1116 ( .A(z_m[16]), .B(n1143), .C(z_m[15]), .D(n1142), .Y(n1144)
         );
  oa211d1_hd U1117 ( .A(n1146), .B(n1242), .C(n1145), .D(n1144), .Y(n401) );
  ao22d1_hd U1118 ( .A(n1241), .B(sum[19]), .C(n873), .D(sum[18]), .Y(n1152)
         );
  ao22d1_hd U1119 ( .A(z_m[15]), .B(n1149), .C(n1148), .D(n1147), .Y(n1150) );
  ao21d1_hd U1120 ( .A(z_m[16]), .B(n1235), .C(n1150), .Y(n1151) );
  oa211d1_hd U1121 ( .A(n1158), .B(n1254), .C(n1152), .D(n1151), .Y(n402) );
  nr2d1_hd U1122 ( .A(n1228), .B(n1153), .Y(n1161) );
  ao21d1_hd U1123 ( .A(n1161), .B(n1158), .C(n1226), .Y(n1157) );
  ao22d1_hd U1124 ( .A(n1241), .B(sum[18]), .C(n873), .D(sum[17]), .Y(n1156)
         );
  ao21d1_hd U1125 ( .A(n1560), .B(n1153), .C(n1229), .Y(n1159) );
  oa21d1_hd U1126 ( .A(z_m[13]), .B(n1228), .C(n1159), .Y(n1154) );
  ao22d1_hd U1127 ( .A(z_m[14]), .B(n1154), .C(z_m[15]), .D(n1235), .Y(n1155)
         );
  oa211d1_hd U1128 ( .A(n1157), .B(n1170), .C(n1156), .D(n1155), .Y(n403) );
  ao22d1_hd U1129 ( .A(n1241), .B(sum[17]), .C(n873), .D(sum[16]), .Y(n1163)
         );
  oa22d1_hd U1130 ( .A(n1159), .B(n1170), .C(n1158), .D(n1242), .Y(n1160) );
  ao21d1_hd U1131 ( .A(n1161), .B(n1170), .C(n1160), .Y(n1162) );
  oa211d1_hd U1132 ( .A(n1164), .B(n1254), .C(n1163), .D(n1162), .Y(n404) );
  ao22d1_hd U1133 ( .A(n1241), .B(sum[16]), .C(n873), .D(sum[15]), .Y(n1169)
         );
  scg20d1_hd U1134 ( .A(n1526), .B(n1165), .C(n1229), .Y(n1173) );
  oa21d1_hd U1135 ( .A(z_m[11]), .B(n1228), .C(n1173), .Y(n1167) );
  oa21d1_hd U1136 ( .A(z_m[12]), .B(n1172), .C(n1254), .Y(n1166) );
  ao22d1_hd U1137 ( .A(z_m[12]), .B(n1167), .C(z_m[11]), .D(n1166), .Y(n1168)
         );
  oa211d1_hd U1138 ( .A(n1170), .B(n1242), .C(n1169), .D(n1168), .Y(n405) );
  ao22d1_hd U1139 ( .A(n1241), .B(sum[15]), .C(n873), .D(sum[14]), .Y(n1176)
         );
  ao22d1_hd U1140 ( .A(z_m[11]), .B(n1173), .C(n1172), .D(n1171), .Y(n1174) );
  ao21d1_hd U1141 ( .A(z_m[12]), .B(n1235), .C(n1174), .Y(n1175) );
  oa211d1_hd U1142 ( .A(n1182), .B(n1254), .C(n1176), .D(n1175), .Y(n406) );
  nr2d1_hd U1143 ( .A(n1228), .B(n1177), .Y(n1185) );
  ao21d1_hd U1144 ( .A(n1185), .B(n1182), .C(n1226), .Y(n1181) );
  ao22d1_hd U1145 ( .A(n1241), .B(sum[14]), .C(n873), .D(sum[13]), .Y(n1180)
         );
  ao21d1_hd U1146 ( .A(n1560), .B(n1177), .C(n1229), .Y(n1183) );
  oa21d1_hd U1147 ( .A(z_m[9]), .B(n1228), .C(n1183), .Y(n1178) );
  ao22d1_hd U1148 ( .A(z_m[10]), .B(n1178), .C(z_m[11]), .D(n1235), .Y(n1179)
         );
  oa211d1_hd U1149 ( .A(n1181), .B(n1194), .C(n1180), .D(n1179), .Y(n407) );
  ao22d1_hd U1150 ( .A(n1241), .B(sum[13]), .C(n873), .D(sum[12]), .Y(n1187)
         );
  oa22d1_hd U1151 ( .A(n1183), .B(n1194), .C(n1182), .D(n1242), .Y(n1184) );
  ao21d1_hd U1152 ( .A(n1185), .B(n1194), .C(n1184), .Y(n1186) );
  oa211d1_hd U1153 ( .A(n1188), .B(n1254), .C(n1187), .D(n1186), .Y(n408) );
  ao22d1_hd U1154 ( .A(n1241), .B(sum[12]), .C(n873), .D(sum[11]), .Y(n1193)
         );
  scg20d1_hd U1155 ( .A(n1526), .B(n1189), .C(n1229), .Y(n1197) );
  oa21d1_hd U1156 ( .A(z_m[7]), .B(n1228), .C(n1197), .Y(n1191) );
  oa21d1_hd U1157 ( .A(z_m[8]), .B(n1196), .C(n1254), .Y(n1190) );
  ao22d1_hd U1158 ( .A(z_m[8]), .B(n1191), .C(z_m[7]), .D(n1190), .Y(n1192) );
  oa211d1_hd U1159 ( .A(n1194), .B(n1242), .C(n1193), .D(n1192), .Y(n409) );
  ao22d1_hd U1160 ( .A(n1241), .B(sum[11]), .C(n873), .D(sum[10]), .Y(n1200)
         );
  ao22d1_hd U1161 ( .A(z_m[7]), .B(n1197), .C(n1196), .D(n1195), .Y(n1198) );
  ao21d1_hd U1162 ( .A(z_m[8]), .B(n1235), .C(n1198), .Y(n1199) );
  oa211d1_hd U1163 ( .A(n1206), .B(n1254), .C(n1200), .D(n1199), .Y(n410) );
  nr2d1_hd U1164 ( .A(n1228), .B(n1201), .Y(n1209) );
  ao21d1_hd U1165 ( .A(n1209), .B(n1206), .C(n1226), .Y(n1205) );
  ao22d1_hd U1166 ( .A(n1241), .B(sum[10]), .C(n873), .D(sum[9]), .Y(n1204) );
  ao21d1_hd U1167 ( .A(n1560), .B(n1201), .C(n1229), .Y(n1207) );
  oa21d1_hd U1168 ( .A(z_m[5]), .B(n1228), .C(n1207), .Y(n1202) );
  ao22d1_hd U1169 ( .A(z_m[6]), .B(n1202), .C(z_m[7]), .D(n1235), .Y(n1203) );
  oa211d1_hd U1170 ( .A(n1205), .B(n1218), .C(n1204), .D(n1203), .Y(n411) );
  ao22d1_hd U1171 ( .A(n1241), .B(sum[9]), .C(n873), .D(sum[8]), .Y(n1211) );
  oa22d1_hd U1172 ( .A(n1207), .B(n1218), .C(n1206), .D(n1242), .Y(n1208) );
  ao21d1_hd U1173 ( .A(n1209), .B(n1218), .C(n1208), .Y(n1210) );
  oa211d1_hd U1174 ( .A(n1212), .B(n1254), .C(n1211), .D(n1210), .Y(n412) );
  ao22d1_hd U1175 ( .A(n1241), .B(sum[8]), .C(n873), .D(sum[7]), .Y(n1217) );
  scg20d1_hd U1176 ( .A(n1526), .B(n1213), .C(n1229), .Y(n1221) );
  oa21d1_hd U1177 ( .A(z_m[3]), .B(n1228), .C(n1221), .Y(n1215) );
  oa21d1_hd U1178 ( .A(z_m[4]), .B(n1220), .C(n1254), .Y(n1214) );
  ao22d1_hd U1179 ( .A(z_m[4]), .B(n1215), .C(z_m[3]), .D(n1214), .Y(n1216) );
  oa211d1_hd U1180 ( .A(n1218), .B(n1242), .C(n1217), .D(n1216), .Y(n413) );
  ao22d1_hd U1181 ( .A(n1241), .B(sum[7]), .C(n873), .D(sum[6]), .Y(n1224) );
  ao22d1_hd U1182 ( .A(z_m[3]), .B(n1221), .C(n1220), .D(n1219), .Y(n1222) );
  ao21d1_hd U1183 ( .A(z_m[4]), .B(n1235), .C(n1222), .Y(n1223) );
  oa211d1_hd U1184 ( .A(n1225), .B(n1254), .C(n1224), .D(n1223), .Y(n414) );
  nr3d1_hd U1185 ( .A(z_m[2]), .B(n1228), .C(n1250), .Y(n1227) );
  nr2d1_hd U1186 ( .A(n1227), .B(n1226), .Y(n1233) );
  ao22d1_hd U1187 ( .A(n1241), .B(sum[6]), .C(n873), .D(sum[5]), .Y(n1232) );
  nr2d1_hd U1188 ( .A(z_m[0]), .B(n1228), .Y(n1246) );
  nr2d1_hd U1189 ( .A(n1229), .B(n1246), .Y(n1239) );
  ao22d1_hd U1190 ( .A(z_m[2]), .B(n1230), .C(z_m[3]), .D(n1235), .Y(n1231) );
  oa211d1_hd U1191 ( .A(n1233), .B(n1243), .C(n1232), .D(n1231), .Y(n415) );
  ao22d1_hd U1192 ( .A(n1241), .B(sum[5]), .C(n873), .D(sum[4]), .Y(n1238) );
  ao22d1_hd U1193 ( .A(z_m[0]), .B(n1236), .C(z_m[2]), .D(n1235), .Y(n1237) );
  oa211d1_hd U1194 ( .A(n1239), .B(n1243), .C(n1238), .D(n1237), .Y(n416) );
  ao22d1_hd U1195 ( .A(n1241), .B(sum[4]), .C(n873), .D(sum[3]), .Y(n1248) );
  oa22d1_hd U1196 ( .A(n1244), .B(n1254), .C(n1243), .D(n1242), .Y(n1245) );
  nr2d1_hd U1197 ( .A(n1246), .B(n1245), .Y(n1247) );
  oa211d1_hd U1198 ( .A(n1250), .B(n1249), .C(n1248), .D(n1247), .Y(n417) );
  ao21d1_hd U1199 ( .A(n1253), .B(n1252), .C(n1251), .Y(n1259) );
  oa21d1_hd U1200 ( .A(z_m[23]), .B(n1255), .C(n1254), .Y(n1256) );
  ao22d1_hd U1201 ( .A(n1268), .B(sum[26]), .C(z_m[22]), .D(n1256), .Y(n1257)
         );
  oa211d1_hd U1202 ( .A(n1259), .B(n1258), .C(n1257), .D(n1266), .Y(n418) );
  nd3d1_hd U1203 ( .A(n1560), .B(n1264), .C(n1263), .Y(n1265) );
  nd4d1_hd U1204 ( .A(n1267), .B(n1525), .C(n1266), .D(n1265), .Y(n1281) );
  nr3d1_hd U1205 ( .A(n1268), .B(state[1]), .C(n1560), .Y(n1269) );
  ao22d1_hd U1206 ( .A(a_e[8]), .B(n1274), .C(n1286), .D(C91_DATA2_8), .Y(
        n1270) );
  ao22d1_hd U1207 ( .A(z_e[7]), .B(n1283), .C(n1286), .D(C91_DATA2_7), .Y(
        n1271) );
  oa21d1_hd U1208 ( .A(n1400), .B(n1525), .C(n1271), .Y(n420) );
  ao22d1_hd U1209 ( .A(z_e[6]), .B(n1283), .C(n1286), .D(C91_DATA2_6), .Y(
        n1272) );
  oa21d1_hd U1210 ( .A(n1273), .B(n1525), .C(n1272), .Y(n421) );
  ao22d1_hd U1211 ( .A(z_e[5]), .B(n1283), .C(n1286), .D(C91_DATA2_5), .Y(
        n1275) );
  oa21d1_hd U1212 ( .A(n1411), .B(n1525), .C(n1275), .Y(n422) );
  ao22d1_hd U1213 ( .A(z_e[4]), .B(n1283), .C(n1286), .D(C91_DATA2_4), .Y(
        n1276) );
  oa21d1_hd U1214 ( .A(n1420), .B(n1525), .C(n1276), .Y(n423) );
  ao22d1_hd U1215 ( .A(z_e[3]), .B(n1283), .C(n1286), .D(C91_DATA2_3), .Y(
        n1277) );
  oa21d1_hd U1216 ( .A(n1427), .B(n1525), .C(n1277), .Y(n424) );
  ao22d1_hd U1217 ( .A(z_e[2]), .B(n1283), .C(n1286), .D(C91_DATA2_2), .Y(
        n1278) );
  oa21d1_hd U1218 ( .A(n1434), .B(n1525), .C(n1278), .Y(n425) );
  ao22d1_hd U1219 ( .A(z_e[1]), .B(n1283), .C(n1286), .D(C91_DATA2_1), .Y(
        n1279) );
  oa21d1_hd U1220 ( .A(n1391), .B(n1525), .C(n1279), .Y(n426) );
  ao22d1_hd U1221 ( .A(a_e[0]), .B(n1274), .C(n1286), .D(n1282), .Y(n1280) );
  oa21d1_hd U1222 ( .A(n1282), .B(n1281), .C(n1280), .Y(n427) );
  ao22d1_hd U1223 ( .A(a_e[9]), .B(n1274), .C(z_e[9]), .D(n1283), .Y(n1289) );
  ivd1_hd U1224 ( .A(z_e[9]), .Y(n1284) );
  ao22d1_hd U1225 ( .A(z_e[9]), .B(n1907), .C(n1535), .D(n1284), .Y(n1287) );
  oa211d1_hd U1226 ( .A(DP_OP_154J2_137_6175_n2), .B(n1287), .C(n1286), .D(
        n1285), .Y(n1288) );
  ao22d1_hd U1227 ( .A(b_m[25]), .B(n1550), .C(n1885), .D(b[21]), .Y(n1290) );
  oa21d1_hd U1228 ( .A(n1291), .B(n1552), .C(n1290), .Y(n429) );
  ao22d1_hd U1229 ( .A(b_m[24]), .B(n1550), .C(n1885), .D(b[20]), .Y(n1292) );
  oa21d1_hd U1230 ( .A(n1293), .B(n1552), .C(n1292), .Y(n430) );
  ao22d1_hd U1231 ( .A(b_m[23]), .B(n1550), .C(n1885), .D(b[19]), .Y(n1294) );
  oa21d1_hd U1232 ( .A(n1295), .B(n1552), .C(n1294), .Y(n431) );
  ao22d1_hd U1233 ( .A(b_m[22]), .B(n1550), .C(n1885), .D(b[18]), .Y(n1296) );
  oa21d1_hd U1234 ( .A(n1297), .B(n1552), .C(n1296), .Y(n432) );
  ao22d1_hd U1235 ( .A(b_m[21]), .B(n1550), .C(n1885), .D(b[17]), .Y(n1298) );
  oa21d1_hd U1236 ( .A(n1299), .B(n1552), .C(n1298), .Y(n433) );
  ao22d1_hd U1237 ( .A(b_m[20]), .B(n1550), .C(n1885), .D(b[16]), .Y(n1300) );
  oa21d1_hd U1238 ( .A(n1301), .B(n1552), .C(n1300), .Y(n434) );
  ao22d1_hd U1239 ( .A(b_m[19]), .B(n1550), .C(n1885), .D(b[15]), .Y(n1302) );
  oa21d1_hd U1240 ( .A(n1304), .B(n1552), .C(n1302), .Y(n435) );
  ao22d1_hd U1241 ( .A(b_m[18]), .B(n1550), .C(n1885), .D(b[14]), .Y(n1305) );
  oa21d1_hd U1242 ( .A(n1306), .B(n1552), .C(n1305), .Y(n436) );
  ao22d1_hd U1243 ( .A(b_m[17]), .B(n1550), .C(n1885), .D(b[13]), .Y(n1307) );
  oa21d1_hd U1244 ( .A(n1308), .B(n1552), .C(n1307), .Y(n437) );
  ao22d1_hd U1245 ( .A(b_m[16]), .B(n1550), .C(n1885), .D(b[12]), .Y(n1309) );
  oa21d1_hd U1246 ( .A(n1310), .B(n1552), .C(n1309), .Y(n438) );
  ao22d1_hd U1247 ( .A(b_m[15]), .B(n1550), .C(n1885), .D(b[11]), .Y(n1311) );
  oa21d1_hd U1248 ( .A(n1312), .B(n1552), .C(n1311), .Y(n439) );
  ao22d1_hd U1249 ( .A(b_m[14]), .B(n1550), .C(n1885), .D(b[10]), .Y(n1313) );
  oa21d1_hd U1250 ( .A(n1314), .B(n1552), .C(n1313), .Y(n440) );
  ao22d1_hd U1251 ( .A(b_m[13]), .B(n1550), .C(n1885), .D(b[9]), .Y(n1315) );
  oa21d1_hd U1252 ( .A(n1316), .B(n1552), .C(n1315), .Y(n441) );
  ao22d1_hd U1253 ( .A(b_m[12]), .B(n1550), .C(n1885), .D(b[8]), .Y(n1317) );
  oa21d1_hd U1254 ( .A(n1318), .B(n1552), .C(n1317), .Y(n442) );
  ao22d1_hd U1255 ( .A(b_m[11]), .B(n1550), .C(n1885), .D(b[7]), .Y(n1319) );
  oa21d1_hd U1256 ( .A(n1320), .B(n1552), .C(n1319), .Y(n443) );
  ao22d1_hd U1257 ( .A(b_m[10]), .B(n1550), .C(n1885), .D(b[6]), .Y(n1321) );
  oa21d1_hd U1258 ( .A(n1322), .B(n1552), .C(n1321), .Y(n444) );
  ao22d1_hd U1259 ( .A(b_m[9]), .B(n1550), .C(n1885), .D(b[5]), .Y(n1323) );
  oa21d1_hd U1260 ( .A(n1324), .B(n1552), .C(n1323), .Y(n445) );
  ao22d1_hd U1261 ( .A(b_m[8]), .B(n1550), .C(n1885), .D(b[4]), .Y(n1325) );
  oa21d1_hd U1262 ( .A(n1326), .B(n1552), .C(n1325), .Y(n446) );
  ao22d1_hd U1263 ( .A(b_m[7]), .B(n1550), .C(n1885), .D(b[3]), .Y(n1327) );
  oa21d1_hd U1264 ( .A(n1328), .B(n1552), .C(n1327), .Y(n447) );
  ao22d1_hd U1265 ( .A(b_m[6]), .B(n1550), .C(n1885), .D(b[2]), .Y(n1329) );
  oa21d1_hd U1266 ( .A(n1330), .B(n1552), .C(n1329), .Y(n448) );
  ao22d1_hd U1267 ( .A(b_m[5]), .B(n1550), .C(n1885), .D(b[1]), .Y(n1331) );
  oa21d1_hd U1268 ( .A(n1332), .B(n1552), .C(n1331), .Y(n449) );
  ao22d1_hd U1269 ( .A(b_m[4]), .B(n1550), .C(n1885), .D(b[0]), .Y(n1333) );
  oa21d1_hd U1270 ( .A(n1334), .B(n1552), .C(n1333), .Y(n450) );
  oa22d1_hd U1271 ( .A(n1335), .B(n1552), .C(n1334), .D(n1336), .Y(n451) );
  oa22d1_hd U1272 ( .A(n1337), .B(n1552), .C(n1335), .D(n1336), .Y(n452) );
  oa22d1_hd U1273 ( .A(n1885), .B(n1338), .C(n1337), .D(n1336), .Y(n453) );
  ao22d1_hd U1274 ( .A(a_m[24]), .B(n874), .C(n1885), .D(a[21]), .Y(n1339) );
  oa21d1_hd U1275 ( .A(n1340), .B(n1388), .C(n1339), .Y(n454) );
  ao22d1_hd U1276 ( .A(a_m[23]), .B(n874), .C(n1885), .D(a[20]), .Y(n1341) );
  oa21d1_hd U1277 ( .A(n1342), .B(n1388), .C(n1341), .Y(n455) );
  ao22d1_hd U1278 ( .A(a_m[22]), .B(n874), .C(n1885), .D(a[19]), .Y(n1343) );
  oa21d1_hd U1279 ( .A(n1344), .B(n1388), .C(n1343), .Y(n456) );
  ao22d1_hd U1280 ( .A(a_m[21]), .B(n874), .C(n1885), .D(a[18]), .Y(n1345) );
  oa21d1_hd U1281 ( .A(n1346), .B(n1388), .C(n1345), .Y(n457) );
  ao22d1_hd U1282 ( .A(a_m[20]), .B(n874), .C(n1885), .D(a[17]), .Y(n1347) );
  oa21d1_hd U1283 ( .A(n1348), .B(n1388), .C(n1347), .Y(n458) );
  ao22d1_hd U1284 ( .A(a_m[19]), .B(n874), .C(n1885), .D(a[16]), .Y(n1349) );
  oa21d1_hd U1285 ( .A(n1350), .B(n1388), .C(n1349), .Y(n459) );
  ao22d1_hd U1286 ( .A(a_m[18]), .B(n874), .C(n1885), .D(a[15]), .Y(n1351) );
  oa21d1_hd U1287 ( .A(n1352), .B(n1388), .C(n1351), .Y(n460) );
  ao22d1_hd U1288 ( .A(a_m[17]), .B(n874), .C(n1885), .D(a[14]), .Y(n1353) );
  oa21d1_hd U1289 ( .A(n1354), .B(n1388), .C(n1353), .Y(n461) );
  ao22d1_hd U1290 ( .A(a_m[16]), .B(n874), .C(n1885), .D(a[13]), .Y(n1355) );
  oa21d1_hd U1291 ( .A(n1356), .B(n1388), .C(n1355), .Y(n462) );
  ao22d1_hd U1292 ( .A(a_m[15]), .B(n874), .C(n1885), .D(a[12]), .Y(n1357) );
  oa21d1_hd U1293 ( .A(n1358), .B(n1388), .C(n1357), .Y(n463) );
  ao22d1_hd U1294 ( .A(a_m[14]), .B(n874), .C(n1885), .D(a[11]), .Y(n1359) );
  oa21d1_hd U1295 ( .A(n1360), .B(n1388), .C(n1359), .Y(n464) );
  ao22d1_hd U1296 ( .A(a_m[13]), .B(n874), .C(n1885), .D(a[10]), .Y(n1361) );
  oa21d1_hd U1297 ( .A(n1362), .B(n1388), .C(n1361), .Y(n465) );
  ao22d1_hd U1298 ( .A(a_m[12]), .B(n874), .C(n1885), .D(a[9]), .Y(n1363) );
  oa21d1_hd U1299 ( .A(n1364), .B(n1388), .C(n1363), .Y(n466) );
  ao22d1_hd U1300 ( .A(a_m[11]), .B(n874), .C(n1885), .D(a[8]), .Y(n1365) );
  oa21d1_hd U1301 ( .A(n1366), .B(n1388), .C(n1365), .Y(n467) );
  ao22d1_hd U1302 ( .A(a_m[10]), .B(n874), .C(n1885), .D(a[7]), .Y(n1367) );
  oa21d1_hd U1303 ( .A(n1368), .B(n1388), .C(n1367), .Y(n468) );
  ao22d1_hd U1304 ( .A(a_m[9]), .B(n874), .C(n1885), .D(a[6]), .Y(n1369) );
  oa21d1_hd U1305 ( .A(n1370), .B(n1388), .C(n1369), .Y(n469) );
  ao22d1_hd U1306 ( .A(a_m[8]), .B(n874), .C(n1885), .D(a[5]), .Y(n1371) );
  oa21d1_hd U1307 ( .A(n1372), .B(n1388), .C(n1371), .Y(n470) );
  ao22d1_hd U1308 ( .A(a_m[7]), .B(n874), .C(n1885), .D(a[4]), .Y(n1373) );
  oa21d1_hd U1309 ( .A(n1374), .B(n1388), .C(n1373), .Y(n471) );
  ao22d1_hd U1310 ( .A(a_m[6]), .B(n874), .C(n1885), .D(a[3]), .Y(n1375) );
  oa21d1_hd U1311 ( .A(n1376), .B(n1388), .C(n1375), .Y(n472) );
  ao22d1_hd U1312 ( .A(a_m[5]), .B(n874), .C(n1885), .D(a[2]), .Y(n1377) );
  oa21d1_hd U1313 ( .A(n1378), .B(n1388), .C(n1377), .Y(n473) );
  ao22d1_hd U1314 ( .A(a_m[4]), .B(n874), .C(n1885), .D(a[1]), .Y(n1379) );
  oa21d1_hd U1315 ( .A(n1380), .B(n1388), .C(n1379), .Y(n474) );
  ao22d1_hd U1316 ( .A(a_m[3]), .B(n874), .C(n1885), .D(a[0]), .Y(n1381) );
  oa21d1_hd U1317 ( .A(n1382), .B(n1388), .C(n1381), .Y(n475) );
  oa22d1_hd U1318 ( .A(n1384), .B(n870), .C(n1383), .D(n1388), .Y(n476) );
  oa22d1_hd U1319 ( .A(n1385), .B(n870), .C(n1384), .D(n1388), .Y(n477) );
  oa22d1_hd U1320 ( .A(n1885), .B(n1386), .C(n1385), .D(n1388), .Y(n478) );
  ao22d1_hd U1321 ( .A(a_m[25]), .B(n874), .C(n1885), .D(a[22]), .Y(n1387) );
  oa21d1_hd U1322 ( .A(n1389), .B(n1388), .C(n1387), .Y(n479) );
  nr2d1_hd U1323 ( .A(n1391), .B(n1445), .Y(n1392) );
  nr2d1_hd U1324 ( .A(n1427), .B(n1426), .Y(n1416) );
  nr2d1_hd U1325 ( .A(n1411), .B(n1410), .Y(n1402) );
  ao21d1_hd U1326 ( .A(n1483), .B(n1395), .C(n1419), .Y(n1401) );
  oa21d1_hd U1327 ( .A(a_e[7]), .B(n1433), .C(n1401), .Y(n1448) );
  nr4d1_hd U1328 ( .A(a_e[8]), .B(n1400), .C(n1433), .D(n1395), .Y(n1393) );
  ivd1_hd U1329 ( .A(n1435), .Y(n1430) );
  ivd1_hd U1330 ( .A(a[27]), .Y(n1418) );
  nr2d1_hd U1331 ( .A(n1429), .B(n1418), .Y(n1417) );
  ivd1_hd U1332 ( .A(a[29]), .Y(n1403) );
  nr2d1_hd U1333 ( .A(n1413), .B(n1403), .Y(n1397) );
  nr2d1_hd U1334 ( .A(n1397), .B(n1518), .Y(n1405) );
  scg17d1_hd U1335 ( .A(a_e[8]), .B(n1448), .C(n1393), .D(n1451), .Y(n480) );
  nr2d1_hd U1336 ( .A(n1518), .B(n1394), .Y(n1398) );
  nr2d1_hd U1337 ( .A(n1433), .B(n1395), .Y(n1396) );
  ao22d1_hd U1338 ( .A(n1398), .B(n1397), .C(n1396), .D(n1400), .Y(n1399) );
  oa211d1_hd U1339 ( .A(n1401), .B(n1400), .C(n1399), .D(n1451), .Y(n481) );
  ao21d1_hd U1340 ( .A(n1483), .B(n1410), .C(n1419), .Y(n1412) );
  ao22d1_hd U1341 ( .A(a_e[6]), .B(n1406), .C(n1405), .D(n1404), .Y(n1407) );
  oa211d1_hd U1342 ( .A(a_e[6]), .B(n1408), .C(n1407), .D(n1452), .Y(n482) );
  oa22d1_hd U1343 ( .A(n1412), .B(n1411), .C(n1410), .D(n1409), .Y(n1415) );
  oa211d1_hd U1344 ( .A(n1417), .B(a[28]), .C(n1885), .D(n1413), .Y(n1414) );
  nd3bd1_hd U1345 ( .AN(n1415), .B(n1452), .C(n1414), .Y(n483) );
  ao211d1_hd U1346 ( .A(n1429), .B(n1418), .C(n1417), .D(n1518), .Y(n1422) );
  ao21d1_hd U1347 ( .A(n1483), .B(n1426), .C(n1419), .Y(n1428) );
  ao21d1_hd U1348 ( .A(n1428), .B(n1425), .C(n1420), .Y(n1421) );
  nr2d1_hd U1349 ( .A(n1422), .B(n1421), .Y(n1423) );
  oa211d1_hd U1350 ( .A(a_e[4]), .B(n1424), .C(n1423), .D(n1452), .Y(n484) );
  oa22d1_hd U1351 ( .A(n1428), .B(n1427), .C(n1426), .D(n1425), .Y(n1432) );
  oa211d1_hd U1352 ( .A(n1430), .B(a[26]), .C(n1885), .D(n1429), .Y(n1431) );
  nd3bd1_hd U1353 ( .AN(n1432), .B(n1452), .C(n1431), .Y(n485) );
  nr2d1_hd U1354 ( .A(a_e[1]), .B(n1433), .Y(n1439) );
  oa21d1_hd U1355 ( .A(n1439), .B(n1440), .C(a_e[2]), .Y(n1438) );
  nd4d1_hd U1356 ( .A(a_e[1]), .B(a_e[0]), .C(n1450), .D(n1434), .Y(n1437) );
  oa211d1_hd U1357 ( .A(n1443), .B(a[25]), .C(n1885), .D(n1435), .Y(n1436) );
  nd4d1_hd U1358 ( .A(n1452), .B(n1438), .C(n1437), .D(n1436), .Y(n486) );
  oa21d1_hd U1359 ( .A(a[23]), .B(a[24]), .C(n1885), .Y(n1442) );
  ao22d1_hd U1360 ( .A(a_e[1]), .B(n1440), .C(a_e[0]), .D(n1439), .Y(n1441) );
  oa211d1_hd U1361 ( .A(n1443), .B(n1442), .C(n1441), .D(n1452), .Y(n487) );
  ao21d1_hd U1362 ( .A(n1450), .B(n1449), .C(n1448), .Y(n1454) );
  oa211d1_hd U1363 ( .A(n1454), .B(n1453), .C(n1452), .D(n1451), .Y(n489) );
  oa21d1_hd U1364 ( .A(n1457), .B(n1456), .C(n1455), .Y(n1458) );
  nr2d1_hd U1365 ( .A(n1510), .B(n1509), .Y(n1498) );
  nr2d1_hd U1366 ( .A(n1459), .B(n1492), .Y(n1488) );
  ao21d1_hd U1367 ( .A(n1488), .B(b_e[4]), .C(n1541), .Y(n1460) );
  nr2d1_hd U1368 ( .A(n1516), .B(n1460), .Y(n1482) );
  oa21d1_hd U1369 ( .A(n1462), .B(n1481), .C(n1483), .Y(n1461) );
  ao21d1_hd U1370 ( .A(n1501), .B(n1466), .C(n1468), .Y(n1554) );
  ivd1_hd U1371 ( .A(b[25]), .Y(n1500) );
  nr2d1_hd U1372 ( .A(n1512), .B(n1500), .Y(n1499) );
  ivd1_hd U1373 ( .A(b[27]), .Y(n1485) );
  nr2d1_hd U1374 ( .A(n1495), .B(n1485), .Y(n1484) );
  ivd1_hd U1375 ( .A(b[29]), .Y(n1471) );
  nr2d1_hd U1376 ( .A(n1478), .B(n1471), .Y(n1465) );
  nr2d1_hd U1377 ( .A(n1465), .B(n1518), .Y(n1473) );
  nr2d1_hd U1378 ( .A(n1462), .B(n1476), .Y(n1467) );
  nd3d1_hd U1379 ( .A(b_e[7]), .B(n1467), .C(n1464), .Y(n1463) );
  oa211d1_hd U1380 ( .A(n1554), .B(n1464), .C(n1556), .D(n1463), .Y(n490) );
  ao22d1_hd U1381 ( .A(b_e[7]), .B(n1468), .C(n1467), .D(n1466), .Y(n1469) );
  oa211d1_hd U1382 ( .A(n1518), .B(n1470), .C(n1469), .D(n1556), .Y(n491) );
  oa21d1_hd U1383 ( .A(b_e[5]), .B(n1555), .C(n1482), .Y(n1474) );
  ao22d1_hd U1384 ( .A(b_e[6]), .B(n1474), .C(n1473), .D(n1472), .Y(n1475) );
  oa211d1_hd U1385 ( .A(b_e[6]), .B(n1476), .C(n1475), .D(n1505), .Y(n492) );
  ao21d1_hd U1386 ( .A(n1477), .B(n1481), .C(n1557), .Y(n1480) );
  oa211d1_hd U1387 ( .A(n1484), .B(b[28]), .C(n1885), .D(n1478), .Y(n1479) );
  oa211d1_hd U1388 ( .A(n1482), .B(n1481), .C(n1480), .D(n1479), .Y(n493) );
  scg6d1_hd U1389 ( .A(n1492), .B(n1483), .C(n1516), .Y(n1494) );
  ao211d1_hd U1390 ( .A(n1495), .B(n1485), .C(n1484), .D(n1518), .Y(n1486) );
  ao211d1_hd U1391 ( .A(b_e[4]), .B(n1494), .C(n1557), .D(n1486), .Y(n1490) );
  nd3d1_hd U1392 ( .A(n1501), .B(n1488), .C(n1487), .Y(n1489) );
  oa211d1_hd U1393 ( .A(b_e[3]), .B(n1491), .C(n1490), .D(n1489), .Y(n494) );
  nr3d1_hd U1394 ( .A(b_e[3]), .B(n1555), .C(n1492), .Y(n1493) );
  ao211d1_hd U1395 ( .A(b_e[3]), .B(n1494), .C(n1557), .D(n1493), .Y(n1497) );
  oa211d1_hd U1396 ( .A(n1499), .B(b[26]), .C(n1885), .D(n1495), .Y(n1496) );
  ao211d1_hd U1397 ( .A(n1512), .B(n1500), .C(n1499), .D(n1518), .Y(n1504) );
  nr2d1_hd U1398 ( .A(b_e[0]), .B(n1555), .Y(n1515) );
  nr2d1_hd U1399 ( .A(n1516), .B(n1515), .Y(n1511) );
  ao21d1_hd U1400 ( .A(n1511), .B(n1508), .C(n1502), .Y(n1503) );
  nr2d1_hd U1401 ( .A(n1504), .B(n1503), .Y(n1506) );
  oa211d1_hd U1402 ( .A(b_e[2]), .B(n1507), .C(n1506), .D(n1505), .Y(n496) );
  oa22d1_hd U1403 ( .A(n1511), .B(n1510), .C(n1509), .D(n1508), .Y(n1514) );
  oa211d1_hd U1404 ( .A(b[23]), .B(b[24]), .C(n1885), .D(n1512), .Y(n1513) );
  scg13d1_hd U1405 ( .A(n1514), .B(n1557), .C(n1513), .Y(n497) );
  ao21d1_hd U1406 ( .A(n1516), .B(b_e[0]), .C(n1515), .Y(n1517) );
  oa21d1_hd U1407 ( .A(b[23]), .B(n1518), .C(n1517), .Y(n498) );
  ao211d1_hd U1408 ( .A(n1519), .B(n871), .C(i_RST), .D(n875), .Y(n499) );
  scg15d1_hd U1409 ( .A(n1563), .B(n1524), .C(n1523), .D(n1522), .Y(n1542) );
  nd3d1_hd U1410 ( .A(n509), .B(o_Z_STB), .C(i_Z_ACK), .Y(n1566) );
  nd4d1_hd U1411 ( .A(N41), .B(n1566), .C(n1526), .D(n1525), .Y(n1533) );
  ivd1_hd U1412 ( .A(n1527), .Y(n1529) );
  oa22d1_hd U1413 ( .A(n1531), .B(n1530), .C(n1529), .D(n1528), .Y(n1532) );
  nr4d1_hd U1414 ( .A(n875), .B(n1542), .C(n1533), .D(n1532), .Y(n1534) );
  ivd1_hd U1415 ( .A(n1562), .Y(n1539) );
  nr2d1_hd U1416 ( .A(n1537), .B(n1545), .Y(n1538) );
  ao22d1_hd U1417 ( .A(state[2]), .B(n1539), .C(N41), .D(n1538), .Y(n1540) );
  oa21d1_hd U1418 ( .A(n1541), .B(n1564), .C(n1540), .Y(n500) );
  nr2d1_hd U1419 ( .A(n1907), .B(n1542), .Y(n1544) );
  oa22d1_hd U1420 ( .A(n1544), .B(n1564), .C(n1543), .D(n1562), .Y(n501) );
  ao21d1_hd U1421 ( .A(state[1]), .B(n1545), .C(state[0]), .Y(n1546) );
  nr2d1_hd U1422 ( .A(n1547), .B(n1546), .Y(n1549) );
  oa22d1_hd U1423 ( .A(n1549), .B(n1564), .C(n1548), .D(n1562), .Y(n502) );
  ao22d1_hd U1424 ( .A(b_m[26]), .B(n1550), .C(n1885), .D(b[22]), .Y(n1551) );
  oa21d1_hd U1425 ( .A(n1553), .B(n1552), .C(n1551), .Y(n503) );
  oa21d1_hd U1426 ( .A(b_e[8]), .B(n1555), .C(n1554), .Y(n1558) );
  scg17d1_hd U1427 ( .A(b_e[9]), .B(n1558), .C(n1557), .D(n1556), .Y(n504) );
  nr3d1_hd U1428 ( .A(n1561), .B(n1560), .C(n1559), .Y(n1565) );
  oa22d1_hd U1429 ( .A(n1565), .B(n1564), .C(n1563), .D(n1562), .Y(n505) );
  ivd1_hd U1430 ( .A(n1566), .Y(n1567) );
  scg21d1_hd U1431 ( .A(n509), .B(o_Z_STB), .C(i_RST), .D(n1567), .Y(n506) );
endmodule


module iir_hpf ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   r_add_AB_STB, w_add_AB_ACK, w_add_Z_STB, r_add_Z_ACK, r_mult_AB_STB,
         w_mult_AB_ACK, w_mult_Z_STB, r_mult_Z_ACK, n_1_net_, N17, r_pstate_0_,
         r_counter_0_, N548, N553, N556, N559, n33, n34, n35, n36, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n221, n223, n260, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n341, n342, n343, n346, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589;
  wire   [31:0] r_add_A;
  wire   [31:0] r_add_B;
  wire   [31:0] w_add_Z;
  wire   [31:0] r_mult_A;
  wire   [31:0] r_mult_B;
  wire   [31:0] w_mult_Z;
  wire   [63:0] r_x_data;
  wire   [31:0] r_y_data;

  float_adder add ( .i_A(r_add_A), .i_B(r_add_B), .i_AB_STB(r_add_AB_STB), 
        .o_AB_ACK(w_add_AB_ACK), .o_Z(w_add_Z), .o_Z_STB(w_add_Z_STB), 
        .i_Z_ACK(r_add_Z_ACK), .i_CLK(i_CLK), .i_RST(N17) );
  float_multiplier mult ( .i_A(r_mult_A), .i_B(r_mult_B), .i_AB_STB(
        r_mult_AB_STB), .o_AB_ACK(w_mult_AB_ACK), .o_Z(w_mult_Z), .o_Z_STB(
        w_mult_Z_STB), .i_Z_ACK(r_mult_Z_ACK), .i_CLK(i_CLK), .i_RST(n_1_net_)
         );
  ivd1_hd I_5 ( .A(i_RSTN), .Y(n_1_net_) );
  fd3qd1_hd r_pstate_reg_1_ ( .D(n212), .CK(i_CLK), .SN(i_RSTN), .Q(n213) );
  fd3qd1_hd r_counter_reg_1_ ( .D(n211), .CK(i_CLK), .SN(i_RSTN), .Q(n221) );
  fd3qd1_hd r_counter_reg_0_ ( .D(n210), .CK(i_CLK), .SN(i_RSTN), .Q(n223) );
  ao22d1_hd U333 ( .A(n457), .B(w_add_Z[31]), .C(n456), .D(w_mult_Z[31]), .Y(
        n293) );
  ao22d1_hd U335 ( .A(n457), .B(w_add_Z[30]), .C(n456), .D(w_mult_Z[30]), .Y(
        n296) );
  ao22d1_hd U337 ( .A(n294), .B(w_add_Z[29]), .C(n456), .D(w_mult_Z[29]), .Y(
        n297) );
  ao22d1_hd U339 ( .A(n294), .B(w_add_Z[28]), .C(n456), .D(w_mult_Z[28]), .Y(
        n298) );
  ao22d1_hd U341 ( .A(n294), .B(w_add_Z[27]), .C(n456), .D(w_mult_Z[27]), .Y(
        n299) );
  ao22d1_hd U343 ( .A(n294), .B(w_add_Z[26]), .C(n456), .D(w_mult_Z[26]), .Y(
        n300) );
  ao22d1_hd U345 ( .A(n294), .B(w_add_Z[25]), .C(n456), .D(w_mult_Z[25]), .Y(
        n301) );
  ao22d1_hd U347 ( .A(n294), .B(w_add_Z[24]), .C(n456), .D(w_mult_Z[24]), .Y(
        n302) );
  ao22d1_hd U349 ( .A(n294), .B(w_add_Z[23]), .C(n456), .D(w_mult_Z[23]), .Y(
        n303) );
  ao22d1_hd U351 ( .A(n294), .B(w_add_Z[22]), .C(n456), .D(w_mult_Z[22]), .Y(
        n304) );
  ao22d1_hd U353 ( .A(n294), .B(w_add_Z[21]), .C(n456), .D(w_mult_Z[21]), .Y(
        n305) );
  ao22d1_hd U355 ( .A(n294), .B(w_add_Z[20]), .C(n456), .D(w_mult_Z[20]), .Y(
        n306) );
  ao22d1_hd U357 ( .A(n294), .B(w_add_Z[19]), .C(n456), .D(w_mult_Z[19]), .Y(
        n307) );
  ao22d1_hd U359 ( .A(n294), .B(w_add_Z[18]), .C(n456), .D(w_mult_Z[18]), .Y(
        n308) );
  ao22d1_hd U361 ( .A(n294), .B(w_add_Z[17]), .C(n295), .D(w_mult_Z[17]), .Y(
        n309) );
  ao22d1_hd U363 ( .A(n294), .B(w_add_Z[16]), .C(n295), .D(w_mult_Z[16]), .Y(
        n310) );
  ao22d1_hd U365 ( .A(n294), .B(w_add_Z[15]), .C(n295), .D(w_mult_Z[15]), .Y(
        n311) );
  ao22d1_hd U367 ( .A(n294), .B(w_add_Z[14]), .C(n295), .D(w_mult_Z[14]), .Y(
        n312) );
  ao22d1_hd U369 ( .A(n294), .B(w_add_Z[13]), .C(n295), .D(w_mult_Z[13]), .Y(
        n313) );
  ao22d1_hd U371 ( .A(n294), .B(w_add_Z[12]), .C(n456), .D(w_mult_Z[12]), .Y(
        n314) );
  ao22d1_hd U373 ( .A(n457), .B(w_add_Z[11]), .C(n456), .D(w_mult_Z[11]), .Y(
        n315) );
  ao22d1_hd U375 ( .A(n457), .B(w_add_Z[10]), .C(n456), .D(w_mult_Z[10]), .Y(
        n316) );
  ao22d1_hd U377 ( .A(n457), .B(w_add_Z[9]), .C(n456), .D(w_mult_Z[9]), .Y(
        n317) );
  ao22d1_hd U379 ( .A(n457), .B(w_add_Z[8]), .C(n456), .D(w_mult_Z[8]), .Y(
        n318) );
  ao22d1_hd U381 ( .A(n457), .B(w_add_Z[7]), .C(n456), .D(w_mult_Z[7]), .Y(
        n319) );
  ao22d1_hd U383 ( .A(n457), .B(w_add_Z[6]), .C(n456), .D(w_mult_Z[6]), .Y(
        n320) );
  ao22d1_hd U385 ( .A(n457), .B(w_add_Z[5]), .C(n456), .D(w_mult_Z[5]), .Y(
        n321) );
  ao22d1_hd U387 ( .A(n457), .B(w_add_Z[4]), .C(n456), .D(w_mult_Z[4]), .Y(
        n322) );
  ao22d1_hd U389 ( .A(n457), .B(w_add_Z[3]), .C(n456), .D(w_mult_Z[3]), .Y(
        n323) );
  ao22d1_hd U391 ( .A(n457), .B(w_add_Z[2]), .C(n456), .D(w_mult_Z[2]), .Y(
        n324) );
  ao22d1_hd U393 ( .A(n457), .B(w_add_Z[1]), .C(n456), .D(w_mult_Z[1]), .Y(
        n325) );
  ao22d1_hd U395 ( .A(n457), .B(w_add_Z[0]), .C(n456), .D(w_mult_Z[0]), .Y(
        n326) );
  scg5d1_hd U402 ( .A(n458), .B(r_add_A[30]), .C(w_mult_Z[30]), .D(n455), .E(
        n34), .F(r_x_data[30]), .Y(n413) );
  scg5d1_hd U403 ( .A(n458), .B(r_add_A[29]), .C(w_mult_Z[29]), .D(n455), .E(
        n34), .F(r_x_data[29]), .Y(n414) );
  scg5d1_hd U404 ( .A(n458), .B(r_add_A[28]), .C(w_mult_Z[28]), .D(n455), .E(
        n34), .F(r_x_data[28]), .Y(n415) );
  scg5d1_hd U405 ( .A(n458), .B(r_add_A[27]), .C(w_mult_Z[27]), .D(n455), .E(
        n34), .F(r_x_data[27]), .Y(n416) );
  scg5d1_hd U406 ( .A(n458), .B(r_add_A[26]), .C(w_mult_Z[26]), .D(n455), .E(
        n34), .F(r_x_data[26]), .Y(n417) );
  scg5d1_hd U407 ( .A(n458), .B(r_add_A[25]), .C(w_mult_Z[25]), .D(n455), .E(
        n34), .F(r_x_data[25]), .Y(n418) );
  scg5d1_hd U408 ( .A(n458), .B(r_add_A[24]), .C(w_mult_Z[24]), .D(n455), .E(
        n34), .F(r_x_data[24]), .Y(n419) );
  scg5d1_hd U409 ( .A(n458), .B(r_add_A[23]), .C(w_mult_Z[23]), .D(n455), .E(
        n34), .F(r_x_data[23]), .Y(n420) );
  scg5d1_hd U410 ( .A(n458), .B(r_add_A[22]), .C(w_mult_Z[22]), .D(n455), .E(
        n34), .F(r_x_data[22]), .Y(n421) );
  scg5d1_hd U411 ( .A(n458), .B(r_add_A[21]), .C(w_mult_Z[21]), .D(n455), .E(
        n34), .F(r_x_data[21]), .Y(n422) );
  scg5d1_hd U412 ( .A(n458), .B(r_add_A[20]), .C(w_mult_Z[20]), .D(n455), .E(
        n34), .F(r_x_data[20]), .Y(n423) );
  scg5d1_hd U413 ( .A(n458), .B(r_add_A[19]), .C(w_mult_Z[19]), .D(n455), .E(
        n34), .F(r_x_data[19]), .Y(n424) );
  scg5d1_hd U414 ( .A(n458), .B(r_add_A[18]), .C(w_mult_Z[18]), .D(n455), .E(
        n34), .F(r_x_data[18]), .Y(n425) );
  scg5d1_hd U415 ( .A(n458), .B(r_add_A[17]), .C(w_mult_Z[17]), .D(n455), .E(
        n34), .F(r_x_data[17]), .Y(n426) );
  scg5d1_hd U416 ( .A(n458), .B(r_add_A[16]), .C(w_mult_Z[16]), .D(n455), .E(
        n34), .F(r_x_data[16]), .Y(n427) );
  scg5d1_hd U417 ( .A(n458), .B(r_add_A[15]), .C(w_mult_Z[15]), .D(n455), .E(
        n34), .F(r_x_data[15]), .Y(n428) );
  scg5d1_hd U418 ( .A(n458), .B(r_add_A[14]), .C(w_mult_Z[14]), .D(n455), .E(
        n34), .F(r_x_data[14]), .Y(n429) );
  scg5d1_hd U419 ( .A(n458), .B(r_add_A[13]), .C(w_mult_Z[13]), .D(n455), .E(
        n34), .F(r_x_data[13]), .Y(n430) );
  scg5d1_hd U420 ( .A(n458), .B(r_add_A[12]), .C(w_mult_Z[12]), .D(n455), .E(
        n34), .F(r_x_data[12]), .Y(n431) );
  scg5d1_hd U421 ( .A(n458), .B(r_add_A[11]), .C(w_mult_Z[11]), .D(n455), .E(
        n34), .F(r_x_data[11]), .Y(n432) );
  scg5d1_hd U422 ( .A(n458), .B(r_add_A[10]), .C(w_mult_Z[10]), .D(n455), .E(
        n34), .F(r_x_data[10]), .Y(n433) );
  scg5d1_hd U423 ( .A(n458), .B(r_add_A[9]), .C(w_mult_Z[9]), .D(n455), .E(n34), .F(r_x_data[9]), .Y(n434) );
  scg5d1_hd U424 ( .A(n458), .B(r_add_A[8]), .C(w_mult_Z[8]), .D(n455), .E(n34), .F(r_x_data[8]), .Y(n435) );
  scg5d1_hd U425 ( .A(n458), .B(r_add_A[7]), .C(w_mult_Z[7]), .D(n455), .E(n34), .F(r_x_data[7]), .Y(n436) );
  scg5d1_hd U426 ( .A(n458), .B(r_add_A[6]), .C(w_mult_Z[6]), .D(n455), .E(n34), .F(r_x_data[6]), .Y(n437) );
  scg5d1_hd U427 ( .A(n458), .B(r_add_A[5]), .C(w_mult_Z[5]), .D(n455), .E(n34), .F(r_x_data[5]), .Y(n438) );
  scg5d1_hd U428 ( .A(n458), .B(r_add_A[4]), .C(w_mult_Z[4]), .D(n455), .E(n34), .F(r_x_data[4]), .Y(n439) );
  scg5d1_hd U429 ( .A(n458), .B(r_add_A[3]), .C(w_mult_Z[3]), .D(n455), .E(n34), .F(r_x_data[3]), .Y(n440) );
  scg5d1_hd U430 ( .A(n458), .B(r_add_A[2]), .C(w_mult_Z[2]), .D(n455), .E(n34), .F(r_x_data[2]), .Y(n441) );
  scg5d1_hd U431 ( .A(n458), .B(r_add_A[1]), .C(w_mult_Z[1]), .D(n455), .E(n34), .F(r_x_data[1]), .Y(n442) );
  scg5d1_hd U442 ( .A(n458), .B(r_add_A[31]), .C(w_mult_Z[31]), .D(n455), .E(
        n34), .F(r_x_data[31]), .Y(n447) );
  scg5d1_hd U443 ( .A(r_add_A[0]), .B(n458), .C(w_mult_Z[0]), .D(n455), .E(n34), .F(r_x_data[0]), .Y(n448) );
  oa211d1_hd U448 ( .A(r_counter_0_), .B(w_add_Z_STB), .C(n221), .D(
        w_mult_Z_STB), .Y(n342) );
  ivd1_hd U456 ( .A(i_RSTN), .Y(N17) );
  fd2qd1_hd r_mult_A_reg_2_ ( .D(n78), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[2]) );
  fd2qd1_hd r_mult_A_reg_3_ ( .D(n77), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[3]) );
  fd2qd1_hd r_mult_A_reg_4_ ( .D(n76), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[4]) );
  fd2qd1_hd r_mult_A_reg_10_ ( .D(n70), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[10]) );
  fd2qd1_hd r_mult_A_reg_12_ ( .D(n68), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[12]) );
  fd2qd1_hd r_mult_A_reg_15_ ( .D(n65), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[15]) );
  fd2qd1_hd r_mult_A_reg_18_ ( .D(n62), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[18]) );
  fd2qd1_hd r_mult_A_reg_19_ ( .D(n61), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[19]) );
  fd2qd1_hd r_mult_A_reg_20_ ( .D(n60), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[20]) );
  fd2qd1_hd r_mult_A_reg_23_ ( .D(n57), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[23]) );
  fd2qd1_hd r_mult_A_reg_30_ ( .D(n50), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[30]) );
  fd2qd1_hd r_mult_A_reg_31_ ( .D(n49), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[31]) );
  fd2qd1_hd r_mult_AB_STB_reg ( .D(n145), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_AB_STB) );
  fd2qd1_hd r_mult_B_reg_31_ ( .D(n214), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[31]) );
  fd2qd1_hd r_mult_B_reg_0_ ( .D(n111), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[0]) );
  fd2qd1_hd r_mult_B_reg_1_ ( .D(n110), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[1]) );
  fd2qd1_hd r_mult_B_reg_2_ ( .D(n109), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[2]) );
  fd2qd1_hd r_mult_B_reg_3_ ( .D(n108), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[3]) );
  fd2qd1_hd r_mult_B_reg_4_ ( .D(n107), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[4]) );
  fd2qd1_hd r_mult_B_reg_5_ ( .D(n106), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[5]) );
  fd2qd1_hd r_mult_B_reg_6_ ( .D(n105), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[6]) );
  fd2qd1_hd r_mult_B_reg_7_ ( .D(n104), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[7]) );
  fd2qd1_hd r_mult_B_reg_8_ ( .D(n103), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[8]) );
  fd2qd1_hd r_mult_B_reg_9_ ( .D(n102), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[9]) );
  fd2qd1_hd r_mult_B_reg_10_ ( .D(n101), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[10]) );
  fd2qd1_hd r_mult_B_reg_11_ ( .D(n100), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[11]) );
  fd2qd1_hd r_mult_B_reg_12_ ( .D(n99), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[12]) );
  fd2qd1_hd r_mult_B_reg_13_ ( .D(n98), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[13]) );
  fd2qd1_hd r_mult_B_reg_14_ ( .D(n97), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[14]) );
  fd2qd1_hd r_mult_B_reg_15_ ( .D(n96), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[15]) );
  fd2qd1_hd r_mult_B_reg_16_ ( .D(n95), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[16]) );
  fd2qd1_hd r_mult_B_reg_17_ ( .D(n94), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[17]) );
  fd2qd1_hd r_mult_B_reg_18_ ( .D(n93), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[18]) );
  fd2qd1_hd r_mult_B_reg_19_ ( .D(n92), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[19]) );
  fd2qd1_hd r_mult_B_reg_20_ ( .D(n91), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[20]) );
  fd2qd1_hd r_mult_B_reg_21_ ( .D(n90), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[21]) );
  fd2qd1_hd r_mult_B_reg_22_ ( .D(n89), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[22]) );
  fd2qd1_hd r_mult_B_reg_23_ ( .D(n88), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[23]) );
  fd2qd1_hd r_mult_B_reg_24_ ( .D(n87), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[24]) );
  fd2qd1_hd r_mult_B_reg_25_ ( .D(n86), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[25]) );
  fd2qd1_hd r_mult_B_reg_26_ ( .D(n85), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[26]) );
  fd2qd1_hd r_mult_B_reg_27_ ( .D(n84), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[27]) );
  fd2qd1_hd r_mult_B_reg_28_ ( .D(n83), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[28]) );
  fd2qd1_hd r_mult_B_reg_29_ ( .D(n82), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[29]) );
  fd2qd1_hd r_mult_B_reg_30_ ( .D(n81), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[30]) );
  fd2qd1_hd r_mult_A_reg_0_ ( .D(n80), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[0]) );
  fd2qd1_hd r_mult_A_reg_1_ ( .D(n79), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[1]) );
  fd2qd1_hd r_mult_A_reg_5_ ( .D(n75), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[5]) );
  fd2qd1_hd r_mult_A_reg_6_ ( .D(n74), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[6]) );
  fd2qd1_hd r_mult_A_reg_7_ ( .D(n73), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[7]) );
  fd2qd1_hd r_mult_A_reg_8_ ( .D(n72), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[8]) );
  fd2qd1_hd r_mult_A_reg_9_ ( .D(n71), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[9]) );
  fd2qd1_hd r_mult_A_reg_11_ ( .D(n69), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[11]) );
  fd2qd1_hd r_mult_A_reg_13_ ( .D(n67), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[13]) );
  fd2qd1_hd r_mult_A_reg_14_ ( .D(n66), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[14]) );
  fd2qd1_hd r_mult_A_reg_16_ ( .D(n64), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[16]) );
  fd2qd1_hd r_mult_A_reg_17_ ( .D(n63), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[17]) );
  fd2qd1_hd r_mult_A_reg_21_ ( .D(n59), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[21]) );
  fd2qd1_hd r_mult_A_reg_22_ ( .D(n58), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[22]) );
  fd2qd1_hd r_mult_A_reg_24_ ( .D(n56), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[24]) );
  fd2qd1_hd r_mult_A_reg_25_ ( .D(n55), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[25]) );
  fd2qd1_hd r_mult_A_reg_26_ ( .D(n54), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[26]) );
  fd2qd1_hd r_mult_A_reg_27_ ( .D(n53), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[27]) );
  fd2qd1_hd r_mult_A_reg_28_ ( .D(n52), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[28]) );
  fd2qd1_hd r_mult_A_reg_29_ ( .D(n51), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[29]) );
  fd2qd1_hd r_mult_Z_ACK_reg ( .D(n144), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_Z_ACK) );
  fd2qd1_hd r_add_A_reg_30_ ( .D(n413), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[30]) );
  fd2qd1_hd r_add_A_reg_29_ ( .D(n414), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[29]) );
  fd2qd1_hd r_add_A_reg_28_ ( .D(n415), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[28]) );
  fd2qd1_hd r_add_A_reg_27_ ( .D(n416), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[27]) );
  fd2qd1_hd r_add_A_reg_26_ ( .D(n417), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[26]) );
  fd2qd1_hd r_add_A_reg_25_ ( .D(n418), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[25]) );
  fd2qd1_hd r_add_A_reg_24_ ( .D(n419), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[24]) );
  fd2qd1_hd r_add_A_reg_23_ ( .D(n420), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[23]) );
  fd2qd1_hd r_add_A_reg_22_ ( .D(n421), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[22]) );
  fd2qd1_hd r_add_A_reg_21_ ( .D(n422), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[21]) );
  fd2qd1_hd r_add_A_reg_20_ ( .D(n423), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[20]) );
  fd2qd1_hd r_add_A_reg_19_ ( .D(n424), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[19]) );
  fd2qd1_hd r_add_A_reg_18_ ( .D(n425), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[18]) );
  fd2qd1_hd r_add_A_reg_17_ ( .D(n426), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[17]) );
  fd2qd1_hd r_add_A_reg_16_ ( .D(n427), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[16]) );
  fd2qd1_hd r_add_A_reg_15_ ( .D(n428), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[15]) );
  fd2qd1_hd r_add_A_reg_14_ ( .D(n429), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[14]) );
  fd2qd1_hd r_add_A_reg_13_ ( .D(n430), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[13]) );
  fd2qd1_hd r_add_A_reg_12_ ( .D(n431), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[12]) );
  fd2qd1_hd r_add_A_reg_11_ ( .D(n432), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[11]) );
  fd2qd1_hd r_add_A_reg_10_ ( .D(n433), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[10]) );
  fd2qd1_hd r_add_A_reg_9_ ( .D(n434), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[9])
         );
  fd2qd1_hd r_add_A_reg_8_ ( .D(n435), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[8])
         );
  fd2qd1_hd r_add_A_reg_7_ ( .D(n436), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[7])
         );
  fd2qd1_hd r_add_A_reg_6_ ( .D(n437), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[6])
         );
  fd2qd1_hd r_add_A_reg_5_ ( .D(n438), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[5])
         );
  fd2qd1_hd r_add_A_reg_4_ ( .D(n439), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[4])
         );
  fd2qd1_hd r_add_A_reg_3_ ( .D(n440), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[3])
         );
  fd2qd1_hd r_add_A_reg_2_ ( .D(n441), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[2])
         );
  fd2qd1_hd r_add_A_reg_1_ ( .D(n442), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[1])
         );
  fd2qd1_hd r_add_A_reg_31_ ( .D(n447), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[31]) );
  fd2qd1_hd r_add_A_reg_0_ ( .D(n448), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[0])
         );
  fd2qd1_hd r_y_data_reg_0_ ( .D(n143), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[0]) );
  fd2qd1_hd r_y_data_reg_1_ ( .D(n142), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[1]) );
  fd2qd1_hd r_y_data_reg_2_ ( .D(n141), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[2]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(n140), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[3]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(n139), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(n138), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(n137), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(n136), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(n135), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(n134), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(n133), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(n132), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(n131), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(n130), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(n129), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(n128), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(n127), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(n126), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(n125), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(n124), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(n123), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(n122), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(n121), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(n120), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(n119), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(n118), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(n117), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(n116), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(n115), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(n114), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(n113), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(n112), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_add_B_reg_31_ ( .D(n348), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[31]) );
  fd2qd1_hd r_add_B_reg_30_ ( .D(n349), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[30]) );
  fd2qd1_hd r_add_B_reg_29_ ( .D(n350), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[29]) );
  fd2qd1_hd r_add_B_reg_28_ ( .D(n351), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[28]) );
  fd2qd1_hd r_add_B_reg_27_ ( .D(n352), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[27]) );
  fd2qd1_hd r_add_B_reg_26_ ( .D(n353), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[26]) );
  fd2qd1_hd r_add_B_reg_25_ ( .D(n354), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[25]) );
  fd2qd1_hd r_add_B_reg_24_ ( .D(n355), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[24]) );
  fd2qd1_hd r_add_B_reg_23_ ( .D(n356), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[23]) );
  fd2qd1_hd r_add_B_reg_22_ ( .D(n357), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[22]) );
  fd2qd1_hd r_add_B_reg_21_ ( .D(n358), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[21]) );
  fd2qd1_hd r_add_B_reg_20_ ( .D(n359), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[20]) );
  fd2qd1_hd r_add_B_reg_19_ ( .D(n360), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[19]) );
  fd2qd1_hd r_add_B_reg_18_ ( .D(n361), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[18]) );
  fd2qd1_hd r_add_B_reg_17_ ( .D(n362), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[17]) );
  fd2qd1_hd r_add_B_reg_16_ ( .D(n363), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[16]) );
  fd2qd1_hd r_add_B_reg_15_ ( .D(n364), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[15]) );
  fd2qd1_hd r_add_B_reg_14_ ( .D(n365), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[14]) );
  fd2qd1_hd r_add_B_reg_13_ ( .D(n366), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[13]) );
  fd2qd1_hd r_add_B_reg_12_ ( .D(n367), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[12]) );
  fd2qd1_hd r_add_B_reg_11_ ( .D(n368), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[11]) );
  fd2qd1_hd r_add_B_reg_10_ ( .D(n369), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[10]) );
  fd2qd1_hd r_add_B_reg_9_ ( .D(n370), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[9])
         );
  fd2qd1_hd r_add_B_reg_8_ ( .D(n371), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[8])
         );
  fd2qd1_hd r_add_B_reg_7_ ( .D(n372), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[7])
         );
  fd2qd1_hd r_add_B_reg_6_ ( .D(n373), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[6])
         );
  fd2qd1_hd r_add_B_reg_5_ ( .D(n374), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[5])
         );
  fd2qd1_hd r_add_B_reg_4_ ( .D(n375), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[4])
         );
  fd2qd1_hd r_add_B_reg_3_ ( .D(n376), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[3])
         );
  fd2qd1_hd r_add_B_reg_2_ ( .D(n377), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[2])
         );
  fd2qd1_hd r_add_B_reg_1_ ( .D(n378), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[1])
         );
  fd2qd1_hd r_add_B_reg_0_ ( .D(n379), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[0])
         );
  fd2qd1_hd r_x_data_reg_32_ ( .D(n177), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[32]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(n176), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(n175), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[34]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(n174), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(n173), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(n172), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[37]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(n171), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(n170), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(n169), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(n168), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(n167), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(n166), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(n165), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(n164), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(n163), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(n162), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(n161), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(n160), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(n159), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(n158), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[51]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(n157), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(n156), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(n155), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(n154), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(n153), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(n152), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(n151), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[58]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(n150), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(n149), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(n148), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(n147), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(n146), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[63]) );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(n411), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[0]) );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(n410), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[1]) );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(n409), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[2]) );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(n408), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[3]) );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(n407), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[4]) );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(n406), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[5]) );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(n405), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[6]) );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(n404), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[7]) );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(n403), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[8]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(n402), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[9]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(n401), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(n400), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(n399), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(n398), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(n397), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(n396), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(n395), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(n394), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(n393), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(n392), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(n391), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(n390), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(n389), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(n388), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(n387), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(n386), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(n385), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(n384), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(n383), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(n382), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(n381), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(n209), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(n208), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(n207), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(n206), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(n205), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(n204), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[5]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(n203), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(n202), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(n201), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(n200), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(n199), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(n198), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(n197), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(n196), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(n195), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(n194), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(n193), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(n192), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(n191), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(n190), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(n189), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(n188), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(n187), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(n186), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(n185), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(n184), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(n183), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(n182), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(n181), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(n180), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(n179), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(n178), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[31]) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(n380), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[31]) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n450), .E(N559), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_add_Z_ACK_reg ( .D(n443), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_Z_ACK) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n444), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_add_AB_STB_reg ( .D(n412), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_AB_STB) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(N553), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_pstate_0_) );
  scg6d1_hd U457 ( .A(n449), .B(n482), .C(n34), .Y(n486) );
  clknd2d1_hd U458 ( .A(n223), .B(n453), .Y(n484) );
  clknd2d1_hd U459 ( .A(w_mult_Z_STB), .B(n221), .Y(n469) );
  clknd2d1_hd U460 ( .A(w_add_AB_ACK), .B(w_mult_AB_ACK), .Y(n471) );
  clknd2d1_hd U461 ( .A(n343), .B(n221), .Y(n470) );
  clknd2d1_hd U462 ( .A(n472), .B(n213), .Y(n474) );
  clknd2d1_hd U463 ( .A(n213), .B(r_pstate_0_), .Y(n481) );
  clknd2d4_hd U464 ( .A(N556), .B(n33), .Y(n460) );
  clknd2d1_hd U465 ( .A(N548), .B(n223), .Y(n480) );
  clknd2d1_hd U466 ( .A(n464), .B(n470), .Y(N548) );
  clknd2d1_hd U467 ( .A(n485), .B(n481), .Y(n475) );
  clknd2d1_hd U468 ( .A(n478), .B(r_add_Z_ACK), .Y(n477) );
  nd2d4_hd U469 ( .A(o_X_DATA_READY), .B(i_X_DATA_VALID), .Y(n450) );
  clknd2d1_hd U470 ( .A(n451), .B(i_X_DATA[31]), .Y(n558) );
  clknd2d1_hd U471 ( .A(n451), .B(i_X_DATA[30]), .Y(n559) );
  clknd2d1_hd U472 ( .A(n451), .B(i_X_DATA[29]), .Y(n560) );
  clknd2d1_hd U473 ( .A(n451), .B(i_X_DATA[28]), .Y(n561) );
  clknd2d1_hd U474 ( .A(n451), .B(i_X_DATA[27]), .Y(n562) );
  clknd2d1_hd U475 ( .A(n451), .B(i_X_DATA[26]), .Y(n563) );
  clknd2d1_hd U476 ( .A(n451), .B(i_X_DATA[25]), .Y(n564) );
  clknd2d1_hd U477 ( .A(n451), .B(i_X_DATA[24]), .Y(n565) );
  clknd2d1_hd U478 ( .A(n451), .B(i_X_DATA[23]), .Y(n566) );
  clknd2d1_hd U479 ( .A(n451), .B(i_X_DATA[22]), .Y(n567) );
  clknd2d1_hd U480 ( .A(n451), .B(i_X_DATA[21]), .Y(n568) );
  clknd2d1_hd U481 ( .A(n451), .B(i_X_DATA[20]), .Y(n569) );
  clknd2d1_hd U482 ( .A(n451), .B(i_X_DATA[19]), .Y(n570) );
  clknd2d1_hd U483 ( .A(n451), .B(i_X_DATA[18]), .Y(n571) );
  clknd2d1_hd U484 ( .A(n451), .B(i_X_DATA[17]), .Y(n572) );
  clknd2d1_hd U485 ( .A(n451), .B(i_X_DATA[16]), .Y(n573) );
  clknd2d1_hd U486 ( .A(n451), .B(i_X_DATA[15]), .Y(n574) );
  clknd2d1_hd U487 ( .A(n451), .B(i_X_DATA[14]), .Y(n575) );
  clknd2d1_hd U488 ( .A(n451), .B(i_X_DATA[13]), .Y(n576) );
  clknd2d1_hd U489 ( .A(n451), .B(i_X_DATA[12]), .Y(n577) );
  clknd2d1_hd U490 ( .A(n451), .B(i_X_DATA[11]), .Y(n578) );
  clknd2d1_hd U491 ( .A(n451), .B(i_X_DATA[10]), .Y(n579) );
  clknd2d1_hd U492 ( .A(n451), .B(i_X_DATA[9]), .Y(n580) );
  clknd2d1_hd U493 ( .A(n451), .B(i_X_DATA[8]), .Y(n581) );
  clknd2d1_hd U494 ( .A(n451), .B(i_X_DATA[7]), .Y(n582) );
  clknd2d1_hd U495 ( .A(n451), .B(i_X_DATA[6]), .Y(n583) );
  clknd2d1_hd U496 ( .A(n451), .B(i_X_DATA[5]), .Y(n584) );
  clknd2d1_hd U497 ( .A(n451), .B(i_X_DATA[4]), .Y(n585) );
  clknd2d1_hd U498 ( .A(n451), .B(i_X_DATA[3]), .Y(n586) );
  clknd2d1_hd U499 ( .A(n451), .B(i_X_DATA[2]), .Y(n587) );
  clknd2d1_hd U500 ( .A(n451), .B(i_X_DATA[1]), .Y(n588) );
  clknd2d1_hd U501 ( .A(n451), .B(i_X_DATA[0]), .Y(n589) );
  nid2_hd U502 ( .A(n295), .Y(n456) );
  ivd6_hd U503 ( .A(n450), .Y(n451) );
  nr2bd2_hd U504 ( .AN(n483), .B(n484), .Y(n294) );
  nd2bd1_hd U505 ( .AN(r_mult_A[29]), .B(n462), .Y(n51) );
  nd2bd1_hd U506 ( .AN(r_mult_A[28]), .B(n462), .Y(n52) );
  nd2bd1_hd U507 ( .AN(r_mult_A[27]), .B(n462), .Y(n53) );
  nd2bd1_hd U508 ( .AN(r_mult_A[9]), .B(n462), .Y(n71) );
  nd2bd1_hd U509 ( .AN(r_mult_A[11]), .B(n462), .Y(n69) );
  nd2bd1_hd U510 ( .AN(r_mult_A[26]), .B(n462), .Y(n54) );
  nd2bd1_hd U511 ( .AN(r_mult_A[7]), .B(n462), .Y(n73) );
  nd2bd1_hd U512 ( .AN(r_mult_A[13]), .B(n462), .Y(n67) );
  nd2bd1_hd U513 ( .AN(r_mult_A[24]), .B(n462), .Y(n56) );
  nd2bd1_hd U514 ( .AN(r_mult_A[25]), .B(n462), .Y(n55) );
  nd2bd1_hd U515 ( .AN(r_mult_A[1]), .B(n462), .Y(n79) );
  nd2bd1_hd U516 ( .AN(r_mult_A[0]), .B(n462), .Y(n80) );
  nd2bd1_hd U517 ( .AN(r_mult_A[22]), .B(n462), .Y(n58) );
  nd2bd1_hd U518 ( .AN(r_mult_A[21]), .B(n462), .Y(n59) );
  nd2bd1_hd U519 ( .AN(r_mult_A[8]), .B(n462), .Y(n72) );
  nd2bd1_hd U520 ( .AN(r_mult_A[17]), .B(n462), .Y(n63) );
  nd2bd1_hd U521 ( .AN(r_mult_A[16]), .B(n462), .Y(n64) );
  nd2bd1_hd U522 ( .AN(r_mult_A[6]), .B(n462), .Y(n74) );
  nd2bd1_hd U523 ( .AN(r_mult_A[14]), .B(n462), .Y(n66) );
  nd2bd1_hd U524 ( .AN(r_mult_A[5]), .B(n462), .Y(n75) );
  nr2d2_hd U525 ( .A(n461), .B(n34), .Y(n462) );
  ivd1_hd U526 ( .A(n34), .Y(n452) );
  ad2d1_hd U527 ( .A(n449), .B(n36), .Y(n548) );
  scg10d1_hd U528 ( .A(n450), .B(r_x_data[2]), .C(r_x_data[34]), .D(n451), .Y(
        n175) );
  scg10d1_hd U529 ( .A(n450), .B(r_x_data[6]), .C(r_x_data[38]), .D(n451), .Y(
        n171) );
  scg10d1_hd U530 ( .A(n450), .B(r_x_data[3]), .C(r_x_data[35]), .D(n451), .Y(
        n174) );
  scg10d1_hd U531 ( .A(n450), .B(r_x_data[7]), .C(r_x_data[39]), .D(n451), .Y(
        n170) );
  scg10d1_hd U532 ( .A(n450), .B(r_x_data[4]), .C(r_x_data[36]), .D(n451), .Y(
        n173) );
  scg10d1_hd U533 ( .A(n450), .B(o_Y_DATA[30]), .C(r_y_data[30]), .D(n451), 
        .Y(n113) );
  scg10d1_hd U534 ( .A(n450), .B(r_x_data[8]), .C(r_x_data[40]), .D(n451), .Y(
        n169) );
  scg10d1_hd U535 ( .A(n450), .B(o_Y_DATA[31]), .C(r_y_data[31]), .D(n451), 
        .Y(n112) );
  scg10d1_hd U536 ( .A(n450), .B(r_x_data[5]), .C(r_x_data[37]), .D(n451), .Y(
        n172) );
  scg10d1_hd U537 ( .A(n450), .B(r_x_data[9]), .C(r_x_data[41]), .D(n451), .Y(
        n168) );
  scg10d1_hd U538 ( .A(n450), .B(r_x_data[0]), .C(r_x_data[32]), .D(n451), .Y(
        n177) );
  scg10d1_hd U539 ( .A(n450), .B(r_x_data[1]), .C(r_x_data[33]), .D(n451), .Y(
        n176) );
  scg10d1_hd U540 ( .A(n450), .B(r_x_data[23]), .C(r_x_data[55]), .D(n451), 
        .Y(n154) );
  scg10d1_hd U541 ( .A(n450), .B(r_x_data[10]), .C(r_x_data[42]), .D(n451), 
        .Y(n167) );
  scg10d1_hd U542 ( .A(n450), .B(r_x_data[11]), .C(r_x_data[43]), .D(n451), 
        .Y(n166) );
  scg10d1_hd U543 ( .A(n450), .B(r_x_data[12]), .C(r_x_data[44]), .D(n451), 
        .Y(n165) );
  scg10d1_hd U544 ( .A(n450), .B(r_x_data[13]), .C(r_x_data[45]), .D(n451), 
        .Y(n164) );
  scg10d1_hd U545 ( .A(n450), .B(r_x_data[14]), .C(r_x_data[46]), .D(n451), 
        .Y(n163) );
  scg10d1_hd U546 ( .A(n450), .B(r_x_data[15]), .C(r_x_data[47]), .D(n451), 
        .Y(n162) );
  scg10d1_hd U547 ( .A(n450), .B(r_x_data[16]), .C(r_x_data[48]), .D(n451), 
        .Y(n161) );
  scg10d1_hd U548 ( .A(n450), .B(r_x_data[17]), .C(r_x_data[49]), .D(n451), 
        .Y(n160) );
  scg10d1_hd U549 ( .A(n450), .B(r_x_data[18]), .C(r_x_data[50]), .D(n451), 
        .Y(n159) );
  scg10d1_hd U550 ( .A(n450), .B(r_x_data[19]), .C(r_x_data[51]), .D(n451), 
        .Y(n158) );
  scg10d1_hd U551 ( .A(n450), .B(r_x_data[20]), .C(r_x_data[52]), .D(n451), 
        .Y(n157) );
  scg10d1_hd U552 ( .A(n450), .B(r_x_data[21]), .C(r_x_data[53]), .D(n451), 
        .Y(n156) );
  scg10d1_hd U553 ( .A(n450), .B(r_x_data[22]), .C(r_x_data[54]), .D(n451), 
        .Y(n155) );
  scg10d1_hd U554 ( .A(n450), .B(r_x_data[24]), .C(r_x_data[56]), .D(n451), 
        .Y(n153) );
  scg10d1_hd U555 ( .A(n450), .B(r_x_data[25]), .C(r_x_data[57]), .D(n451), 
        .Y(n152) );
  scg10d1_hd U556 ( .A(n450), .B(r_x_data[26]), .C(r_x_data[58]), .D(n451), 
        .Y(n151) );
  scg10d1_hd U557 ( .A(n450), .B(r_x_data[27]), .C(r_x_data[59]), .D(n451), 
        .Y(n150) );
  scg10d1_hd U558 ( .A(n450), .B(r_x_data[28]), .C(r_x_data[60]), .D(n451), 
        .Y(n149) );
  scg10d1_hd U559 ( .A(n450), .B(r_x_data[29]), .C(r_x_data[61]), .D(n451), 
        .Y(n148) );
  scg10d1_hd U560 ( .A(n450), .B(r_x_data[30]), .C(r_x_data[62]), .D(n451), 
        .Y(n147) );
  scg10d1_hd U561 ( .A(n450), .B(r_x_data[31]), .C(r_x_data[63]), .D(n451), 
        .Y(n146) );
  scg10d1_hd U562 ( .A(n450), .B(o_Y_DATA[0]), .C(r_y_data[0]), .D(n451), .Y(
        n143) );
  scg10d1_hd U563 ( .A(n450), .B(o_Y_DATA[1]), .C(r_y_data[1]), .D(n451), .Y(
        n142) );
  scg10d1_hd U564 ( .A(n450), .B(o_Y_DATA[2]), .C(r_y_data[2]), .D(n451), .Y(
        n141) );
  scg10d1_hd U565 ( .A(n450), .B(o_Y_DATA[4]), .C(r_y_data[4]), .D(n451), .Y(
        n139) );
  scg10d1_hd U566 ( .A(n450), .B(o_Y_DATA[5]), .C(r_y_data[5]), .D(n451), .Y(
        n138) );
  scg10d1_hd U567 ( .A(n450), .B(o_Y_DATA[6]), .C(r_y_data[6]), .D(n451), .Y(
        n137) );
  scg10d1_hd U568 ( .A(n450), .B(o_Y_DATA[7]), .C(r_y_data[7]), .D(n451), .Y(
        n136) );
  scg10d1_hd U569 ( .A(n450), .B(o_Y_DATA[8]), .C(r_y_data[8]), .D(n451), .Y(
        n135) );
  scg10d1_hd U570 ( .A(n450), .B(o_Y_DATA[9]), .C(r_y_data[9]), .D(n451), .Y(
        n134) );
  scg10d1_hd U571 ( .A(n450), .B(o_Y_DATA[10]), .C(r_y_data[10]), .D(n451), 
        .Y(n133) );
  scg10d1_hd U572 ( .A(n450), .B(o_Y_DATA[11]), .C(r_y_data[11]), .D(n451), 
        .Y(n132) );
  scg10d1_hd U573 ( .A(n450), .B(o_Y_DATA[12]), .C(r_y_data[12]), .D(n451), 
        .Y(n131) );
  scg10d1_hd U574 ( .A(n450), .B(o_Y_DATA[13]), .C(r_y_data[13]), .D(n451), 
        .Y(n130) );
  scg10d1_hd U575 ( .A(n450), .B(o_Y_DATA[14]), .C(r_y_data[14]), .D(n451), 
        .Y(n129) );
  scg10d1_hd U576 ( .A(n450), .B(o_Y_DATA[15]), .C(r_y_data[15]), .D(n451), 
        .Y(n128) );
  scg10d1_hd U577 ( .A(n450), .B(o_Y_DATA[16]), .C(r_y_data[16]), .D(n451), 
        .Y(n127) );
  scg10d1_hd U578 ( .A(n450), .B(o_Y_DATA[17]), .C(r_y_data[17]), .D(n451), 
        .Y(n126) );
  scg10d1_hd U579 ( .A(n450), .B(o_Y_DATA[18]), .C(r_y_data[18]), .D(n451), 
        .Y(n125) );
  scg10d1_hd U580 ( .A(n450), .B(o_Y_DATA[28]), .C(r_y_data[28]), .D(n451), 
        .Y(n115) );
  scg10d1_hd U581 ( .A(n450), .B(o_Y_DATA[26]), .C(r_y_data[26]), .D(n451), 
        .Y(n117) );
  scg10d1_hd U582 ( .A(n450), .B(o_Y_DATA[22]), .C(r_y_data[22]), .D(n451), 
        .Y(n121) );
  scg10d1_hd U583 ( .A(n450), .B(o_Y_DATA[19]), .C(r_y_data[19]), .D(n451), 
        .Y(n124) );
  scg10d1_hd U584 ( .A(n450), .B(o_Y_DATA[24]), .C(r_y_data[24]), .D(n451), 
        .Y(n119) );
  scg10d1_hd U585 ( .A(n450), .B(o_Y_DATA[3]), .C(r_y_data[3]), .D(n451), .Y(
        n140) );
  scg10d1_hd U586 ( .A(n450), .B(o_Y_DATA[20]), .C(r_y_data[20]), .D(n451), 
        .Y(n123) );
  scg10d1_hd U587 ( .A(n450), .B(o_Y_DATA[21]), .C(r_y_data[21]), .D(n451), 
        .Y(n122) );
  scg10d1_hd U588 ( .A(n450), .B(o_Y_DATA[23]), .C(r_y_data[23]), .D(n451), 
        .Y(n120) );
  scg10d1_hd U589 ( .A(n450), .B(o_Y_DATA[25]), .C(r_y_data[25]), .D(n451), 
        .Y(n118) );
  scg10d1_hd U590 ( .A(n450), .B(o_Y_DATA[27]), .C(r_y_data[27]), .D(n451), 
        .Y(n116) );
  scg10d1_hd U591 ( .A(n450), .B(o_Y_DATA[29]), .C(r_y_data[29]), .D(n451), 
        .Y(n114) );
  nid6_hd U592 ( .A(n459), .Y(n34) );
  nid2_hd U593 ( .A(n486), .Y(n453) );
  nid2_hd U594 ( .A(n548), .Y(n455) );
  scg14d1_hd U595 ( .A(n463), .B(n341), .C(n481), .Y(n36) );
  ivd1_hd U596 ( .A(n485), .Y(n463) );
  nr3d1_hd U597 ( .A(n555), .B(n485), .C(n484), .Y(n295) );
  nid2_hd U598 ( .A(n294), .Y(n457) );
  ivd1_hd U599 ( .A(n449), .Y(n485) );
  nid4_hd U600 ( .A(n260), .Y(n458) );
  nd2d1_hd U601 ( .A(n36), .B(n33), .Y(n260) );
  ivd2_hd U602 ( .A(n548), .Y(n454) );
  nr2d1_hd U603 ( .A(r_counter_0_), .B(n470), .Y(n459) );
  nr2d1_hd U604 ( .A(n481), .B(n471), .Y(n343) );
  ivd1_hd U605 ( .A(w_add_Z_STB), .Y(n215) );
  ivd1_hd U606 ( .A(n223), .Y(r_counter_0_) );
  nr2d1_hd U607 ( .A(n213), .B(r_pstate_0_), .Y(n449) );
  scg6d1_hd U608 ( .A(o_Y_DATA_VALID), .B(n475), .C(n551), .Y(n444) );
  ivd1_hd U609 ( .A(n481), .Y(n466) );
  ivd1_hd U610 ( .A(n471), .Y(n35) );
  ivd1_hd U611 ( .A(o_Y_DATA[13]), .Y(n514) );
  ivd1_hd U612 ( .A(o_Y_DATA[17]), .Y(n522) );
  ivd1_hd U613 ( .A(o_Y_DATA[16]), .Y(n520) );
  ivd1_hd U614 ( .A(o_Y_DATA[15]), .Y(n518) );
  ivd1_hd U615 ( .A(o_Y_DATA[14]), .Y(n516) );
  ivd1_hd U616 ( .A(o_Y_DATA[26]), .Y(n540) );
  ivd1_hd U617 ( .A(o_Y_DATA[25]), .Y(n538) );
  ivd1_hd U618 ( .A(o_Y_DATA[29]), .Y(n546) );
  ivd1_hd U619 ( .A(o_Y_DATA[28]), .Y(n544) );
  ivd1_hd U620 ( .A(o_Y_DATA[27]), .Y(n542) );
  ivd1_hd U621 ( .A(o_Y_DATA[21]), .Y(n530) );
  ivd1_hd U622 ( .A(o_Y_DATA[20]), .Y(n528) );
  ivd1_hd U623 ( .A(o_Y_DATA[24]), .Y(n536) );
  ivd1_hd U624 ( .A(o_Y_DATA[22]), .Y(n532) );
  ivd1_hd U625 ( .A(o_Y_DATA[12]), .Y(n512) );
  ivd1_hd U626 ( .A(o_Y_DATA[19]), .Y(n526) );
  ivd1_hd U627 ( .A(o_Y_DATA[18]), .Y(n524) );
  ivd1_hd U628 ( .A(o_Y_DATA[30]), .Y(n549) );
  ivd1_hd U629 ( .A(o_Y_DATA[0]), .Y(n488) );
  ivd1_hd U630 ( .A(o_Y_DATA[7]), .Y(n502) );
  ivd1_hd U631 ( .A(o_Y_DATA[5]), .Y(n498) );
  ivd1_hd U632 ( .A(o_Y_DATA[2]), .Y(n492) );
  ivd1_hd U633 ( .A(o_Y_DATA[1]), .Y(n490) );
  ivd1_hd U634 ( .A(o_Y_DATA[4]), .Y(n496) );
  ivd1_hd U635 ( .A(o_Y_DATA[3]), .Y(n494) );
  ivd1_hd U636 ( .A(o_Y_DATA[6]), .Y(n500) );
  ivd1_hd U637 ( .A(o_Y_DATA[23]), .Y(n534) );
  ivd1_hd U638 ( .A(o_Y_DATA[11]), .Y(n510) );
  ivd1_hd U639 ( .A(o_Y_DATA[9]), .Y(n506) );
  ivd1_hd U640 ( .A(o_Y_DATA[10]), .Y(n508) );
  ivd1_hd U641 ( .A(n221), .Y(n555) );
  ivd1_hd U642 ( .A(o_Y_DATA[8]), .Y(n504) );
  ao211d1_hd U643 ( .A(n221), .B(n346), .C(r_counter_0_), .D(n215), .Y(n482)
         );
  ivd1_hd U644 ( .A(w_mult_Z_STB), .Y(n346) );
  scg22d1_hd U645 ( .A(n221), .B(n35), .C(r_counter_0_), .D(n466), .Y(n33) );
  nr2d1_hd U646 ( .A(n469), .B(n223), .Y(n341) );
  nr2d1_hd U647 ( .A(n221), .B(n485), .Y(n483) );
  scg22d1_hd U648 ( .A(n468), .B(n463), .C(r_counter_0_), .D(n481), .Y(N556)
         );
  ad2d2_hd U649 ( .A(N556), .B(n463), .Y(n461) );
  scg2d1_hd U650 ( .A(n481), .B(r_mult_Z_ACK), .C(n463), .D(n467), .Y(n144) );
  scg5d1_hd U651 ( .A(n460), .B(r_mult_B[12]), .C(n34), .D(r_y_data[12]), .E(
        n461), .F(w_add_Z[12]), .Y(n99) );
  scg5d1_hd U652 ( .A(n460), .B(r_mult_B[13]), .C(n34), .D(r_y_data[13]), .E(
        n461), .F(w_add_Z[13]), .Y(n98) );
  scg5d1_hd U653 ( .A(n460), .B(r_mult_B[14]), .C(n34), .D(r_y_data[14]), .E(
        n461), .F(w_add_Z[14]), .Y(n97) );
  scg5d1_hd U654 ( .A(n460), .B(r_mult_B[15]), .C(n34), .D(r_y_data[15]), .E(
        n461), .F(w_add_Z[15]), .Y(n96) );
  scg5d1_hd U655 ( .A(n460), .B(r_mult_B[16]), .C(n34), .D(r_y_data[16]), .E(
        n461), .F(w_add_Z[16]), .Y(n95) );
  scg5d1_hd U656 ( .A(n460), .B(r_mult_B[17]), .C(n34), .D(r_y_data[17]), .E(
        n461), .F(w_add_Z[17]), .Y(n94) );
  scg5d1_hd U657 ( .A(n460), .B(r_mult_B[18]), .C(n34), .D(r_y_data[18]), .E(
        n461), .F(w_add_Z[18]), .Y(n93) );
  scg5d1_hd U658 ( .A(n460), .B(r_mult_B[19]), .C(n34), .D(r_y_data[19]), .E(
        n461), .F(w_add_Z[19]), .Y(n92) );
  scg5d1_hd U659 ( .A(n460), .B(r_mult_B[20]), .C(n34), .D(r_y_data[20]), .E(
        n461), .F(w_add_Z[20]), .Y(n91) );
  scg5d1_hd U660 ( .A(n460), .B(r_mult_B[21]), .C(n34), .D(r_y_data[21]), .E(
        n461), .F(w_add_Z[21]), .Y(n90) );
  scg5d1_hd U661 ( .A(n460), .B(r_mult_B[22]), .C(n34), .D(r_y_data[22]), .E(
        n461), .F(w_add_Z[22]), .Y(n89) );
  scg5d1_hd U662 ( .A(n460), .B(r_mult_B[23]), .C(n34), .D(r_y_data[23]), .E(
        n461), .F(w_add_Z[23]), .Y(n88) );
  scg5d1_hd U663 ( .A(n460), .B(r_mult_B[24]), .C(n34), .D(r_y_data[24]), .E(
        n461), .F(w_add_Z[24]), .Y(n87) );
  scg5d1_hd U664 ( .A(n460), .B(r_mult_B[25]), .C(n34), .D(r_y_data[25]), .E(
        n461), .F(w_add_Z[25]), .Y(n86) );
  scg5d1_hd U665 ( .A(n460), .B(r_mult_B[26]), .C(n34), .D(r_y_data[26]), .E(
        n461), .F(w_add_Z[26]), .Y(n85) );
  scg5d1_hd U666 ( .A(n460), .B(r_mult_B[27]), .C(n34), .D(r_y_data[27]), .E(
        n461), .F(w_add_Z[27]), .Y(n84) );
  scg5d1_hd U667 ( .A(n460), .B(r_mult_B[28]), .C(n34), .D(r_y_data[28]), .E(
        n461), .F(w_add_Z[28]), .Y(n83) );
  scg5d1_hd U668 ( .A(n460), .B(r_mult_B[29]), .C(n34), .D(r_y_data[29]), .E(
        n461), .F(w_add_Z[29]), .Y(n82) );
  scg5d1_hd U669 ( .A(n460), .B(r_mult_B[30]), .C(n34), .D(r_y_data[30]), .E(
        n461), .F(w_add_Z[30]), .Y(n81) );
  ad2d1_hd U670 ( .A(r_mult_A[2]), .B(n460), .Y(n78) );
  ad2d1_hd U671 ( .A(r_mult_A[3]), .B(n460), .Y(n77) );
  ad2d1_hd U672 ( .A(r_mult_A[4]), .B(n460), .Y(n76) );
  ad2d1_hd U673 ( .A(r_mult_A[10]), .B(n460), .Y(n70) );
  ad2d1_hd U674 ( .A(r_mult_A[12]), .B(n460), .Y(n68) );
  ad2d1_hd U675 ( .A(r_mult_A[15]), .B(n460), .Y(n65) );
  ad2d1_hd U676 ( .A(r_mult_A[18]), .B(n460), .Y(n62) );
  ad2d1_hd U677 ( .A(r_mult_A[19]), .B(n460), .Y(n61) );
  ad2d1_hd U678 ( .A(r_mult_A[20]), .B(n460), .Y(n60) );
  ad2d1_hd U679 ( .A(r_mult_A[23]), .B(n460), .Y(n57) );
  ad2d1_hd U680 ( .A(r_mult_A[30]), .B(n460), .Y(n50) );
  ad2d1_hd U681 ( .A(r_mult_A[31]), .B(n460), .Y(n49) );
  scg5d1_hd U682 ( .A(n460), .B(r_mult_B[31]), .C(n34), .D(r_y_data[31]), .E(
        n461), .F(w_add_Z[31]), .Y(n214) );
  scg14d1_hd U683 ( .A(r_mult_AB_STB), .B(n464), .C(n465), .Y(n145) );
  oa211d1_hd U684 ( .A(n35), .B(n463), .C(n466), .D(n221), .Y(n465) );
  scg13d1_hd U685 ( .A(n468), .B(n341), .C(n481), .Y(n467) );
  scg5d1_hd U686 ( .A(n460), .B(r_mult_B[0]), .C(n34), .D(r_y_data[0]), .E(
        n461), .F(w_add_Z[0]), .Y(n111) );
  scg5d1_hd U687 ( .A(n460), .B(r_mult_B[1]), .C(n34), .D(r_y_data[1]), .E(
        n461), .F(w_add_Z[1]), .Y(n110) );
  scg5d1_hd U688 ( .A(n460), .B(r_mult_B[2]), .C(n34), .D(r_y_data[2]), .E(
        n461), .F(w_add_Z[2]), .Y(n109) );
  scg5d1_hd U689 ( .A(n460), .B(r_mult_B[3]), .C(n34), .D(r_y_data[3]), .E(
        n461), .F(w_add_Z[3]), .Y(n108) );
  scg5d1_hd U690 ( .A(n460), .B(r_mult_B[4]), .C(n34), .D(r_y_data[4]), .E(
        n461), .F(w_add_Z[4]), .Y(n107) );
  scg5d1_hd U691 ( .A(n460), .B(r_mult_B[5]), .C(n34), .D(r_y_data[5]), .E(
        n461), .F(w_add_Z[5]), .Y(n106) );
  scg5d1_hd U692 ( .A(n460), .B(r_mult_B[6]), .C(n34), .D(r_y_data[6]), .E(
        n461), .F(w_add_Z[6]), .Y(n105) );
  scg5d1_hd U693 ( .A(n460), .B(r_mult_B[7]), .C(n34), .D(r_y_data[7]), .E(
        n461), .F(w_add_Z[7]), .Y(n104) );
  scg5d1_hd U694 ( .A(n460), .B(r_mult_B[8]), .C(n34), .D(r_y_data[8]), .E(
        n461), .F(w_add_Z[8]), .Y(n103) );
  scg5d1_hd U695 ( .A(n460), .B(r_mult_B[9]), .C(n34), .D(r_y_data[9]), .E(
        n461), .F(w_add_Z[9]), .Y(n102) );
  scg5d1_hd U696 ( .A(n460), .B(r_mult_B[10]), .C(n34), .D(r_y_data[10]), .E(
        n461), .F(w_add_Z[10]), .Y(n101) );
  scg5d1_hd U697 ( .A(n460), .B(r_mult_B[11]), .C(n34), .D(r_y_data[11]), .E(
        n461), .F(w_add_Z[11]), .Y(n100) );
  nr2d1_hd U698 ( .A(n469), .B(n215), .Y(n468) );
  ao21d1_hd U699 ( .A(n343), .B(n223), .C(n463), .Y(n464) );
  ivd1_hd U700 ( .A(r_pstate_0_), .Y(n472) );
  ivd1_hd U701 ( .A(n474), .Y(n553) );
  oa21d1_hd U702 ( .A(n341), .B(n482), .C(n449), .Y(n552) );
  ivd1_hd U703 ( .A(n552), .Y(n554) );
  ao211d1_hd U704 ( .A(i_Y_ACK), .B(o_Y_DATA_VALID), .C(n213), .D(n472), .Y(
        n551) );
  ao211d1_hd U705 ( .A(n553), .B(n451), .C(n554), .D(n551), .Y(n473) );
  oa21d1_hd U706 ( .A(n35), .B(n481), .C(n473), .Y(N553) );
  nr2d1_hd U707 ( .A(N17), .B(n474), .Y(N559) );
  nr2d1_hd U708 ( .A(r_counter_0_), .B(n215), .Y(n476) );
  ao21d1_hd U709 ( .A(n476), .B(n483), .C(N556), .Y(n478) );
  oa21d1_hd U710 ( .A(n485), .B(n478), .C(n477), .Y(n443) );
  ivd1_hd U711 ( .A(r_add_AB_STB), .Y(n479) );
  oa22d1_hd U712 ( .A(n481), .B(n480), .C(N548), .D(n479), .Y(n412) );
  oa21d1_hd U713 ( .A(n488), .B(n453), .C(n326), .Y(n411) );
  oa21d1_hd U714 ( .A(n453), .B(n490), .C(n325), .Y(n410) );
  oa21d1_hd U715 ( .A(n453), .B(n492), .C(n324), .Y(n409) );
  oa21d1_hd U716 ( .A(n453), .B(n494), .C(n323), .Y(n408) );
  oa21d1_hd U717 ( .A(n453), .B(n496), .C(n322), .Y(n407) );
  oa21d1_hd U718 ( .A(n453), .B(n498), .C(n321), .Y(n406) );
  oa21d1_hd U719 ( .A(n453), .B(n500), .C(n320), .Y(n405) );
  oa21d1_hd U720 ( .A(n453), .B(n502), .C(n319), .Y(n404) );
  oa21d1_hd U721 ( .A(n486), .B(n504), .C(n318), .Y(n403) );
  oa21d1_hd U722 ( .A(n486), .B(n506), .C(n317), .Y(n402) );
  oa21d1_hd U723 ( .A(n486), .B(n508), .C(n316), .Y(n401) );
  oa21d1_hd U724 ( .A(n486), .B(n510), .C(n315), .Y(n400) );
  oa21d1_hd U725 ( .A(n486), .B(n512), .C(n314), .Y(n399) );
  oa21d1_hd U726 ( .A(n486), .B(n514), .C(n313), .Y(n398) );
  oa21d1_hd U727 ( .A(n486), .B(n516), .C(n312), .Y(n397) );
  oa21d1_hd U728 ( .A(n486), .B(n518), .C(n311), .Y(n396) );
  oa21d1_hd U729 ( .A(n486), .B(n520), .C(n310), .Y(n395) );
  oa21d1_hd U730 ( .A(n486), .B(n522), .C(n309), .Y(n394) );
  oa21d1_hd U731 ( .A(n486), .B(n524), .C(n308), .Y(n393) );
  oa21d1_hd U732 ( .A(n453), .B(n526), .C(n307), .Y(n392) );
  oa21d1_hd U733 ( .A(n453), .B(n528), .C(n306), .Y(n391) );
  oa21d1_hd U734 ( .A(n453), .B(n530), .C(n305), .Y(n390) );
  oa21d1_hd U735 ( .A(n453), .B(n532), .C(n304), .Y(n389) );
  oa21d1_hd U736 ( .A(n486), .B(n534), .C(n303), .Y(n388) );
  oa21d1_hd U737 ( .A(n453), .B(n536), .C(n302), .Y(n387) );
  oa21d1_hd U738 ( .A(n453), .B(n538), .C(n301), .Y(n386) );
  oa21d1_hd U739 ( .A(n453), .B(n540), .C(n300), .Y(n385) );
  oa21d1_hd U740 ( .A(n453), .B(n542), .C(n299), .Y(n384) );
  oa21d1_hd U741 ( .A(n453), .B(n544), .C(n298), .Y(n383) );
  oa21d1_hd U742 ( .A(n453), .B(n546), .C(n297), .Y(n382) );
  oa21d1_hd U743 ( .A(n453), .B(n549), .C(n296), .Y(n381) );
  scg16d1_hd U744 ( .A(o_Y_DATA[31]), .B(n453), .C(n293), .Y(n380) );
  ao22d1_hd U745 ( .A(n34), .B(r_x_data[32]), .C(r_add_B[0]), .D(n458), .Y(
        n487) );
  oa21d1_hd U746 ( .A(n488), .B(n454), .C(n487), .Y(n379) );
  ao22d1_hd U747 ( .A(n34), .B(r_x_data[33]), .C(r_add_B[1]), .D(n260), .Y(
        n489) );
  oa21d1_hd U748 ( .A(n490), .B(n454), .C(n489), .Y(n378) );
  ao22d1_hd U749 ( .A(n34), .B(r_x_data[34]), .C(r_add_B[2]), .D(n260), .Y(
        n491) );
  oa21d1_hd U750 ( .A(n492), .B(n454), .C(n491), .Y(n377) );
  ao22d1_hd U751 ( .A(n34), .B(r_x_data[35]), .C(r_add_B[3]), .D(n260), .Y(
        n493) );
  oa21d1_hd U752 ( .A(n494), .B(n454), .C(n493), .Y(n376) );
  ao22d1_hd U753 ( .A(n34), .B(r_x_data[36]), .C(r_add_B[4]), .D(n260), .Y(
        n495) );
  oa21d1_hd U754 ( .A(n496), .B(n454), .C(n495), .Y(n375) );
  ao22d1_hd U755 ( .A(n34), .B(r_x_data[37]), .C(r_add_B[5]), .D(n260), .Y(
        n497) );
  oa21d1_hd U756 ( .A(n498), .B(n454), .C(n497), .Y(n374) );
  ao22d1_hd U757 ( .A(n34), .B(r_x_data[38]), .C(r_add_B[6]), .D(n260), .Y(
        n499) );
  oa21d1_hd U758 ( .A(n500), .B(n454), .C(n499), .Y(n373) );
  ao22d1_hd U759 ( .A(n34), .B(r_x_data[39]), .C(r_add_B[7]), .D(n260), .Y(
        n501) );
  oa21d1_hd U760 ( .A(n502), .B(n454), .C(n501), .Y(n372) );
  ao22d1_hd U761 ( .A(n34), .B(r_x_data[40]), .C(r_add_B[8]), .D(n260), .Y(
        n503) );
  oa21d1_hd U762 ( .A(n504), .B(n454), .C(n503), .Y(n371) );
  ao22d1_hd U763 ( .A(n34), .B(r_x_data[41]), .C(r_add_B[9]), .D(n260), .Y(
        n505) );
  oa21d1_hd U764 ( .A(n506), .B(n454), .C(n505), .Y(n370) );
  ao22d1_hd U765 ( .A(n34), .B(r_x_data[42]), .C(r_add_B[10]), .D(n458), .Y(
        n507) );
  oa21d1_hd U766 ( .A(n508), .B(n454), .C(n507), .Y(n369) );
  ao22d1_hd U767 ( .A(n34), .B(r_x_data[43]), .C(r_add_B[11]), .D(n458), .Y(
        n509) );
  oa21d1_hd U768 ( .A(n510), .B(n454), .C(n509), .Y(n368) );
  ao22d1_hd U769 ( .A(n34), .B(r_x_data[44]), .C(r_add_B[12]), .D(n458), .Y(
        n511) );
  oa21d1_hd U770 ( .A(n512), .B(n454), .C(n511), .Y(n367) );
  ao22d1_hd U771 ( .A(n34), .B(r_x_data[45]), .C(r_add_B[13]), .D(n458), .Y(
        n513) );
  oa21d1_hd U772 ( .A(n514), .B(n454), .C(n513), .Y(n366) );
  ao22d1_hd U773 ( .A(n34), .B(r_x_data[46]), .C(r_add_B[14]), .D(n458), .Y(
        n515) );
  oa21d1_hd U774 ( .A(n516), .B(n454), .C(n515), .Y(n365) );
  ao22d1_hd U775 ( .A(n34), .B(r_x_data[47]), .C(r_add_B[15]), .D(n458), .Y(
        n517) );
  oa21d1_hd U776 ( .A(n518), .B(n454), .C(n517), .Y(n364) );
  ao22d1_hd U777 ( .A(n34), .B(r_x_data[48]), .C(r_add_B[16]), .D(n458), .Y(
        n519) );
  oa21d1_hd U778 ( .A(n520), .B(n454), .C(n519), .Y(n363) );
  ao22d1_hd U779 ( .A(n34), .B(r_x_data[49]), .C(r_add_B[17]), .D(n458), .Y(
        n521) );
  oa21d1_hd U780 ( .A(n522), .B(n454), .C(n521), .Y(n362) );
  ao22d1_hd U781 ( .A(n34), .B(r_x_data[50]), .C(r_add_B[18]), .D(n458), .Y(
        n523) );
  oa21d1_hd U782 ( .A(n524), .B(n454), .C(n523), .Y(n361) );
  ao22d1_hd U783 ( .A(n34), .B(r_x_data[51]), .C(r_add_B[19]), .D(n458), .Y(
        n525) );
  oa21d1_hd U784 ( .A(n526), .B(n454), .C(n525), .Y(n360) );
  ao22d1_hd U785 ( .A(n34), .B(r_x_data[52]), .C(r_add_B[20]), .D(n458), .Y(
        n527) );
  oa21d1_hd U786 ( .A(n528), .B(n454), .C(n527), .Y(n359) );
  ao22d1_hd U787 ( .A(n34), .B(r_x_data[53]), .C(r_add_B[21]), .D(n458), .Y(
        n529) );
  oa21d1_hd U788 ( .A(n530), .B(n454), .C(n529), .Y(n358) );
  ao22d1_hd U789 ( .A(n34), .B(r_x_data[54]), .C(r_add_B[22]), .D(n458), .Y(
        n531) );
  oa21d1_hd U790 ( .A(n532), .B(n454), .C(n531), .Y(n357) );
  ao22d1_hd U791 ( .A(n34), .B(r_x_data[55]), .C(r_add_B[23]), .D(n458), .Y(
        n533) );
  oa21d1_hd U792 ( .A(n534), .B(n454), .C(n533), .Y(n356) );
  ao22d1_hd U793 ( .A(n34), .B(r_x_data[56]), .C(r_add_B[24]), .D(n458), .Y(
        n535) );
  oa21d1_hd U794 ( .A(n536), .B(n454), .C(n535), .Y(n355) );
  ao22d1_hd U795 ( .A(n34), .B(r_x_data[57]), .C(r_add_B[25]), .D(n458), .Y(
        n537) );
  oa21d1_hd U796 ( .A(n538), .B(n454), .C(n537), .Y(n354) );
  ao22d1_hd U797 ( .A(n34), .B(r_x_data[58]), .C(r_add_B[26]), .D(n458), .Y(
        n539) );
  oa21d1_hd U798 ( .A(n540), .B(n454), .C(n539), .Y(n353) );
  ao22d1_hd U799 ( .A(n34), .B(r_x_data[59]), .C(r_add_B[27]), .D(n458), .Y(
        n541) );
  oa21d1_hd U800 ( .A(n542), .B(n454), .C(n541), .Y(n352) );
  ao22d1_hd U801 ( .A(n34), .B(r_x_data[60]), .C(r_add_B[28]), .D(n458), .Y(
        n543) );
  oa21d1_hd U802 ( .A(n544), .B(n454), .C(n543), .Y(n351) );
  ao22d1_hd U803 ( .A(n34), .B(r_x_data[61]), .C(r_add_B[29]), .D(n458), .Y(
        n545) );
  oa21d1_hd U804 ( .A(n546), .B(n454), .C(n545), .Y(n350) );
  ao22d1_hd U805 ( .A(n34), .B(r_x_data[62]), .C(r_add_B[30]), .D(n458), .Y(
        n547) );
  oa21d1_hd U806 ( .A(n549), .B(n454), .C(n547), .Y(n349) );
  ao22d1_hd U807 ( .A(o_Y_DATA[31]), .B(n548), .C(r_add_B[31]), .D(n458), .Y(
        n550) );
  oa21d1_hd U808 ( .A(r_x_data[63]), .B(n452), .C(n550), .Y(n348) );
  ao211d1_hd U809 ( .A(n449), .B(n342), .C(n551), .D(n343), .Y(n212) );
  nr2d1_hd U810 ( .A(n555), .B(n552), .Y(n557) );
  nr2d1_hd U811 ( .A(n554), .B(n553), .Y(n556) );
  ao22d1_hd U812 ( .A(n557), .B(r_counter_0_), .C(n556), .D(n555), .Y(n211) );
  ao22d1_hd U813 ( .A(n223), .B(n557), .C(n556), .D(r_counter_0_), .Y(n210) );
  scg14d1_hd U814 ( .A(r_x_data[31]), .B(n450), .C(n558), .Y(n178) );
  scg14d1_hd U815 ( .A(r_x_data[30]), .B(n450), .C(n559), .Y(n179) );
  scg14d1_hd U816 ( .A(r_x_data[29]), .B(n450), .C(n560), .Y(n180) );
  scg14d1_hd U817 ( .A(r_x_data[28]), .B(n450), .C(n561), .Y(n181) );
  scg14d1_hd U818 ( .A(r_x_data[27]), .B(n450), .C(n562), .Y(n182) );
  scg14d1_hd U819 ( .A(r_x_data[26]), .B(n450), .C(n563), .Y(n183) );
  scg14d1_hd U820 ( .A(r_x_data[25]), .B(n450), .C(n564), .Y(n184) );
  scg14d1_hd U821 ( .A(r_x_data[24]), .B(n450), .C(n565), .Y(n185) );
  scg14d1_hd U822 ( .A(r_x_data[23]), .B(n450), .C(n566), .Y(n186) );
  scg14d1_hd U823 ( .A(r_x_data[22]), .B(n450), .C(n567), .Y(n187) );
  scg14d1_hd U824 ( .A(r_x_data[21]), .B(n450), .C(n568), .Y(n188) );
  scg14d1_hd U825 ( .A(r_x_data[20]), .B(n450), .C(n569), .Y(n189) );
  scg14d1_hd U826 ( .A(r_x_data[19]), .B(n450), .C(n570), .Y(n190) );
  scg14d1_hd U827 ( .A(r_x_data[18]), .B(n450), .C(n571), .Y(n191) );
  scg14d1_hd U828 ( .A(r_x_data[17]), .B(n450), .C(n572), .Y(n192) );
  scg14d1_hd U829 ( .A(r_x_data[16]), .B(n450), .C(n573), .Y(n193) );
  scg14d1_hd U830 ( .A(r_x_data[15]), .B(n450), .C(n574), .Y(n194) );
  scg14d1_hd U831 ( .A(r_x_data[14]), .B(n450), .C(n575), .Y(n195) );
  scg14d1_hd U832 ( .A(r_x_data[13]), .B(n450), .C(n576), .Y(n196) );
  scg14d1_hd U833 ( .A(r_x_data[12]), .B(n450), .C(n577), .Y(n197) );
  scg14d1_hd U834 ( .A(r_x_data[11]), .B(n450), .C(n578), .Y(n198) );
  scg14d1_hd U835 ( .A(r_x_data[10]), .B(n450), .C(n579), .Y(n199) );
  scg14d1_hd U836 ( .A(r_x_data[9]), .B(n450), .C(n580), .Y(n200) );
  scg14d1_hd U837 ( .A(r_x_data[8]), .B(n450), .C(n581), .Y(n201) );
  scg14d1_hd U838 ( .A(r_x_data[7]), .B(n450), .C(n582), .Y(n202) );
  scg14d1_hd U839 ( .A(r_x_data[6]), .B(n450), .C(n583), .Y(n203) );
  scg14d1_hd U840 ( .A(r_x_data[5]), .B(n450), .C(n584), .Y(n204) );
  scg14d1_hd U841 ( .A(r_x_data[4]), .B(n450), .C(n585), .Y(n205) );
  scg14d1_hd U842 ( .A(r_x_data[3]), .B(n450), .C(n586), .Y(n206) );
  scg14d1_hd U843 ( .A(r_x_data[2]), .B(n450), .C(n587), .Y(n207) );
  scg14d1_hd U844 ( .A(r_x_data[1]), .B(n450), .C(n588), .Y(n208) );
  scg14d1_hd U845 ( .A(r_x_data[0]), .B(n450), .C(n589), .Y(n209) );
endmodule

