
module async_rstn_synchronizer ( i_CLK, i_RSTN, o_RSTN );
  input i_CLK, i_RSTN;
  output o_RSTN;
  wire   r_ff;

  fd2qd1_hd:1 o_RSTN_reg ( .D(r_ff), .CK(i_CLK), .RN(i_RSTN), .Q(o_RSTN) );
  fd2qd1_hd:1 r_ff_reg ( .D(1'b1), .CK(i_CLK), .RN(i_RSTN), .Q(r_ff) );
endmodule


module async_rstn_glitch_synchronizer ( i_CLK, i_RSTN, o_RSTN );
  input i_CLK, i_RSTN;
  output o_RSTN;
  wire   w_or_1, eco_net, eco_net_1, eco_net_2, eco_net_3;

  or2d8_hd u__tmp100 ( .A(eco_net), .B(i_RSTN), .Y(w_or_1) );
  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        w_or_1), .o_RSTN(o_RSTN) );
  nid1_hd eco_cell ( .A(eco_net_1), .Y(eco_net) );
  nid1_hd eco_cell_1 ( .A(eco_net_2), .Y(eco_net_1) );
  nid1_hd eco_cell_2 ( .A(eco_net_3), .Y(eco_net_2) );
  nid1_hd eco_cell_3 ( .A(i_RSTN), .Y(eco_net_3) );
endmodule


module divider_by_2 ( i_CLK, i_RSTN, o_CLK_DIV_2 );
  input i_CLK, i_RSTN;
  output o_CLK_DIV_2;


  fj4d1_hd o_CLK_DIV_2_reg ( .J(1'b1), .K(1'b1), .CK(i_CLK), .SN(i_RSTN), .RN(
        1'b1), .Q(o_CLK_DIV_2) );
endmodule


module async_rst_synchronizer ( i_CLK, i_RSTN, o_RST );
  input i_CLK, i_RSTN;
  output o_RST;
  wire   r_ff;

  fd3qd1_hd r_ff_reg ( .D(1'b0), .CK(i_CLK), .SN(i_RSTN), .Q(r_ff) );
  fd3qd1_hd o_RST_reg ( .D(r_ff), .CK(i_CLK), .SN(i_RSTN), .Q(o_RST) );
endmodule


module uart_tx_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  had1_hd U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  had1_hd U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  had1_hd U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  had1_hd U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  had1_hd U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  had1_hd U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  xo2d1_hd U11 ( .A(n1), .B(A[7]), .Y(SUM[7]) );
  ivd1_hd U12 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_uart_tx_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_uart_tx_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module uart_tx ( i_CLK, i_RSTN, i_Tx_DV, i_Tx_Byte, o_Tx_Serial, o_Tx_Done );
  input [7:0] i_Tx_Byte;
  input i_CLK, i_RSTN, i_Tx_DV;
  output o_Tx_Serial, o_Tx_Done;
  wire   w_rst, N21, N22, N23, N24, N25, N26, N29, N32, N35, N42, N44, N45,
         N46, N47, N48, N49, N50, N51, N62, N77, N78, N95, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N130, N131, N132, N134, N135, N141, add_x_3_n1, lt_x_2_n9,
         lt_x_2_n7, lt_x_2_n5, n1, n2, n4, n5, n6, n7, n9, n10, n11, n30, n34,
         n35, n36, n37, n38, n39, n40, n41, n48, n51, n72, n73, n74, n75, n76,
         n77, n78, n79, n80;
  wire   [2:0] r_SM_Main;
  wire   [7:0] r_Clock_Count;
  wire   [2:0] r_Bit_Index;
  wire   [7:0] r_Tx_Data;

  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  had1_hd add_x_3_U2 ( .A(r_Bit_Index[1]), .B(r_Bit_Index[0]), .CO(add_x_3_n1), 
        .S(N77) );
  nr2d1_hd lt_x_2_U9 ( .A(lt_x_2_n9), .B(lt_x_2_n7), .Y(lt_x_2_n5) );
  ao22d1_hd U8 ( .A(N95), .B(n35), .C(n30), .D(N42), .Y(n1) );
  ad2d1_hd U10 ( .A(N25), .B(i_Tx_DV), .Y(N132) );
  nr2bd1_hd U11 ( .AN(N78), .B(n6), .Y(N128) );
  nr2bd1_hd U12 ( .AN(N77), .B(n6), .Y(N127) );
  nr2d1_hd U13 ( .A(r_Bit_Index[0]), .B(n6), .Y(N126) );
  or2d1_hd U14 ( .A(n38), .B(n2), .Y(n6) );
  or2d1_hd U15 ( .A(N25), .B(n4), .Y(N125) );
  nr2d1_hd U16 ( .A(N42), .B(n2), .Y(n4) );
  ad2d1_hd U17 ( .A(N51), .B(n7), .Y(N124) );
  ad2d1_hd U18 ( .A(N50), .B(n7), .Y(N123) );
  ad2d1_hd U19 ( .A(N49), .B(n7), .Y(N122) );
  ad2d1_hd U20 ( .A(N48), .B(n7), .Y(N121) );
  ad2d1_hd U21 ( .A(N47), .B(n7), .Y(N120) );
  ad2d1_hd U22 ( .A(N46), .B(n7), .Y(N119) );
  ad2d1_hd U23 ( .A(N45), .B(n7), .Y(N118) );
  ad2d1_hd U24 ( .A(N44), .B(n7), .Y(N117) );
  oa21d1_hd U25 ( .A(N95), .B(n2), .C(n5), .Y(n7) );
  oa21d1_hd U26 ( .A(n30), .B(n35), .C(N42), .Y(n5) );
  ivd1_hd U27 ( .A(n36), .Y(n2) );
  or2d1_hd U28 ( .A(N131), .B(N141), .Y(N115) );
  nr2bd1_hd U29 ( .AN(n30), .B(N42), .Y(N131) );
  scg6d1_hd U31 ( .A(N62), .B(n36), .C(N135), .Y(N114) );
  or2d1_hd U54 ( .A(N21), .B(r_SM_Main[1]), .Y(N35) );
  ad2d1_hd U55 ( .A(N24), .B(N23), .Y(N25) );
  ad2d1_hd U56 ( .A(N21), .B(N22), .Y(N24) );
  or2d1_hd U57 ( .A(r_SM_Main[2]), .B(r_SM_Main[1]), .Y(N26) );
  or2d1_hd U58 ( .A(r_SM_Main[2]), .B(N22), .Y(N32) );
  or2d1_hd U59 ( .A(r_SM_Main[2]), .B(N22), .Y(N29) );
  or4d1_hd U60 ( .A(N25), .B(n35), .C(n36), .D(n30), .Y(N113) );
  or2d1_hd U78 ( .A(n30), .B(n37), .Y(N116) );
  clknd2d1_hd U79 ( .A(n1), .B(n2), .Y(N130) );
  mx2d1_hd U80 ( .D0(r_Bit_Index[1]), .D1(N127), .S(N125), .Y(n9) );
  mx2d1_hd U81 ( .D0(r_Bit_Index[0]), .D1(N126), .S(N125), .Y(n10) );
  mx2d1_hd U82 ( .D0(o_Tx_Serial), .D1(N114), .S(N134), .Y(n34) );
  ad2d1_hd U83 ( .A(N113), .B(n51), .Y(N134) );
  mx2d1_hd U84 ( .D0(n39), .D1(n40), .S(r_Bit_Index[2]), .Y(N62) );
  mx2d1_hd U85 ( .D0(r_Bit_Index[2]), .D1(N128), .S(N125), .Y(n11) );
  xo2d1_hd U86 ( .A(add_x_3_n1), .B(r_Bit_Index[2]), .Y(N78) );
  nr2d1_hd U88 ( .A(N32), .B(N23), .Y(n30) );
  ivd1_hd U89 ( .A(r_Bit_Index[1]), .Y(lt_x_2_n9) );
  nr2d1_hd U93 ( .A(N26), .B(N23), .Y(n35) );
  ivd1_hd U94 ( .A(N42), .Y(N95) );
  nr2d1_hd U95 ( .A(N29), .B(r_SM_Main[0]), .Y(n36) );
  nr2d1_hd U96 ( .A(N35), .B(r_SM_Main[0]), .Y(n37) );
  or2d1_hd U97 ( .A(N25), .B(n37), .Y(N141) );
  ad2d1_hd U98 ( .A(lt_x_2_n5), .B(r_Bit_Index[0]), .Y(n38) );
  or2d1_hd U99 ( .A(N25), .B(n30), .Y(N135) );
  mx4d1_hd U100 ( .D0(r_Tx_Data[0]), .D1(r_Tx_Data[1]), .D2(r_Tx_Data[2]), 
        .D3(r_Tx_Data[3]), .S0(r_Bit_Index[0]), .S1(r_Bit_Index[1]), .Y(n39)
         );
  mx4d1_hd U101 ( .D0(r_Tx_Data[4]), .D1(r_Tx_Data[5]), .D2(r_Tx_Data[6]), 
        .D3(r_Tx_Data[7]), .S0(r_Bit_Index[0]), .S1(r_Bit_Index[1]), .Y(n40)
         );
  ad2d1_hd U102 ( .A(r_Clock_Count[3]), .B(r_Clock_Count[4]), .Y(n41) );
  oa211d1_hd U103 ( .A(n41), .B(r_Clock_Count[5]), .C(r_Clock_Count[6]), .D(
        r_Clock_Count[7]), .Y(N42) );
  ivd1_hd U36 ( .A(w_rst), .Y(n48) );
  ivd1_hd U39 ( .A(w_rst), .Y(n51) );
  uart_tx_DW01_inc_0 add_x_1 ( .A(r_Clock_Count), .SUM({N51, N50, N49, N48, 
        N47, N46, N45, N44}) );
  SNPS_CLOCK_GATE_HIGH_uart_tx_4 clk_gate_r_Clock_Count_reg_6__0 ( .CLK(i_CLK), 
        .EN(N113), .ENCLK(n73), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_uart_tx_5 clk_gate_r_Tx_Data_reg_7__0 ( .CLK(i_CLK), 
        .EN(N132), .ENCLK(n72), .TE(1'b0) );
  fd2qd1_hd r_Bit_Index_reg_1_ ( .D(n9), .CK(n73), .RN(n51), .Q(r_Bit_Index[1]) );
  fd2qd1_hd r_Bit_Index_reg_0_ ( .D(n10), .CK(n73), .RN(n51), .Q(
        r_Bit_Index[0]) );
  fd1qd1_hd o_Tx_Serial_reg ( .D(n34), .CK(n73), .Q(o_Tx_Serial) );
  fd2qd1_hd r_SM_Main_reg_2_ ( .D(N131), .CK(i_CLK), .RN(n48), .Q(r_SM_Main[2]) );
  fd2qd1_hd r_SM_Main_reg_1_ ( .D(N130), .CK(i_CLK), .RN(n48), .Q(r_SM_Main[1]) );
  fd2qd1_hd r_Tx_Done_reg ( .D(n74), .CK(i_CLK), .RN(n51), .Q(o_Tx_Done) );
  fd2qd1_hd r_Bit_Index_reg_2_ ( .D(n11), .CK(n73), .RN(n51), .Q(
        r_Bit_Index[2]) );
  fd2qd1_hd r_Clock_Count_reg_7_ ( .D(N124), .CK(n73), .RN(n48), .Q(
        r_Clock_Count[7]) );
  fd2qd1_hd r_Clock_Count_reg_6_ ( .D(N123), .CK(n73), .RN(n51), .Q(
        r_Clock_Count[6]) );
  fd2qd1_hd r_Clock_Count_reg_5_ ( .D(N122), .CK(n73), .RN(n48), .Q(
        r_Clock_Count[5]) );
  fd2qd1_hd r_Clock_Count_reg_4_ ( .D(N121), .CK(n73), .RN(n51), .Q(
        r_Clock_Count[4]) );
  fd2qd1_hd r_Clock_Count_reg_3_ ( .D(N120), .CK(n73), .RN(n48), .Q(
        r_Clock_Count[3]) );
  fd2qd1_hd r_Clock_Count_reg_2_ ( .D(N119), .CK(n73), .RN(n48), .Q(
        r_Clock_Count[2]) );
  fd2qd1_hd r_Clock_Count_reg_1_ ( .D(N118), .CK(n73), .RN(n48), .Q(
        r_Clock_Count[1]) );
  fd2qd1_hd r_Clock_Count_reg_0_ ( .D(N117), .CK(n73), .RN(n51), .Q(
        r_Clock_Count[0]) );
  fd2qd1_hd r_Tx_Data_reg_7_ ( .D(i_Tx_Byte[7]), .CK(n72), .RN(n48), .Q(
        r_Tx_Data[7]) );
  fd2qd1_hd r_Tx_Data_reg_6_ ( .D(i_Tx_Byte[6]), .CK(n72), .RN(n48), .Q(
        r_Tx_Data[6]) );
  fd2qd1_hd r_Tx_Data_reg_5_ ( .D(i_Tx_Byte[5]), .CK(n72), .RN(n48), .Q(
        r_Tx_Data[5]) );
  fd2qd1_hd r_Tx_Data_reg_4_ ( .D(i_Tx_Byte[4]), .CK(n72), .RN(n48), .Q(
        r_Tx_Data[4]) );
  fd2qd1_hd r_Tx_Data_reg_3_ ( .D(i_Tx_Byte[3]), .CK(n72), .RN(n48), .Q(
        r_Tx_Data[3]) );
  fd2qd1_hd r_Tx_Data_reg_2_ ( .D(i_Tx_Byte[2]), .CK(n72), .RN(n51), .Q(
        r_Tx_Data[2]) );
  fd2qd1_hd r_Tx_Data_reg_1_ ( .D(i_Tx_Byte[1]), .CK(n72), .RN(n51), .Q(
        r_Tx_Data[1]) );
  fd2qd1_hd r_Tx_Data_reg_0_ ( .D(i_Tx_Byte[0]), .CK(n72), .RN(n51), .Q(
        r_Tx_Data[0]) );
  fd2qd1_hd r_SM_Main_reg_0_ ( .D(n75), .CK(i_CLK), .RN(n51), .Q(r_SM_Main[0])
         );
  ivd1_hd U1 ( .A(r_SM_Main[2]), .Y(N21) );
  ivd1_hd U2 ( .A(r_SM_Main[0]), .Y(N23) );
  ivd1_hd U3 ( .A(r_Bit_Index[2]), .Y(lt_x_2_n7) );
  mx2d1_hd U4 ( .D0(r_SM_Main[0]), .D1(n79), .S(n80), .Y(n75) );
  mx2d1_hd U5 ( .D0(o_Tx_Done), .D1(N116), .S(N115), .Y(n74) );
  ivd1_hd U6 ( .A(r_SM_Main[1]), .Y(N22) );
  ao211d1_hd U7 ( .A(r_SM_Main[1]), .B(n76), .C(r_SM_Main[2]), .D(n77), .Y(n79) );
  ao21d1_hd U9 ( .A(n78), .B(i_Tx_DV), .C(r_SM_Main[1]), .Y(n77) );
  nd2bd1_hd U30 ( .AN(N42), .B(r_SM_Main[0]), .Y(n78) );
  scg13d1_hd U32 ( .A(r_SM_Main[0]), .B(N42), .C(n38), .Y(n76) );
  scg17d1_hd U33 ( .A(i_Tx_DV), .B(N22), .C(r_SM_Main[2]), .D(N42), .Y(n80) );
endmodule


module uart_rx_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  had1_hd U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  had1_hd U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  had1_hd U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  had1_hd U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  had1_hd U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  had1_hd U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  xo2d1_hd U11 ( .A(n1), .B(A[7]), .Y(SUM[7]) );
  ivd1_hd U12 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_uart_rx_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module uart_rx ( i_CLK, i_RSTN, i_Rx_Serial, o_Rx_DV, o_Rx_Byte );
  output [7:0] o_Rx_Byte;
  input i_CLK, i_RSTN, i_Rx_Serial;
  output o_Rx_DV;
  wire   w_rst, r_Rx_Data, r_Rx_Data_R, N31, N32, N33, N34, N35, N36, N39, N42,
         N45, N52, N53, N54, N55, N56, N57, N58, N59, N71, N72, N85, N86, N129,
         N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140,
         N141, N142, N143, N144, N146, N147, N148, N149, N150, N151, N152,
         N153, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N169, N172, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, add_x_3_n1, lt_x_2_n13,
         lt_x_2_n9, lt_x_2_n7, lt_x_2_n5, n2, n4, n5, n6, n7, n8, n9, n11, n12,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n31, n33, n36, n37,
         n38, n39, n40, n41, n42, n43, n52, n55, n77, n78;
  wire   [2:0] r_SM_Main;
  wire   [7:0] r_Clock_Count;
  wire   [2:0] r_Bit_Index;

  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  had1_hd add_x_3_U2 ( .A(r_Bit_Index[1]), .B(r_Bit_Index[0]), .CO(add_x_3_n1), 
        .S(N85) );
  nr2d1_hd lt_x_2_U9 ( .A(lt_x_2_n9), .B(lt_x_2_n7), .Y(lt_x_2_n5) );
  ad2d1_hd U8 ( .A(N176), .B(n2), .Y(N153) );
  ad2d1_hd U9 ( .A(N178), .B(n2), .Y(N152) );
  ad2d1_hd U10 ( .A(N180), .B(n2), .Y(N151) );
  ad2d1_hd U11 ( .A(N182), .B(n2), .Y(N150) );
  ad2d1_hd U12 ( .A(N184), .B(n2), .Y(N149) );
  ad2d1_hd U13 ( .A(N186), .B(n2), .Y(N148) );
  ad2d1_hd U14 ( .A(N188), .B(n2), .Y(N147) );
  ad2d1_hd U15 ( .A(N190), .B(n2), .Y(N146) );
  oa211d1_hd U16 ( .A(n39), .B(n4), .C(n5), .D(n6), .Y(N144) );
  scg7d1_hd U18 ( .A(n2), .B(n42), .C(N35), .D(n7), .E(n8), .Y(N143) );
  nr2bd1_hd U19 ( .AN(N86), .B(n9), .Y(N142) );
  nr2bd1_hd U20 ( .AN(N85), .B(n9), .Y(N141) );
  nr2d1_hd U21 ( .A(r_Bit_Index[0]), .B(n9), .Y(N140) );
  or2d1_hd U22 ( .A(n42), .B(n6), .Y(n9) );
  or2d1_hd U23 ( .A(n2), .B(N35), .Y(N139) );
  nr2d1_hd U24 ( .A(N71), .B(n6), .Y(n2) );
  ivd1_hd U25 ( .A(n40), .Y(n6) );
  nr2bd1_hd U26 ( .AN(N59), .B(n11), .Y(N138) );
  nr2bd1_hd U27 ( .AN(N58), .B(n11), .Y(N137) );
  nr2bd1_hd U28 ( .AN(N57), .B(n11), .Y(N136) );
  nr2bd1_hd U29 ( .AN(N56), .B(n11), .Y(N135) );
  nr2bd1_hd U30 ( .AN(N55), .B(n11), .Y(N134) );
  nr2bd1_hd U31 ( .AN(N54), .B(n11), .Y(N133) );
  nr2bd1_hd U32 ( .AN(N53), .B(n11), .Y(N132) );
  nr2bd1_hd U33 ( .AN(N52), .B(n11), .Y(N131) );
  ao21d1_hd U34 ( .A(n40), .B(N71), .C(n8), .Y(n11) );
  scg17d1_hd U38 ( .A(n37), .B(n7), .C(N172), .D(n12), .Y(N130) );
  or2d1_hd U41 ( .A(N169), .B(n38), .Y(N129) );
  or2d1_hd U66 ( .A(r_Clock_Count[4]), .B(N160), .Y(N161) );
  or2d1_hd U67 ( .A(N156), .B(N159), .Y(N160) );
  or2d1_hd U68 ( .A(N155), .B(r_Clock_Count[7]), .Y(N159) );
  ivd1_hd U69 ( .A(r_SM_Main[2]), .Y(N31) );
  ivd1_hd U70 ( .A(r_SM_Main[1]), .Y(N32) );
  clknd2d1_hd U71 ( .A(n37), .B(n39), .Y(n12) );
  or2d1_hd U72 ( .A(r_SM_Main[2]), .B(N32), .Y(N39) );
  clknd2d1_hd U73 ( .A(n5), .B(n12), .Y(n8) );
  or2d1_hd U74 ( .A(r_Clock_Count[1]), .B(N163), .Y(N164) );
  or2d1_hd U75 ( .A(N158), .B(N162), .Y(N163) );
  or2d1_hd U76 ( .A(N157), .B(N161), .Y(N162) );
  clknd2d1_hd U77 ( .A(n36), .B(N71), .Y(n5) );
  or2d1_hd U78 ( .A(r_SM_Main[2]), .B(r_SM_Main[1]), .Y(N36) );
  or2d1_hd U79 ( .A(N31), .B(r_SM_Main[1]), .Y(N45) );
  ad2d1_hd U80 ( .A(N34), .B(N33), .Y(N35) );
  ad2d1_hd U81 ( .A(N31), .B(N32), .Y(N34) );
  or2d1_hd U82 ( .A(r_SM_Main[2]), .B(N32), .Y(N42) );
  mx2d1_hd U83 ( .D0(r_Clock_Count[0]), .D1(N131), .S(N130), .Y(n31) );
  mx2d1_hd U87 ( .D0(o_Rx_Byte[0]), .D1(r_Rx_Data), .S(N146), .Y(n15) );
  ad2d1_hd U88 ( .A(N189), .B(lt_x_2_n7), .Y(N190) );
  ad2d1_hd U89 ( .A(lt_x_2_n13), .B(lt_x_2_n9), .Y(N189) );
  mx2d1_hd U90 ( .D0(o_Rx_Byte[1]), .D1(r_Rx_Data), .S(N147), .Y(n16) );
  ad2d1_hd U91 ( .A(N187), .B(lt_x_2_n7), .Y(N188) );
  ad2d1_hd U92 ( .A(r_Bit_Index[0]), .B(lt_x_2_n9), .Y(N187) );
  mx2d1_hd U93 ( .D0(o_Rx_Byte[2]), .D1(r_Rx_Data), .S(N148), .Y(n17) );
  ad2d1_hd U94 ( .A(N185), .B(lt_x_2_n7), .Y(N186) );
  ad2d1_hd U95 ( .A(lt_x_2_n13), .B(r_Bit_Index[1]), .Y(N185) );
  mx2d1_hd U96 ( .D0(o_Rx_Byte[3]), .D1(r_Rx_Data), .S(N149), .Y(n18) );
  ad2d1_hd U97 ( .A(N183), .B(lt_x_2_n7), .Y(N184) );
  ad2d1_hd U98 ( .A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Y(N183) );
  mx2d1_hd U99 ( .D0(o_Rx_Byte[4]), .D1(r_Rx_Data), .S(N150), .Y(n19) );
  ad2d1_hd U100 ( .A(N181), .B(r_Bit_Index[2]), .Y(N182) );
  ad2d1_hd U101 ( .A(lt_x_2_n13), .B(lt_x_2_n9), .Y(N181) );
  mx2d1_hd U102 ( .D0(o_Rx_Byte[5]), .D1(r_Rx_Data), .S(N151), .Y(n20) );
  ad2d1_hd U103 ( .A(N179), .B(r_Bit_Index[2]), .Y(N180) );
  ad2d1_hd U104 ( .A(r_Bit_Index[0]), .B(lt_x_2_n9), .Y(N179) );
  mx2d1_hd U105 ( .D0(o_Rx_Byte[6]), .D1(r_Rx_Data), .S(N152), .Y(n21) );
  ad2d1_hd U106 ( .A(N177), .B(r_Bit_Index[2]), .Y(N178) );
  ad2d1_hd U107 ( .A(lt_x_2_n13), .B(r_Bit_Index[1]), .Y(N177) );
  mx2d1_hd U108 ( .D0(o_Rx_Byte[7]), .D1(r_Rx_Data), .S(N153), .Y(n22) );
  ad2d1_hd U109 ( .A(N175), .B(r_Bit_Index[2]), .Y(N176) );
  ad2d1_hd U110 ( .A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Y(N175) );
  clknd2d1_hd U111 ( .A(n37), .B(n7), .Y(n4) );
  mx2d1_hd U113 ( .D0(r_Bit_Index[2]), .D1(N142), .S(N139), .Y(n23) );
  xo2d1_hd U114 ( .A(add_x_3_n1), .B(r_Bit_Index[2]), .Y(N86) );
  mx2d1_hd U115 ( .D0(r_Bit_Index[1]), .D1(N141), .S(N139), .Y(n24) );
  mx2d1_hd U116 ( .D0(r_Bit_Index[0]), .D1(N140), .S(N139), .Y(n33) );
  ivd1_hd U122 ( .A(r_SM_Main[0]), .Y(N33) );
  ivd1_hd U123 ( .A(r_Rx_Data), .Y(n7) );
  ivd1_hd U124 ( .A(N71), .Y(N72) );
  nr2d1_hd U125 ( .A(N42), .B(N33), .Y(n36) );
  nr2d1_hd U126 ( .A(N36), .B(N33), .Y(n37) );
  ad2d1_hd U127 ( .A(N72), .B(n36), .Y(n38) );
  or2d1_hd U128 ( .A(r_Clock_Count[0]), .B(N164), .Y(n39) );
  nr2d1_hd U129 ( .A(N39), .B(r_SM_Main[0]), .Y(n40) );
  or3d1_hd U130 ( .A(N35), .B(n40), .C(n36), .Y(N172) );
  nr2d1_hd U131 ( .A(N45), .B(r_SM_Main[0]), .Y(n41) );
  or2d1_hd U132 ( .A(N35), .B(n41), .Y(N169) );
  ad2d1_hd U133 ( .A(lt_x_2_n5), .B(r_Bit_Index[0]), .Y(n42) );
  ad2d1_hd U134 ( .A(r_Clock_Count[3]), .B(r_Clock_Count[4]), .Y(n43) );
  oa211d1_hd U135 ( .A(n43), .B(r_Clock_Count[5]), .C(r_Clock_Count[6]), .D(
        r_Clock_Count[7]), .Y(N71) );
  fd3qd1_hd r_Rx_Data_reg ( .D(r_Rx_Data_R), .CK(i_CLK), .SN(n52), .Q(
        r_Rx_Data) );
  fd3qd1_hd r_Rx_Data_R_reg ( .D(i_Rx_Serial), .CK(i_CLK), .SN(n52), .Q(
        r_Rx_Data_R) );
  ivd1_hd U42 ( .A(w_rst), .Y(n52) );
  ivd1_hd U45 ( .A(w_rst), .Y(n55) );
  uart_rx_DW01_inc_0 add_x_1 ( .A(r_Clock_Count), .SUM({N59, N58, N57, N56, 
        N55, N54, N53, N52}) );
  SNPS_CLOCK_GATE_HIGH_uart_rx_2 clk_gate_r_Clock_Count_reg_7__0 ( .CLK(i_CLK), 
        .EN(N130), .ENCLK(n77), .TE(1'b0) );
  fd2qd1_hd r_SM_Main_reg_2_ ( .D(n38), .CK(i_CLK), .RN(n52), .Q(r_SM_Main[2])
         );
  fd2qd1_hd r_Rx_DV_reg ( .D(n78), .CK(i_CLK), .RN(n52), .Q(o_Rx_DV) );
  fd2qd1_hd r_SM_Main_reg_1_ ( .D(N144), .CK(i_CLK), .RN(n55), .Q(r_SM_Main[1]) );
  fd2qd1_hd r_Rx_Byte_reg_7_ ( .D(n22), .CK(n77), .RN(n52), .Q(o_Rx_Byte[7])
         );
  fd2qd1_hd r_Rx_Byte_reg_6_ ( .D(n21), .CK(n77), .RN(n52), .Q(o_Rx_Byte[6])
         );
  fd2qd1_hd r_Rx_Byte_reg_5_ ( .D(n20), .CK(n77), .RN(n55), .Q(o_Rx_Byte[5])
         );
  fd2qd1_hd r_Rx_Byte_reg_4_ ( .D(n19), .CK(n77), .RN(n55), .Q(o_Rx_Byte[4])
         );
  fd2qd1_hd r_Rx_Byte_reg_3_ ( .D(n18), .CK(n77), .RN(n55), .Q(o_Rx_Byte[3])
         );
  fd2qd1_hd r_Rx_Byte_reg_2_ ( .D(n17), .CK(n77), .RN(n52), .Q(o_Rx_Byte[2])
         );
  fd2qd1_hd r_Rx_Byte_reg_1_ ( .D(n16), .CK(n77), .RN(n55), .Q(o_Rx_Byte[1])
         );
  fd2qd1_hd r_Rx_Byte_reg_0_ ( .D(n15), .CK(n77), .RN(n55), .Q(o_Rx_Byte[0])
         );
  fd2qd1_hd r_Bit_Index_reg_2_ ( .D(n23), .CK(n77), .RN(n55), .Q(
        r_Bit_Index[2]) );
  fd2qd1_hd r_Bit_Index_reg_1_ ( .D(n24), .CK(n77), .RN(n55), .Q(
        r_Bit_Index[1]) );
  fd2qd1_hd r_Bit_Index_reg_0_ ( .D(n33), .CK(n77), .RN(n52), .Q(
        r_Bit_Index[0]) );
  fd2qd1_hd r_SM_Main_reg_0_ ( .D(N143), .CK(i_CLK), .RN(n55), .Q(r_SM_Main[0]) );
  fd2qd1_hd r_Clock_Count_reg_7_ ( .D(N138), .CK(n77), .RN(n55), .Q(
        r_Clock_Count[7]) );
  fd2qd1_hd r_Clock_Count_reg_6_ ( .D(N137), .CK(n77), .RN(n52), .Q(
        r_Clock_Count[6]) );
  fd2qd1_hd r_Clock_Count_reg_5_ ( .D(N136), .CK(n77), .RN(n55), .Q(
        r_Clock_Count[5]) );
  fd2qd1_hd r_Clock_Count_reg_4_ ( .D(N135), .CK(n77), .RN(n52), .Q(
        r_Clock_Count[4]) );
  fd2qd1_hd r_Clock_Count_reg_3_ ( .D(N134), .CK(n77), .RN(n55), .Q(
        r_Clock_Count[3]) );
  fd2qd1_hd r_Clock_Count_reg_2_ ( .D(N133), .CK(n77), .RN(n55), .Q(
        r_Clock_Count[2]) );
  fd2qd1_hd r_Clock_Count_reg_1_ ( .D(N132), .CK(n77), .RN(n52), .Q(
        r_Clock_Count[1]) );
  fd2qd1_hd r_Clock_Count_reg_0_ ( .D(n31), .CK(i_CLK), .RN(n52), .Q(
        r_Clock_Count[0]) );
  ivd1_hd U1 ( .A(r_Clock_Count[6]), .Y(N155) );
  ivd1_hd U2 ( .A(r_Clock_Count[5]), .Y(N156) );
  ivd1_hd U3 ( .A(r_Clock_Count[3]), .Y(N157) );
  ivd1_hd U4 ( .A(r_Bit_Index[2]), .Y(lt_x_2_n7) );
  ivd1_hd U5 ( .A(r_Bit_Index[1]), .Y(lt_x_2_n9) );
  ivd1_hd U6 ( .A(r_Bit_Index[0]), .Y(lt_x_2_n13) );
  ivd1_hd U7 ( .A(r_Clock_Count[2]), .Y(N158) );
  mx2d1_hd U17 ( .D0(o_Rx_DV), .D1(n36), .S(N129), .Y(n78) );
endmodule


module SNPS_CLOCK_GATE_HIGH_uart_controller_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_uart_controller_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_uart_controller_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_uart_controller_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module uart_controller ( i_UART_DATA_TX, i_UART_DATA_TX_VALID, 
        o_UART_DATA_TX_READY, o_UART_DATA_RX, o_UART_DATA_RX_VALID, 
        i_CORE_BUSY, i_UART_RXD, o_UART_TXD, i_CLK, i_RSTN );
  input [55:0] i_UART_DATA_TX;
  output [15:0] o_UART_DATA_RX;
  input i_UART_DATA_TX_VALID, i_CORE_BUSY, i_UART_RXD, i_CLK, i_RSTN;
  output o_UART_DATA_TX_READY, o_UART_DATA_RX_VALID, o_UART_TXD;
  wire   w_rst, w_rstn, r_uart_data_tx_valid, w_uart_data_tx_done,
         w_uart_data_rx_valid, N34, N35, N36, N37, N38, N39, N42, N47, N50,
         N51, N54, N60, N62, N120, N121, N122, N127, N128, N129, N130, N131,
         N132, N133, N134, N194, N199, N200, N214, N215, N223, N225, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N305, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N321, N322, N325, N326,
         N327, N328, N329, N330, N333, N334, N335, N336, N337, N338, N339,
         N340, N343, N344, N345, N346, N347, N348, N349, N350, N351, N354,
         N355, N356, N357, N358, N359, N360, N361, N364, N365, N366, N367,
         N368, N369, N370, N371, N372, N375, N376, N377, N378, N379, N380,
         N386, N396, N397, alt45_n18, alt45_n61, alt45_n63, gt_x_3_n7,
         gt_x_3_n5, add_x_2_n1, gt_x_1_n9, gt_x_1_n7, gt_x_1_n5, n1, n5, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n23,
         n109, n110, n111, n112, n113, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331;
  wire   [7:0] r_uart_data_tx;
  wire   [2:0] r_pstate;
  wire   [55:0] r_uart_data_tx_shift;
  wire   [1:0] r_data_counter;
  wire   [1:0] r_lstate;

  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  uart_tx uart_tx ( .i_CLK(i_CLK), .i_RSTN(w_rstn), .i_Tx_DV(
        r_uart_data_tx_valid), .i_Tx_Byte(r_uart_data_tx), .o_Tx_Serial(
        o_UART_TXD), .o_Tx_Done(w_uart_data_tx_done) );
  uart_rx uart_rx ( .i_CLK(i_CLK), .i_RSTN(w_rstn), .i_Rx_Serial(i_UART_RXD), 
        .o_Rx_DV(w_uart_data_rx_valid), .o_Rx_Byte({N134, N133, N132, N131, 
        N130, N129, N128, N127}) );
  nr2d1_hd gt_x_3_U9 ( .A(gt_x_1_n9), .B(gt_x_3_n7), .Y(gt_x_3_n5) );
  had1_hd add_x_2_U2 ( .A(r_data_counter[1]), .B(r_data_counter[0]), .CO(
        add_x_2_n1), .S(N199) );
  nr2d1_hd gt_x_1_U9 ( .A(gt_x_1_n9), .B(gt_x_1_n7), .Y(gt_x_1_n5) );
  nr3d1_hd U5 ( .A(n117), .B(n120), .C(n125), .Y(n1) );
  nr3d1_hd U8 ( .A(r_pstate[1]), .B(r_pstate[0]), .C(N34), .Y(N50) );
  scg12d1_hd U10 ( .A(r_pstate[1]), .B(r_pstate[0]), .C(r_pstate[2]), .Y(N47)
         );
  scg15d1_hd U14 ( .A(n120), .B(n130), .C(n8), .D(n9), .Y(N302) );
  nd2bd1_hd U15 ( .AN(n10), .B(n11), .Y(N301) );
  scg18d1_hd U16 ( .A(n12), .B(N121), .C(n13), .D(n8), .E(n11), .Y(N300) );
  ao22d1_hd U17 ( .A(N194), .B(n120), .C(n14), .D(n15), .Y(n11) );
  ivd1_hd U18 ( .A(N321), .Y(n15) );
  scg17d1_hd U20 ( .A(n14), .B(n131), .C(N397), .D(n9), .Y(N299) );
  scg16d1_hd U21 ( .A(n16), .B(N215), .C(n122), .Y(n9) );
  ad2d1_hd U23 ( .A(n122), .B(w_uart_data_tx_done), .Y(n14) );
  scg14d1_hd U24 ( .A(n12), .B(N122), .C(n17), .Y(N298) );
  ivd1_hd U25 ( .A(n18), .Y(N297) );
  nr2bd1_hd U26 ( .AN(N200), .B(n8), .Y(N296) );
  nr2bd1_hd U27 ( .AN(N199), .B(n8), .Y(N295) );
  nr2d1_hd U28 ( .A(n8), .B(r_data_counter[0]), .Y(N294) );
  ad2d1_hd U77 ( .A(i_UART_DATA_TX[7]), .B(n10), .Y(N244) );
  ad2d1_hd U78 ( .A(i_UART_DATA_TX[6]), .B(n10), .Y(N243) );
  ad2d1_hd U79 ( .A(i_UART_DATA_TX[5]), .B(n10), .Y(N242) );
  ad2d1_hd U80 ( .A(i_UART_DATA_TX[4]), .B(n10), .Y(N241) );
  ad2d1_hd U81 ( .A(i_UART_DATA_TX[3]), .B(n10), .Y(N240) );
  ad2d1_hd U82 ( .A(i_UART_DATA_TX[2]), .B(n10), .Y(N239) );
  ad2d1_hd U83 ( .A(i_UART_DATA_TX[1]), .B(n10), .Y(N238) );
  ad2d1_hd U84 ( .A(i_UART_DATA_TX[0]), .B(n10), .Y(N237) );
  ao21d1_hd U86 ( .A(N60), .B(i_CORE_BUSY), .C(N307), .Y(n20) );
  ad2d1_hd U88 ( .A(r_uart_data_tx_shift[55]), .B(n125), .Y(N235) );
  ad2d1_hd U89 ( .A(r_uart_data_tx_shift[54]), .B(n125), .Y(N234) );
  ad2d1_hd U90 ( .A(r_uart_data_tx_shift[53]), .B(n125), .Y(N233) );
  ad2d1_hd U91 ( .A(r_uart_data_tx_shift[52]), .B(n125), .Y(N232) );
  ad2d1_hd U92 ( .A(r_uart_data_tx_shift[51]), .B(n125), .Y(N231) );
  ad2d1_hd U93 ( .A(r_uart_data_tx_shift[50]), .B(n125), .Y(N230) );
  ad2d1_hd U94 ( .A(r_uart_data_tx_shift[49]), .B(n125), .Y(N229) );
  ad2d1_hd U95 ( .A(r_uart_data_tx_shift[48]), .B(n125), .Y(N228) );
  scg17d1_hd U96 ( .A(n122), .B(N215), .C(N38), .D(n8), .Y(N227) );
  ao22d1_hd U97 ( .A(N214), .B(N50), .C(N47), .D(n21), .Y(n8) );
  ivd1_hd U98 ( .A(n116), .Y(n21) );
  nd4d1_hd U100 ( .A(N38), .B(i_CORE_BUSY), .C(n128), .D(w_uart_data_rx_valid), 
        .Y(n17) );
  nr2bd1_hd U101 ( .AN(N305), .B(n19), .Y(n12) );
  ivd1_hd U107 ( .A(N38), .Y(n19) );
  ao22d1_hd U108 ( .A(N47), .B(n116), .C(N50), .D(n118), .Y(n23) );
  ivd1_hd U202 ( .A(N132), .Y(N364) );
  ivd1_hd U203 ( .A(r_uart_data_tx_shift[54]), .Y(N308) );
  ivd1_hd U204 ( .A(N133), .Y(N343) );
  ivd1_hd U205 ( .A(N134), .Y(N354) );
  ivd1_hd U206 ( .A(N131), .Y(N344) );
  or2d1_hd U207 ( .A(N131), .B(N368), .Y(N369) );
  or2d1_hd U208 ( .A(N364), .B(N367), .Y(N368) );
  or2d1_hd U209 ( .A(N343), .B(N134), .Y(N367) );
  or2d1_hd U210 ( .A(N364), .B(N375), .Y(N376) );
  or2d1_hd U211 ( .A(N343), .B(N134), .Y(N375) );
  ivd1_hd U212 ( .A(i_CORE_BUSY), .Y(alt45_n63) );
  or2d1_hd U213 ( .A(N309), .B(N325), .Y(N326) );
  or2d1_hd U214 ( .A(N308), .B(r_uart_data_tx_shift[55]), .Y(N325) );
  or2d1_hd U215 ( .A(N310), .B(N315), .Y(N316) );
  or2d1_hd U216 ( .A(r_uart_data_tx_shift[52]), .B(N314), .Y(N315) );
  or2d1_hd U217 ( .A(N309), .B(N313), .Y(N314) );
  or2d1_hd U218 ( .A(N308), .B(r_uart_data_tx_shift[55]), .Y(N313) );
  ad2d1_hd U219 ( .A(alt45_n63), .B(N62), .Y(alt45_n61) );
  or2d1_hd U220 ( .A(N344), .B(N347), .Y(N348) );
  or2d1_hd U221 ( .A(N132), .B(N346), .Y(N347) );
  or2d1_hd U222 ( .A(N343), .B(N134), .Y(N346) );
  or2d1_hd U223 ( .A(N130), .B(N358), .Y(N359) );
  or2d1_hd U224 ( .A(N344), .B(N357), .Y(N358) );
  or2d1_hd U225 ( .A(N132), .B(N356), .Y(N357) );
  or2d1_hd U226 ( .A(N133), .B(N354), .Y(N356) );
  ivd1_hd U227 ( .A(N128), .Y(N345) );
  ivd1_hd U228 ( .A(r_pstate[1]), .Y(N35) );
  or2d1_hd U229 ( .A(r_uart_data_tx_shift[54]), .B(N333), .Y(N335) );
  ivd1_hd U230 ( .A(r_uart_data_tx_shift[55]), .Y(N333) );
  ivd1_hd U231 ( .A(r_uart_data_tx_shift[53]), .Y(N309) );
  ivd1_hd U232 ( .A(r_uart_data_tx_shift[51]), .Y(N310) );
  or2d1_hd U233 ( .A(N366), .B(N370), .Y(N371) );
  ivd1_hd U234 ( .A(N129), .Y(N366) );
  or2d1_hd U235 ( .A(N365), .B(N369), .Y(N370) );
  ivd1_hd U236 ( .A(N130), .Y(N365) );
  or2d1_hd U237 ( .A(N128), .B(N379), .Y(N380) );
  or2d1_hd U238 ( .A(N129), .B(N378), .Y(N379) );
  or2d1_hd U239 ( .A(N130), .B(N377), .Y(N378) );
  or2d1_hd U240 ( .A(N131), .B(N376), .Y(N377) );
  ivd1_hd U241 ( .A(N127), .Y(N355) );
  or2d1_hd U242 ( .A(r_uart_data_tx_shift[49]), .B(N329), .Y(N330) );
  or2d1_hd U243 ( .A(r_uart_data_tx_shift[50]), .B(N328), .Y(N329) );
  or2d1_hd U244 ( .A(r_uart_data_tx_shift[51]), .B(N327), .Y(N328) );
  or2d1_hd U245 ( .A(r_uart_data_tx_shift[52]), .B(N326), .Y(N327) );
  ivd1_hd U246 ( .A(r_uart_data_tx_shift[48]), .Y(N312) );
  or2d1_hd U247 ( .A(r_uart_data_tx_shift[49]), .B(N317), .Y(N318) );
  or2d1_hd U248 ( .A(N311), .B(N316), .Y(N317) );
  ivd1_hd U249 ( .A(r_uart_data_tx_shift[50]), .Y(N311) );
  ad2d1_hd U250 ( .A(r_lstate[0]), .B(r_lstate[1]), .Y(N321) );
  clknd2d1_hd U251 ( .A(n19), .B(n1), .Y(N396) );
  ad2d1_hd U252 ( .A(r_pstate[2]), .B(r_pstate[1]), .Y(N54) );
  ad2d1_hd U255 ( .A(i_UART_DATA_TX_VALID), .B(N62), .Y(N60) );
  ad2d1_hd U256 ( .A(i_UART_DATA_TX_VALID), .B(alt45_n61), .Y(N307) );
  or2d1_hd U257 ( .A(n126), .B(N121), .Y(N122) );
  or2d1_hd U258 ( .A(N345), .B(N350), .Y(N351) );
  or2d1_hd U259 ( .A(N129), .B(N349), .Y(N350) );
  or2d1_hd U260 ( .A(N130), .B(N348), .Y(N349) );
  or2d1_hd U261 ( .A(N345), .B(N360), .Y(N361) );
  or2d1_hd U262 ( .A(N129), .B(N359), .Y(N360) );
  ad2d1_hd U263 ( .A(N37), .B(N36), .Y(N38) );
  ad2d1_hd U264 ( .A(N34), .B(N35), .Y(N37) );
  or2d1_hd U265 ( .A(r_pstate[2]), .B(N35), .Y(N42) );
  or2d1_hd U266 ( .A(r_uart_data_tx_shift[50]), .B(N338), .Y(N339) );
  or2d1_hd U267 ( .A(N310), .B(N337), .Y(N338) );
  or2d1_hd U268 ( .A(r_uart_data_tx_shift[52]), .B(N336), .Y(N337) );
  or2d1_hd U269 ( .A(N309), .B(N335), .Y(N336) );
  ivd1_hd U270 ( .A(r_uart_data_tx_shift[49]), .Y(N334) );
  clknd2d1_hd U271 ( .A(N321), .B(w_uart_data_tx_done), .Y(n16) );
  or3d1_hd U272 ( .A(N38), .B(N47), .C(N50), .Y(N293) );
  or2d1_hd U273 ( .A(n127), .B(n119), .Y(N121) );
  or2d1_hd U274 ( .A(N128), .B(N371), .Y(N372) );
  or2d1_hd U275 ( .A(r_pstate[2]), .B(r_pstate[1]), .Y(N39) );
  or2d1_hd U277 ( .A(N34), .B(r_pstate[1]), .Y(N51) );
  or2d1_hd U278 ( .A(n129), .B(n121), .Y(N194) );
  or2d1_hd U279 ( .A(N396), .B(N54), .Y(N397) );
  ivd1_hd U280 ( .A(r_lstate[1]), .Y(N322) );
  mx2d1_hd U385 ( .D0(r_pstate[1]), .D1(N301), .S(N299), .Y(n111) );
  clknd2d1_hd U395 ( .A(n19), .B(n18), .Y(N225) );
  clknd2d1_hd U397 ( .A(n23), .B(n19), .Y(N223) );
  mx2d1_hd U398 ( .D0(r_pstate[2]), .D1(N302), .S(N299), .Y(n110) );
  or2d1_hd U399 ( .A(N334), .B(N339), .Y(N340) );
  mx2d1_hd U410 ( .D0(r_data_counter[1]), .D1(N295), .S(N293), .Y(n109) );
  mx2d1_hd U411 ( .D0(gt_x_1_n7), .D1(N296), .S(N293), .Y(n113) );
  xo2d1_hd U412 ( .A(add_x_2_n1), .B(gt_x_1_n7), .Y(N200) );
  mx2d1_hd U422 ( .D0(r_pstate[0]), .D1(N300), .S(N299), .Y(n112) );
  scg2d1_hd U423 ( .A(N62), .B(n117), .C(n122), .D(N215), .Y(n13) );
  or2d1_hd U424 ( .A(w_uart_data_rx_valid), .B(i_CORE_BUSY), .Y(alt45_n18) );
  clknd2d1_hd U425 ( .A(n117), .B(w_uart_data_rx_valid), .Y(n18) );
  ivd1_hd U426 ( .A(w_uart_data_rx_valid), .Y(N62) );
  ad2d1_hd U427 ( .A(w_uart_data_rx_valid), .B(alt45_n63), .Y(N305) );
  ivd4_hd U428 ( .A(w_rst), .Y(n5) );
  scg6d1_hd U431 ( .A(gt_x_1_n5), .B(r_data_counter[0]), .C(gt_x_1_n7), .Y(
        n116) );
  nr2d1_hd U432 ( .A(N39), .B(N36), .Y(n117) );
  or2d1_hd U433 ( .A(N305), .B(n123), .Y(N386) );
  ad2d1_hd U434 ( .A(gt_x_3_n5), .B(r_data_counter[0]), .Y(n118) );
  nr2d1_hd U435 ( .A(N355), .B(N380), .Y(n119) );
  nr2d1_hd U436 ( .A(N42), .B(r_pstate[0]), .Y(n120) );
  nr2d1_hd U437 ( .A(N312), .B(N318), .Y(n121) );
  nr2d1_hd U438 ( .A(i_UART_DATA_TX_VALID), .B(alt45_n18), .Y(n123) );
  nr2d1_hd U439 ( .A(i_UART_DATA_TX_VALID), .B(w_uart_data_rx_valid), .Y(n124)
         );
  or2d1_hd U440 ( .A(w_uart_data_rx_valid), .B(n124), .Y(N120) );
  or2d1_hd U441 ( .A(N47), .B(N50), .Y(n125) );
  ivd1_hd U442 ( .A(r_pstate[2]), .Y(N34) );
  nr2d1_hd U443 ( .A(N127), .B(N351), .Y(n126) );
  nr2d1_hd U444 ( .A(N355), .B(N372), .Y(n127) );
  nr2d1_hd U445 ( .A(N355), .B(N361), .Y(n128) );
  ivd1_hd U446 ( .A(r_data_counter[1]), .Y(gt_x_1_n9) );
  ivd1_hd U447 ( .A(w_uart_data_tx_done), .Y(N215) );
  nr2d1_hd U448 ( .A(N312), .B(N330), .Y(n129) );
  ivd1_hd U449 ( .A(gt_x_1_n7), .Y(gt_x_3_n7) );
  nr2d1_hd U450 ( .A(r_uart_data_tx_shift[48]), .B(N340), .Y(n130) );
  ivd1_hd U451 ( .A(n118), .Y(N214) );
  nr2d1_hd U452 ( .A(r_lstate[0]), .B(N322), .Y(n131) );
  SNPS_CLOCK_GATE_HIGH_uart_controller_8 clk_gate_o_UART_DATA_RX_reg_15__0 ( 
        .CLK(i_CLK), .EN(N298), .ENCLK(n268), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_uart_controller_9 clk_gate_o_UART_DATA_RX_reg_7__0 ( 
        .CLK(i_CLK), .EN(N297), .ENCLK(n267), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_uart_controller_10 clk_gate_r_uart_data_tx_valid_reg_0 ( 
        .CLK(i_CLK), .EN(N227), .ENCLK(n266), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_uart_controller_11 clk_gate_r_uart_data_tx_shift_reg_7__0 ( 
        .CLK(i_CLK), .EN(N236), .ENCLK(n265), .TE(1'b0) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(n112), .CK(i_CLK), .RN(n5), .Q(r_pstate[0])
         );
  fd2qd1_hd o_UART_DATA_RX_reg_15_ ( .D(N134), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[15]) );
  fd2qd1_hd o_UART_DATA_RX_reg_14_ ( .D(N133), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[14]) );
  fd2qd1_hd o_UART_DATA_RX_reg_13_ ( .D(N132), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[13]) );
  fd2qd1_hd o_UART_DATA_RX_reg_12_ ( .D(N131), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[12]) );
  fd2qd1_hd o_UART_DATA_RX_reg_11_ ( .D(N130), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[11]) );
  fd2qd1_hd o_UART_DATA_RX_reg_10_ ( .D(N129), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[10]) );
  fd2qd1_hd o_UART_DATA_RX_reg_9_ ( .D(N128), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[9]) );
  fd2qd1_hd o_UART_DATA_RX_reg_8_ ( .D(N127), .CK(n268), .RN(n5), .Q(
        o_UART_DATA_RX[8]) );
  fd2qd1_hd o_UART_DATA_RX_reg_7_ ( .D(N134), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[7]) );
  fd2qd1_hd o_UART_DATA_RX_reg_6_ ( .D(N133), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[6]) );
  fd2qd1_hd o_UART_DATA_RX_reg_3_ ( .D(N130), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[3]) );
  fd2qd1_hd o_UART_DATA_RX_reg_2_ ( .D(N129), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[2]) );
  fd2qd1_hd o_UART_DATA_RX_reg_5_ ( .D(N132), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[5]) );
  fd2qd1_hd o_UART_DATA_RX_reg_4_ ( .D(N131), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[4]) );
  fd2qd1_hd o_UART_DATA_RX_reg_1_ ( .D(N128), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[1]) );
  fd2qd1_hd o_UART_DATA_RX_reg_0_ ( .D(N127), .CK(n267), .RN(n5), .Q(
        o_UART_DATA_RX[0]) );
  fd2qd1_hd r_uart_data_tx_valid_reg ( .D(n125), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx_valid) );
  fd2qd1_hd r_lstate_reg_1_ ( .D(n269), .CK(i_CLK), .RN(n5), .Q(r_lstate[1])
         );
  fd2qd1_hd r_uart_data_tx_reg_7_ ( .D(N235), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[7]) );
  fd2qd1_hd r_uart_data_tx_reg_6_ ( .D(N234), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[6]) );
  fd2qd1_hd r_uart_data_tx_reg_5_ ( .D(N233), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[5]) );
  fd2qd1_hd r_uart_data_tx_reg_4_ ( .D(N232), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[4]) );
  fd2qd1_hd r_uart_data_tx_reg_3_ ( .D(N231), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[3]) );
  fd2qd1_hd r_uart_data_tx_reg_2_ ( .D(N230), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[2]) );
  fd2qd1_hd r_uart_data_tx_reg_1_ ( .D(N229), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[1]) );
  fd2qd1_hd r_uart_data_tx_reg_0_ ( .D(N228), .CK(n266), .RN(n5), .Q(
        r_uart_data_tx[0]) );
  fd2qd1_hd r_lstate_reg_0_ ( .D(n270), .CK(i_CLK), .RN(n5), .Q(r_lstate[0])
         );
  fd2qd1_hd r_uart_data_tx_shift_reg_52_ ( .D(n328), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[52]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_23_ ( .D(n299), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[23]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_22_ ( .D(n298), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[22]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_21_ ( .D(n297), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[21]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_20_ ( .D(n296), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[20]) );
  fd2qd1_hd r_data_counter_reg_0_ ( .D(n271), .CK(i_CLK), .RN(n5), .Q(
        r_data_counter[0]) );
  fd2qd1_hd r_data_counter_reg_2_ ( .D(n113), .CK(i_CLK), .RN(n5), .Q(
        gt_x_1_n7) );
  fd2qd1_hd r_data_counter_reg_1_ ( .D(n109), .CK(i_CLK), .RN(n5), .Q(
        r_data_counter[1]) );
  fd2qd1_hd o_UART_DATA_RX_VALID_reg ( .D(n273), .CK(i_CLK), .RN(n5), .Q(
        o_UART_DATA_RX_VALID) );
  fd2qd1_hd r_pstate_reg_2_ ( .D(n110), .CK(i_CLK), .RN(n5), .Q(r_pstate[2])
         );
  fd2qd1_hd o_UART_DATA_TX_READY_reg ( .D(n272), .CK(i_CLK), .RN(n5), .Q(
        o_UART_DATA_TX_READY) );
  fd2qd1_hd r_uart_data_tx_shift_reg_55_ ( .D(n331), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[55]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_54_ ( .D(n330), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[54]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_53_ ( .D(n329), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[53]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_51_ ( .D(n327), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[51]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_50_ ( .D(n326), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[50]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_49_ ( .D(n325), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[49]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_48_ ( .D(n324), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[48]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_47_ ( .D(n323), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[47]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_46_ ( .D(n322), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[46]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_45_ ( .D(n321), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[45]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_44_ ( .D(n320), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[44]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_43_ ( .D(n319), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[43]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_42_ ( .D(n318), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[42]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_41_ ( .D(n317), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[41]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_40_ ( .D(n316), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[40]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_39_ ( .D(n315), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[39]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_38_ ( .D(n314), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[38]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_37_ ( .D(n313), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[37]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_36_ ( .D(n312), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[36]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_35_ ( .D(n311), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[35]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_34_ ( .D(n310), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[34]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_33_ ( .D(n309), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[33]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_32_ ( .D(n308), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[32]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_31_ ( .D(n307), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[31]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_30_ ( .D(n306), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[30]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_29_ ( .D(n305), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[29]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_28_ ( .D(n304), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[28]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_27_ ( .D(n303), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[27]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_26_ ( .D(n302), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[26]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_25_ ( .D(n301), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[25]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_24_ ( .D(n300), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[24]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_19_ ( .D(n295), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[19]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_18_ ( .D(n294), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[18]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_17_ ( .D(n293), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[17]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_16_ ( .D(n292), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[16]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_15_ ( .D(n291), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[15]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_14_ ( .D(n290), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[14]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_13_ ( .D(n289), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[13]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_12_ ( .D(n288), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[12]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_11_ ( .D(n287), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[11]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_10_ ( .D(n286), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[10]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_9_ ( .D(n285), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[9]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_8_ ( .D(n284), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[8]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_7_ ( .D(N244), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[7]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_5_ ( .D(N242), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[5]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_4_ ( .D(N241), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[4]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_3_ ( .D(N240), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[3]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_1_ ( .D(N238), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[1]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_0_ ( .D(N237), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[0]) );
  fd2qd1_hd r_pstate_reg_1_ ( .D(n111), .CK(i_CLK), .RN(n5), .Q(r_pstate[1])
         );
  fd2qd1_hd r_uart_data_tx_shift_reg_2_ ( .D(N239), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[2]) );
  fd2qd1_hd r_uart_data_tx_shift_reg_6_ ( .D(N243), .CK(n265), .RN(n5), .Q(
        r_uart_data_tx_shift[6]) );
  nr2d4_hd U1 ( .A(n19), .B(n20), .Y(n10) );
  nr2d1_hd U2 ( .A(N51), .B(N36), .Y(n122) );
  scg6d1_hd U3 ( .A(n122), .B(w_uart_data_tx_done), .C(N38), .Y(N236) );
  scg2d1_hd U4 ( .A(i_UART_DATA_TX[8]), .B(n10), .C(r_uart_data_tx_shift[0]), 
        .D(n277), .Y(n284) );
  scg2d1_hd U6 ( .A(i_UART_DATA_TX[9]), .B(n10), .C(r_uart_data_tx_shift[1]), 
        .D(n277), .Y(n285) );
  scg2d1_hd U7 ( .A(i_UART_DATA_TX[10]), .B(n10), .C(r_uart_data_tx_shift[2]), 
        .D(n277), .Y(n286) );
  scg2d1_hd U9 ( .A(i_UART_DATA_TX[11]), .B(n10), .C(r_uart_data_tx_shift[3]), 
        .D(n276), .Y(n287) );
  scg2d1_hd U11 ( .A(i_UART_DATA_TX[12]), .B(n10), .C(r_uart_data_tx_shift[4]), 
        .D(n276), .Y(n288) );
  scg2d1_hd U12 ( .A(i_UART_DATA_TX[13]), .B(n10), .C(r_uart_data_tx_shift[5]), 
        .D(n277), .Y(n289) );
  scg2d1_hd U13 ( .A(i_UART_DATA_TX[14]), .B(n10), .C(r_uart_data_tx_shift[6]), 
        .D(n278), .Y(n290) );
  scg2d1_hd U19 ( .A(i_UART_DATA_TX[15]), .B(n10), .C(r_uart_data_tx_shift[7]), 
        .D(n278), .Y(n291) );
  scg2d1_hd U22 ( .A(i_UART_DATA_TX[16]), .B(n10), .C(r_uart_data_tx_shift[8]), 
        .D(n278), .Y(n292) );
  scg2d1_hd U29 ( .A(i_UART_DATA_TX[17]), .B(n10), .C(r_uart_data_tx_shift[9]), 
        .D(n276), .Y(n293) );
  scg2d1_hd U30 ( .A(i_UART_DATA_TX[18]), .B(n10), .C(r_uart_data_tx_shift[10]), .D(n277), .Y(n294) );
  scg2d1_hd U31 ( .A(i_UART_DATA_TX[19]), .B(n10), .C(r_uart_data_tx_shift[11]), .D(n276), .Y(n295) );
  scg2d1_hd U32 ( .A(i_UART_DATA_TX[24]), .B(n10), .C(r_uart_data_tx_shift[16]), .D(n278), .Y(n300) );
  scg2d1_hd U33 ( .A(i_UART_DATA_TX[25]), .B(n10), .C(r_uart_data_tx_shift[17]), .D(n277), .Y(n301) );
  scg2d1_hd U34 ( .A(i_UART_DATA_TX[26]), .B(n10), .C(r_uart_data_tx_shift[18]), .D(n278), .Y(n302) );
  scg2d1_hd U35 ( .A(i_UART_DATA_TX[27]), .B(n10), .C(r_uart_data_tx_shift[19]), .D(n277), .Y(n303) );
  scg2d1_hd U36 ( .A(i_UART_DATA_TX[28]), .B(n10), .C(r_uart_data_tx_shift[20]), .D(n278), .Y(n304) );
  scg2d1_hd U37 ( .A(i_UART_DATA_TX[29]), .B(n10), .C(r_uart_data_tx_shift[21]), .D(n278), .Y(n305) );
  scg2d1_hd U38 ( .A(i_UART_DATA_TX[30]), .B(n10), .C(r_uart_data_tx_shift[22]), .D(n276), .Y(n306) );
  scg2d1_hd U39 ( .A(i_UART_DATA_TX[31]), .B(n10), .C(r_uart_data_tx_shift[23]), .D(n278), .Y(n307) );
  scg2d1_hd U40 ( .A(i_UART_DATA_TX[32]), .B(n10), .C(r_uart_data_tx_shift[24]), .D(n278), .Y(n308) );
  scg2d1_hd U41 ( .A(i_UART_DATA_TX[33]), .B(n10), .C(r_uart_data_tx_shift[25]), .D(n276), .Y(n309) );
  scg2d1_hd U42 ( .A(i_UART_DATA_TX[34]), .B(n10), .C(r_uart_data_tx_shift[26]), .D(n277), .Y(n310) );
  scg2d1_hd U43 ( .A(i_UART_DATA_TX[35]), .B(n10), .C(r_uart_data_tx_shift[27]), .D(n278), .Y(n311) );
  scg2d1_hd U44 ( .A(i_UART_DATA_TX[36]), .B(n10), .C(r_uart_data_tx_shift[28]), .D(n278), .Y(n312) );
  scg2d1_hd U45 ( .A(i_UART_DATA_TX[37]), .B(n10), .C(r_uart_data_tx_shift[29]), .D(n276), .Y(n313) );
  scg2d1_hd U46 ( .A(i_UART_DATA_TX[38]), .B(n10), .C(r_uart_data_tx_shift[30]), .D(n276), .Y(n314) );
  scg2d1_hd U47 ( .A(i_UART_DATA_TX[39]), .B(n10), .C(r_uart_data_tx_shift[31]), .D(n276), .Y(n315) );
  scg2d1_hd U48 ( .A(i_UART_DATA_TX[40]), .B(n10), .C(r_uart_data_tx_shift[32]), .D(n276), .Y(n316) );
  scg2d1_hd U49 ( .A(i_UART_DATA_TX[41]), .B(n10), .C(r_uart_data_tx_shift[33]), .D(n278), .Y(n317) );
  scg2d1_hd U50 ( .A(i_UART_DATA_TX[42]), .B(n10), .C(r_uart_data_tx_shift[34]), .D(n276), .Y(n318) );
  scg2d1_hd U51 ( .A(i_UART_DATA_TX[43]), .B(n10), .C(r_uart_data_tx_shift[35]), .D(n278), .Y(n319) );
  scg2d1_hd U52 ( .A(i_UART_DATA_TX[44]), .B(n10), .C(r_uart_data_tx_shift[36]), .D(n277), .Y(n320) );
  scg2d1_hd U53 ( .A(i_UART_DATA_TX[45]), .B(n10), .C(r_uart_data_tx_shift[37]), .D(n277), .Y(n321) );
  scg2d1_hd U54 ( .A(i_UART_DATA_TX[46]), .B(n10), .C(r_uart_data_tx_shift[38]), .D(n277), .Y(n322) );
  scg2d1_hd U55 ( .A(i_UART_DATA_TX[47]), .B(n10), .C(r_uart_data_tx_shift[39]), .D(n276), .Y(n323) );
  scg2d1_hd U56 ( .A(i_UART_DATA_TX[48]), .B(n10), .C(r_uart_data_tx_shift[40]), .D(n277), .Y(n324) );
  scg2d1_hd U57 ( .A(i_UART_DATA_TX[49]), .B(n10), .C(r_uart_data_tx_shift[41]), .D(n277), .Y(n325) );
  scg2d1_hd U58 ( .A(i_UART_DATA_TX[50]), .B(n10), .C(r_uart_data_tx_shift[42]), .D(n278), .Y(n326) );
  scg2d1_hd U59 ( .A(i_UART_DATA_TX[51]), .B(n10), .C(r_uart_data_tx_shift[43]), .D(n277), .Y(n327) );
  scg2d1_hd U60 ( .A(i_UART_DATA_TX[53]), .B(n10), .C(r_uart_data_tx_shift[45]), .D(n277), .Y(n329) );
  scg2d1_hd U61 ( .A(i_UART_DATA_TX[54]), .B(n10), .C(r_uart_data_tx_shift[46]), .D(n276), .Y(n330) );
  scg2d1_hd U62 ( .A(i_UART_DATA_TX[55]), .B(n10), .C(r_uart_data_tx_shift[47]), .D(n276), .Y(n331) );
  mx2d1_hd U63 ( .D0(o_UART_DATA_TX_READY), .D1(n280), .S(N223), .Y(n272) );
  mx2d1_hd U64 ( .D0(o_UART_DATA_RX_VALID), .D1(n279), .S(N225), .Y(n273) );
  mx2d1_hd U65 ( .D0(r_data_counter[0]), .D1(N294), .S(N293), .Y(n271) );
  scg2d1_hd U66 ( .A(i_UART_DATA_TX[20]), .B(n10), .C(r_uart_data_tx_shift[12]), .D(n277), .Y(n296) );
  scg2d1_hd U67 ( .A(i_UART_DATA_TX[21]), .B(n10), .C(r_uart_data_tx_shift[13]), .D(n278), .Y(n297) );
  scg2d1_hd U68 ( .A(i_UART_DATA_TX[22]), .B(n10), .C(r_uart_data_tx_shift[14]), .D(n278), .Y(n298) );
  scg2d1_hd U69 ( .A(i_UART_DATA_TX[23]), .B(n10), .C(r_uart_data_tx_shift[15]), .D(n276), .Y(n299) );
  scg2d1_hd U70 ( .A(i_UART_DATA_TX[52]), .B(n10), .C(r_uart_data_tx_shift[44]), .D(n276), .Y(n328) );
  mx2d1_hd U71 ( .D0(r_lstate[0]), .D1(N35), .S(n125), .Y(n270) );
  clknd2d1_hd U72 ( .A(n264), .B(N322), .Y(n269) );
  ivd1_hd U73 ( .A(n125), .Y(n264) );
  ivd1_hd U74 ( .A(r_pstate[0]), .Y(N36) );
  scg17d1_hd U75 ( .A(N305), .B(n126), .C(n117), .D(n274), .Y(n279) );
  nd3d1_hd U76 ( .A(w_uart_data_rx_valid), .B(i_CORE_BUSY), .C(n128), .Y(n274)
         );
  scg17d1_hd U85 ( .A(i_CORE_BUSY), .B(N120), .C(N50), .D(n275), .Y(n280) );
  nr2d1_hd U87 ( .A(N47), .B(N386), .Y(n275) );
  ivd1_hd U99 ( .A(N36), .Y(n276) );
  ivd1_hd U102 ( .A(N36), .Y(n277) );
  ivd1_hd U103 ( .A(N36), .Y(n278) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_sensor_core_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module sensor_core ( o_UART_DATA_TX, o_UART_DATA_TX_VALID, 
        i_UART_DATA_TX_READY, i_UART_DATA_RX, i_UART_DATA_RX_VALID, 
        i_MPR121_DATA_OUT, o_MPR121_REG_ADDR, o_MPR121_DATA_IN, 
        o_MPR121_WRITE_ENABLE, o_MPR121_READ_ENABLE, i_MPR121_INIT_SET, 
        i_MPR121_BUSY, i_MPR121_FAIL, o_MPR121_ERROR, 
        i_ADS1292_FILTERED_DATA_OUT, o_ADS1292_CONTROL, o_ADS1292_REG_ADDR, 
        o_ADS1292_DATA_IN, i_ADS1292_REG_DATA_OUT, i_ADS1292_INIT_SET, 
        i_ADS1292_FILTERED_DATA_VALID, o_ADS1292_FILTERED_DATA_ACK, 
        i_ADS1292_BUSY, i_CLK, i_RSTN );
  output [55:0] o_UART_DATA_TX;
  input [15:0] i_UART_DATA_RX;
  input [7:0] i_MPR121_DATA_OUT;
  output [7:0] o_MPR121_REG_ADDR;
  output [7:0] o_MPR121_DATA_IN;
  input [23:0] i_ADS1292_FILTERED_DATA_OUT;
  output [2:0] o_ADS1292_CONTROL;
  output [7:0] o_ADS1292_REG_ADDR;
  output [7:0] o_ADS1292_DATA_IN;
  input [7:0] i_ADS1292_REG_DATA_OUT;
  input i_UART_DATA_TX_READY, i_UART_DATA_RX_VALID, i_MPR121_INIT_SET,
         i_MPR121_BUSY, i_MPR121_FAIL, i_ADS1292_INIT_SET,
         i_ADS1292_FILTERED_DATA_VALID, i_ADS1292_BUSY, i_CLK, i_RSTN;
  output o_UART_DATA_TX_VALID, o_MPR121_WRITE_ENABLE, o_MPR121_READ_ENABLE,
         o_MPR121_ERROR, o_ADS1292_FILTERED_DATA_ACK;
  wire   n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n597, n598, n599, n619, N8, N63, N68, w_rst, r_run_mode, N153,
         N154, N155, N158, N164, N165, N166, N167, N168, N169, N170,
         r_ads_data_send_ready, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N215, N216, N217, N219, N224,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N243, N250, N251, N252, N253, N254,
         N255, r_chip_set, r_ads_chip_set_done, r_run_set, r_mpr_run_set_done,
         r_ads_run_set_done, r_mpr_chip_set, r_mpr_run_set, r_mpr_read_reg,
         r_ads_chip_set, r_ads_read_reg, N274, N275, N276, N277, N279, N282,
         N283, N285, N286, N288, N297, N298, N302, N303, N304, N308, N309,
         N314, N316, N318, N319, N322, N326, N330, N331, N332, N333, N343,
         N344, N345, N346, N347, N350, N351, N352, N353, N354, N355, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N370,
         N371, N372, N373, N374, N377, N378, N379, N380, N383, N384, N385,
         N386, N389, N390, N391, N392, N395, N396, N397, N398, N399, N402,
         N403, N404, N405, N408, N409, N410, N411, N414, N415, N416, N417,
         N420, N421, N422, N423, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N438, N439, N440, N441, N444, N445, N446, N447,
         N448, N451, N452, N453, N454, N457, N458, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N475, N476, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N596, N597,
         N598, N603, N607, N608, N616, N617, N618, N626, N627, N631, N635,
         N636, N637, N638, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N657, N658, N659, N660,
         N661, N662, N663, N664, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N680, N681, N682, N683, N691, N692,
         N693, N694, N695, N696, N697, N698, N700, N701, N702, N703, N707,
         N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N725,
         N728, N741, N742, N743, N744, N747, N748, N749, N751, N752, N753,
         N756, N757, N760, N761, N764, N765, N766, N767, N768, N769, N770,
         N773, N774, N777, N778, N781, N782, N785, N786, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N801, N802, N803, N804,
         N805, N806, N807, N808, N809, N810, N811, N812, N905, N906, N907,
         N914, N915, N921, N922, N923, N929, N932, N933, N936, N937, N938,
         N939, N940, N941, N942, N943, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N958, N959, N960, N961, N962,
         N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973,
         N974, N975, N976, N977, N978, N979, N980, N981, N985, N986, N987,
         N988, N990, N991, N992, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1013, N1014, N1016, N1017, N1018, N1019, N1020, N1021,
         N1022, N1023, N1024, N1025, N1026, N1027, N1029, N1030, N1032, N1038,
         N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1049, N1050,
         N1052, N1055, N1056, N1059, N1064, N1065, N1068, N1069, N1070, N1071,
         N1072, N1073, N1075, N1076, N1077, N1078, N1079, N1087, N1088, N1091,
         N1092, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1104,
         N1105, N1106, N1108, N1109, N1110, N1111, N1113, N1114, N1115, N1116,
         N1117, N1118, N1119, N1120, N1123, N1124, N1125, N1126, N1127, N1128,
         N1131, N1132, N1133, N1134, N1136, N1137, N1140, N1141, N1142, N1144,
         N1145, N1146, N1149, N1150, N1151, N1153, N1154, N1155, N1157, N1158,
         N1159, N1161, N1162, N1163, N1165, N1166, N1167, N1169, N1170, N1171,
         N1172, N1173, N1174, N1175, N1177, N1178, N1181, N1182, N1183, N1185,
         N1186, N1187, N1189, N1190, N1191, N1193, N1194, N1195, N1197, N1198,
         N1199, N1201, N1202, N1205, N1206, N1207, N1209, N1210, N1211, N1213,
         N1214, N1229, N1238, N1239, N1240, N1243, N1244, N1256, N1257, N1258,
         N1259, N1270, N1271, N1273, N1275, N1278, N1282, N1286, N1289, N1290,
         N1291, N1294, N1299, N1303, N1311, N1312, N1313, N1314, N1315, N1316,
         N1317, N1318, N1319, alt36_n60, alt36_n63, alt36_n127, alt36_n128,
         alt36_n129, alt36_n159, alt36_n287, alt36_n288, alt36_n298,
         alt36_n301, alt36_n329, alt36_n332, alt36_n508, alt36_n509,
         alt36_n510, alt36_n511, alt36_n513, add_x_150_n2, add_x_150_n1,
         gt_x_149_n18, gt_x_149_n17, gt_x_149_n15, gt_x_149_n14, gt_x_149_n13,
         gt_x_149_n12, gt_x_149_n10, gt_x_149_n9, add_x_148_n2, add_x_148_n1,
         gt_x_147_n15, gt_x_147_n13, gt_x_147_n12, add_x_62_n2, add_x_62_n1,
         gt_x_61_n18, gt_x_61_n17, gt_x_61_n15, gt_x_61_n14, gt_x_61_n13,
         gt_x_61_n12, gt_x_61_n7, add_x_60_n2, add_x_60_n1, add_x_1_n2,
         add_x_1_n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15,
         n16, n18, n20, n21, n22, n23, n36, n37, n38, n39, n40, n42, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n68, n69, n70, n71, n72, n73, n74, n76,
         n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n166, n168, n170, n174, n178, n180, n182, n184, n185,
         n186, n187, n188, n190, n191, n192, n193, n195, n196, n197, n198,
         n199, n200, n202, n203, n204, n205, n206, n208, n209, n210, n211,
         n212, n213, n491, n492, n512, n513, n514, n516, n517, n518, n519,
         n520, n521, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n565,
         n566, n569, n570, n571, n572, n573, n574, r_mpr_lstate_1_, n67, n75,
         n78, n92, n154, n175, n177, n183, n189, n194, n201, n207, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n290, n291, n292, n293, n294, n295, n296, n297, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n337, n338, n339, n340,
         n341, n342, n343, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n390, n391, n392, n393, n394, n395, n404, n405,
         n406, n407, n408, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n636, n767, n768, n906, n908, n909, n910, n911, n912, n914,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n961;
  wire   [1:0] r_uart_pstate;
  wire   [3:0] r_uart_clk_counter;
  wire   [11:0] r_mpr_touch_status;
  wire   [7:0] r_ads_reg_addr;
  wire   [7:0] r_mpr_reg_addr;
  wire   [2:1] r_core_pstate;
  wire   [5:0] r_mpr_pstate;
  wire   [3:0] r_mpr_set_counter;
  wire   [7:0] r_mpr_first_param;
  wire   [2:0] r_mpr_clk_counter;
  wire   [7:0] r_mpr_second_param;
  wire   [3:0] r_ads_set_counter;
  wire   [7:0] r_ads_first_param;
  wire   [2:0] r_ads_clk_counter;
  wire   [7:0] r_ads_second_param;

  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  had1_hd add_x_150_U3 ( .A(n407), .B(n404), .CO(add_x_150_n2), .S(N921) );
  had1_hd add_x_150_U2 ( .A(n406), .B(add_x_150_n2), .CO(add_x_150_n1), .S(
        N922) );
  nr2d1_hd gt_x_149_U17 ( .A(n407), .B(gt_x_149_n15), .Y(gt_x_149_n13) );
  ao21d1_hd gt_x_149_U16 ( .A(gt_x_149_n13), .B(n404), .C(gt_x_149_n14), .Y(
        gt_x_149_n12) );
  had1_hd add_x_148_U3 ( .A(n342), .B(n337), .CO(add_x_148_n2), .S(N905) );
  had1_hd add_x_148_U2 ( .A(n207), .B(add_x_148_n2), .CO(add_x_148_n1), .S(
        N906) );
  nr2d1_hd gt_x_147_U17 ( .A(N1076), .B(n207), .Y(gt_x_147_n13) );
  ao21d1_hd gt_x_147_U16 ( .A(gt_x_147_n13), .B(n337), .C(n207), .Y(
        gt_x_147_n12) );
  had1_hd add_x_62_U3 ( .A(n394), .B(n390), .CO(add_x_62_n2), .S(N616) );
  had1_hd add_x_62_U2 ( .A(n393), .B(add_x_62_n2), .CO(add_x_62_n1), .S(N617)
         );
  nr2d1_hd gt_x_61_U17 ( .A(n394), .B(gt_x_61_n15), .Y(gt_x_61_n13) );
  ao21d1_hd gt_x_61_U16 ( .A(gt_x_61_n13), .B(n390), .C(gt_x_61_n14), .Y(
        gt_x_61_n12) );
  had1_hd add_x_60_U3 ( .A(n214), .B(n408), .CO(add_x_60_n2), .S(N596) );
  had1_hd add_x_60_U2 ( .A(n340), .B(add_x_60_n2), .CO(add_x_60_n1), .S(N597)
         );
  had1_hd add_x_1_U3 ( .A(n351), .B(n352), .CO(add_x_1_n2), .S(N164) );
  had1_hd add_x_1_U2 ( .A(n353), .B(add_x_1_n2), .CO(add_x_1_n1), .S(N165) );
  or2d1_hd U5 ( .A(N462), .B(o_MPR121_ERROR), .Y(n599) );
  or2d1_hd U6 ( .A(n3), .B(n468), .Y(r_ads_chip_set_done) );
  nd2bd1_hd U12 ( .AN(n516), .B(n4), .Y(N992) );
  or3d1_hd U13 ( .A(n5), .B(n513), .C(n546), .Y(N991) );
  nr2d1_hd U15 ( .A(n545), .B(n5), .Y(n4) );
  nd3d1_hd U16 ( .A(n202), .B(n7), .C(N767), .Y(n5) );
  ivd1_hd U17 ( .A(n2), .Y(N603) );
  nr2d1_hd U18 ( .A(N1068), .B(n561), .Y(n2) );
  ivd1_hd U19 ( .A(N355), .Y(N63) );
  scg22d1_hd U22 ( .A(n9), .B(n10), .C(n154), .D(i_UART_DATA_TX_READY), .Y(
        n192) );
  ivd1_hd U28 ( .A(n447), .Y(n10) );
  or4d1_hd U30 ( .A(N431), .B(n534), .C(n553), .D(n13), .Y(N1289) );
  or4d1_hd U31 ( .A(n535), .B(n14), .C(n516), .D(n513), .Y(N1282) );
  scg13d1_hd U32 ( .A(n545), .B(N751), .C(n15), .Y(N1275) );
  nd4d1_hd U33 ( .A(n16), .B(n148), .C(N430), .D(n18), .Y(N1270) );
  ivd1_hd U34 ( .A(n548), .Y(n18) );
  scg13d1_hd U36 ( .A(N462), .B(n519), .C(n11), .Y(N1258) );
  nr3d1_hd U37 ( .A(N431), .B(n549), .C(n532), .Y(n11) );
  nr4d1_hd U38 ( .A(n463), .B(N458), .C(N457), .D(N357), .Y(N462) );
  or4d1_hd U40 ( .A(n534), .B(n521), .C(n512), .D(n20), .Y(N1257) );
  ivd1_hd U41 ( .A(n12), .Y(n20) );
  nr2d1_hd U42 ( .A(n548), .B(n514), .Y(n12) );
  nd3bd1_hd U43 ( .AN(n553), .B(N355), .C(n21), .Y(N1256) );
  nd3d1_hd U44 ( .A(n148), .B(n139), .C(n22), .Y(N1244) );
  nr3d1_hd U45 ( .A(n532), .B(n519), .C(n548), .Y(n22) );
  nr2bd1_hd U47 ( .AN(n95), .B(n13), .Y(n21) );
  nd2bd1_hd U48 ( .AN(n544), .B(N362), .Y(n13) );
  nr2d1_hd U49 ( .A(n534), .B(n518), .Y(n16) );
  ivd1_hd U51 ( .A(N751), .Y(n193) );
  nr4d1_hd U54 ( .A(n516), .B(n545), .C(n513), .D(n491), .Y(n23) );
  nd3bd1_hd U56 ( .AN(n535), .B(n203), .C(n15), .Y(N1229) );
  nr2d1_hd U57 ( .A(n530), .B(n14), .Y(n15) );
  ivd1_hd U59 ( .A(n546), .Y(n6) );
  ivd1_hd U60 ( .A(n527), .Y(n7) );
  oa21d1_hd U62 ( .A(gt_x_147_n12), .B(N1075), .C(N751), .Y(n62) );
  nr2d1_hd U63 ( .A(N748), .B(N749), .Y(N751) );
  scg17d1_hd U102 ( .A(n491), .B(N805), .C(n36), .D(n37), .Y(N999) );
  oa21d1_hd U103 ( .A(n541), .B(n38), .C(n39), .Y(n37) );
  ao21d1_hd U104 ( .A(n40), .B(N1155), .C(n523), .Y(n38) );
  oa21d1_hd U105 ( .A(N1172), .B(n42), .C(N1163), .Y(n40) );
  nr2bd1_hd U106 ( .AN(N923), .B(n44), .Y(N988) );
  nr2bd1_hd U107 ( .AN(N922), .B(n44), .Y(N987) );
  nr2bd1_hd U108 ( .AN(N921), .B(n44), .Y(N986) );
  nr2d1_hd U109 ( .A(n404), .B(n44), .Y(N985) );
  ad2d1_hd U110 ( .A(i_ADS1292_FILTERED_DATA_OUT[23]), .B(n542), .Y(N981) );
  ad2d1_hd U111 ( .A(i_ADS1292_FILTERED_DATA_OUT[22]), .B(n542), .Y(N980) );
  ad2d1_hd U112 ( .A(i_ADS1292_FILTERED_DATA_OUT[21]), .B(n542), .Y(N979) );
  ad2d1_hd U113 ( .A(i_ADS1292_FILTERED_DATA_OUT[20]), .B(n542), .Y(N978) );
  ad2d1_hd U114 ( .A(i_ADS1292_FILTERED_DATA_OUT[19]), .B(n542), .Y(N977) );
  ad2d1_hd U115 ( .A(i_ADS1292_FILTERED_DATA_OUT[18]), .B(n542), .Y(N976) );
  ad2d1_hd U116 ( .A(i_ADS1292_FILTERED_DATA_OUT[17]), .B(n542), .Y(N975) );
  ad2d1_hd U117 ( .A(i_ADS1292_FILTERED_DATA_OUT[16]), .B(n542), .Y(N974) );
  ad2d1_hd U118 ( .A(i_ADS1292_FILTERED_DATA_OUT[15]), .B(n542), .Y(N973) );
  ad2d1_hd U119 ( .A(i_ADS1292_FILTERED_DATA_OUT[14]), .B(n542), .Y(N972) );
  ad2d1_hd U120 ( .A(i_ADS1292_FILTERED_DATA_OUT[13]), .B(n542), .Y(N971) );
  ad2d1_hd U121 ( .A(i_ADS1292_FILTERED_DATA_OUT[12]), .B(n542), .Y(N970) );
  ad2d1_hd U122 ( .A(i_ADS1292_FILTERED_DATA_OUT[11]), .B(n542), .Y(N969) );
  ad2d1_hd U123 ( .A(i_ADS1292_FILTERED_DATA_OUT[10]), .B(n542), .Y(N968) );
  ad2d1_hd U124 ( .A(i_ADS1292_FILTERED_DATA_OUT[9]), .B(n542), .Y(N967) );
  ad2d1_hd U125 ( .A(i_ADS1292_FILTERED_DATA_OUT[8]), .B(n542), .Y(N966) );
  ad2d1_hd U126 ( .A(i_ADS1292_FILTERED_DATA_OUT[7]), .B(n542), .Y(N965) );
  ad2d1_hd U127 ( .A(i_ADS1292_FILTERED_DATA_OUT[6]), .B(n542), .Y(N964) );
  ad2d1_hd U128 ( .A(i_ADS1292_FILTERED_DATA_OUT[5]), .B(n542), .Y(N963) );
  ad2d1_hd U129 ( .A(i_ADS1292_FILTERED_DATA_OUT[4]), .B(n542), .Y(N962) );
  ad2d1_hd U130 ( .A(i_ADS1292_FILTERED_DATA_OUT[3]), .B(n542), .Y(N961) );
  ad2d1_hd U131 ( .A(i_ADS1292_FILTERED_DATA_OUT[2]), .B(n542), .Y(N960) );
  ad2d1_hd U132 ( .A(i_ADS1292_FILTERED_DATA_OUT[1]), .B(n542), .Y(N959) );
  ad2d1_hd U133 ( .A(i_ADS1292_FILTERED_DATA_OUT[0]), .B(n542), .Y(N958) );
  nr3d1_hd U134 ( .A(n45), .B(n46), .C(n42), .Y(N956) );
  ad3d1_hd U135 ( .A(N1079), .B(n47), .C(N751), .Y(N955) );
  oa21d1_hd U136 ( .A(n48), .B(n49), .C(N1111), .Y(n47) );
  nr2d1_hd U137 ( .A(n541), .B(n50), .Y(N954) );
  scg9d1_hd U138 ( .A(n46), .B(n48), .C(n51), .Y(n50) );
  nr4d1_hd U140 ( .A(N1171), .B(n54), .C(n45), .D(n55), .Y(N953) );
  ivd1_hd U141 ( .A(n56), .Y(N952) );
  oa21d1_hd U142 ( .A(N1195), .B(n57), .C(n56), .Y(N951) );
  oa22ad1_hd U143 ( .A(n523), .B(n57), .C(n541), .D(n52), .Y(N950) );
  or2d1_hd U144 ( .A(n58), .B(n46), .Y(n57) );
  nr4d1_hd U145 ( .A(n45), .B(n46), .C(n517), .D(n59), .Y(N949) );
  ivd1_hd U146 ( .A(n60), .Y(n59) );
  nr2bd1_hd U148 ( .AN(N907), .B(n62), .Y(N948) );
  nr2bd1_hd U149 ( .AN(N906), .B(n62), .Y(N947) );
  nr2bd1_hd U150 ( .AN(N905), .B(n62), .Y(N946) );
  nr2d1_hd U151 ( .A(n337), .B(n62), .Y(N945) );
  ad2d1_hd U152 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[7]), .Y(N943) );
  ad2d1_hd U153 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[6]), .Y(N942) );
  ad2d1_hd U154 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[5]), .Y(N941) );
  ad2d1_hd U155 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[4]), .Y(N940) );
  ad2d1_hd U156 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[3]), .Y(N939) );
  ad2d1_hd U157 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[2]), .Y(N938) );
  ad2d1_hd U158 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[1]), .Y(N937) );
  ad2d1_hd U159 ( .A(n527), .B(i_ADS1292_REG_DATA_OUT[0]), .Y(N936) );
  ivd1_hd U160 ( .A(n63), .Y(N812) );
  ivd1_hd U161 ( .A(n64), .Y(N811) );
  nr2d1_hd U162 ( .A(n65), .B(n66), .Y(N805) );
  ao22d1_hd U169 ( .A(N627), .B(n531), .C(N608), .D(n74), .Y(n72) );
  ivd1_hd U172 ( .A(n77), .Y(n74) );
  scg18d1_hd U175 ( .A(n529), .B(N607), .C(N1294), .D(n80), .E(n81), .Y(n79)
         );
  ao211d1_hd U177 ( .A(n521), .B(n533), .C(n83), .D(n76), .Y(n81) );
  ivd1_hd U179 ( .A(n70), .Y(n83) );
  ao211d1_hd U181 ( .A(n518), .B(N607), .C(n68), .D(N1291), .Y(n82) );
  scg18d1_hd U183 ( .A(n531), .B(N626), .C(N1271), .D(n87), .E(n80), .Y(n86)
         );
  nd2bd1_hd U184 ( .AN(n556), .B(n519), .Y(n87) );
  ao211d1_hd U186 ( .A(n562), .B(n521), .C(n90), .D(n91), .Y(n89) );
  oa211d1_hd U187 ( .A(n77), .B(alt36_n159), .C(n80), .D(n84), .Y(n91) );
  nr2d1_hd U189 ( .A(n529), .B(n518), .Y(n77) );
  nr2d1_hd U190 ( .A(n555), .B(n95), .Y(n90) );
  nr2d1_hd U191 ( .A(n69), .B(N1286), .Y(n88) );
  ivd1_hd U192 ( .A(n73), .Y(n69) );
  oa21d1_hd U196 ( .A(n93), .B(n94), .C(n95), .Y(N716) );
  ivd1_hd U200 ( .A(n95), .Y(N713) );
  ivd1_hd U201 ( .A(n71), .Y(N712) );
  nr2d1_hd U203 ( .A(n98), .B(n99), .Y(n97) );
  nr3d1_hd U204 ( .A(n558), .B(n100), .C(n101), .Y(n98) );
  scg14d1_hd U206 ( .A(n529), .B(n96), .C(n95), .Y(N710) );
  nr2d1_hd U211 ( .A(n95), .B(n102), .Y(N698) );
  oa21d1_hd U212 ( .A(n95), .B(n103), .C(n104), .Y(N697) );
  ao22d1_hd U216 ( .A(N63), .B(n100), .C(n526), .D(N486), .Y(n107) );
  scg15d1_hd U218 ( .A(n526), .B(N485), .C(n104), .D(n110), .Y(N694) );
  nd3d1_hd U219 ( .A(N63), .B(n111), .C(n112), .Y(n110) );
  ao211d1_hd U220 ( .A(N63), .B(n113), .C(N1299), .D(N644), .Y(n104) );
  oa211d1_hd U221 ( .A(n114), .B(N355), .C(n108), .D(n115), .Y(N693) );
  ao211d1_hd U223 ( .A(N1134), .B(n116), .C(n117), .D(n118), .Y(n114) );
  oa211d1_hd U224 ( .A(n119), .B(n120), .C(N1142), .D(N1151), .Y(n116) );
  nd2bd1_hd U226 ( .AN(n121), .B(n122), .Y(n101) );
  ivd1_hd U227 ( .A(n123), .Y(n111) );
  scg17d1_hd U228 ( .A(n526), .B(N483), .C(n124), .D(n108), .Y(N692) );
  ivd1_hd U229 ( .A(N1299), .Y(n108) );
  ao211d1_hd U230 ( .A(N1134), .B(n125), .C(n117), .D(n126), .Y(n124) );
  oa211d1_hd U231 ( .A(n127), .B(n119), .C(N1142), .D(N1151), .Y(n125) );
  ao21d1_hd U232 ( .A(n122), .B(n121), .C(n123), .Y(n127) );
  nr2d1_hd U234 ( .A(n128), .B(n129), .Y(n122) );
  oa21d1_hd U235 ( .A(n130), .B(N355), .C(n131), .Y(N691) );
  ao22d1_hd U236 ( .A(n392), .B(n519), .C(n526), .D(N482), .Y(n131) );
  ao211d1_hd U237 ( .A(N1106), .B(n132), .C(n133), .D(n118), .Y(n130) );
  ad4d1_hd U238 ( .A(N1151), .B(N1167), .C(N1106), .D(n134), .Y(n133) );
  oa21d1_hd U239 ( .A(n135), .B(n136), .C(N1175), .Y(n134) );
  ao211d1_hd U240 ( .A(N1199), .B(N1211), .C(n137), .D(n128), .Y(n135) );
  oa211d1_hd U241 ( .A(N1159), .B(n138), .C(N1142), .D(N1134), .Y(n132) );
  ivd1_hd U242 ( .A(N1151), .Y(n138) );
  nr2bd1_hd U243 ( .AN(N618), .B(n80), .Y(N683) );
  nr2bd1_hd U244 ( .AN(N617), .B(n80), .Y(N682) );
  nr2bd1_hd U245 ( .AN(N616), .B(n80), .Y(N681) );
  nr2d1_hd U246 ( .A(n390), .B(n80), .Y(N680) );
  ad2d1_hd U248 ( .A(n264), .B(N68), .Y(N678) );
  ad2d1_hd U249 ( .A(n265), .B(N68), .Y(N677) );
  ad2d1_hd U250 ( .A(n266), .B(N68), .Y(N676) );
  ad2d1_hd U251 ( .A(n267), .B(N68), .Y(N675) );
  ad2d1_hd U252 ( .A(n268), .B(N68), .Y(N674) );
  ad2d1_hd U253 ( .A(n269), .B(N68), .Y(N673) );
  ad2d1_hd U254 ( .A(n215), .B(N68), .Y(N672) );
  ad2d1_hd U255 ( .A(n216), .B(N68), .Y(N671) );
  ad2d1_hd U256 ( .A(n217), .B(N68), .Y(N670) );
  ad2d1_hd U257 ( .A(n218), .B(N68), .Y(N669) );
  ad2d1_hd U258 ( .A(n219), .B(N68), .Y(N668) );
  ad2d1_hd U259 ( .A(n220), .B(N68), .Y(N667) );
  nr2d1_hd U260 ( .A(n139), .B(n140), .Y(N664) );
  nr2d1_hd U261 ( .A(n139), .B(n141), .Y(N663) );
  nr2d1_hd U262 ( .A(n139), .B(n142), .Y(N662) );
  nr2d1_hd U263 ( .A(n139), .B(n143), .Y(N661) );
  nr2d1_hd U264 ( .A(n139), .B(n144), .Y(N660) );
  nr2d1_hd U265 ( .A(n139), .B(n145), .Y(N659) );
  nr2d1_hd U266 ( .A(n139), .B(n146), .Y(N658) );
  nr2d1_hd U267 ( .A(n139), .B(n147), .Y(N657) );
  ivd1_hd U268 ( .A(n531), .Y(n139) );
  ivd1_hd U269 ( .A(n85), .Y(N654) );
  nr2d1_hd U272 ( .A(n148), .B(n140), .Y(N653) );
  ivd1_hd U273 ( .A(i_MPR121_DATA_OUT[7]), .Y(n140) );
  nr2d1_hd U274 ( .A(n148), .B(n141), .Y(N652) );
  ivd1_hd U275 ( .A(i_MPR121_DATA_OUT[6]), .Y(n141) );
  nr2d1_hd U276 ( .A(n148), .B(n142), .Y(N651) );
  ivd1_hd U277 ( .A(i_MPR121_DATA_OUT[5]), .Y(n142) );
  nr2d1_hd U278 ( .A(n148), .B(n143), .Y(N650) );
  ivd1_hd U279 ( .A(i_MPR121_DATA_OUT[4]), .Y(n143) );
  nr2d1_hd U280 ( .A(n148), .B(n144), .Y(N649) );
  ivd1_hd U281 ( .A(i_MPR121_DATA_OUT[3]), .Y(n144) );
  nr2d1_hd U282 ( .A(n148), .B(n145), .Y(N648) );
  ivd1_hd U283 ( .A(i_MPR121_DATA_OUT[2]), .Y(n145) );
  nr2d1_hd U284 ( .A(n148), .B(n146), .Y(N647) );
  ivd1_hd U285 ( .A(i_MPR121_DATA_OUT[1]), .Y(n146) );
  nr2d1_hd U286 ( .A(n148), .B(n147), .Y(N646) );
  ivd1_hd U287 ( .A(i_MPR121_DATA_OUT[0]), .Y(n147) );
  ivd1_hd U288 ( .A(n529), .Y(n148) );
  ao21d1_hd U289 ( .A(N1073), .B(N1106), .C(N355), .Y(N644) );
  oa21d1_hd U290 ( .A(N355), .B(n149), .C(n150), .Y(N643) );
  oa211d1_hd U292 ( .A(n152), .B(n136), .C(N1175), .D(n153), .Y(n151) );
  ivd1_hd U293 ( .A(N1183), .Y(n136) );
  oa21d1_hd U294 ( .A(n126), .B(n149), .C(N362), .Y(N641) );
  ad2d1_hd U297 ( .A(n137), .B(N1191), .Y(n152) );
  nr2d1_hd U298 ( .A(N1207), .B(n129), .Y(n137) );
  ivd1_hd U299 ( .A(N1199), .Y(n129) );
  nr2d1_hd U300 ( .A(n123), .B(n155), .Y(n109) );
  ivd1_hd U301 ( .A(n105), .Y(n126) );
  nr2d1_hd U302 ( .A(N355), .B(n118), .Y(n105) );
  ivd1_hd U303 ( .A(N1073), .Y(n118) );
  scg16d1_hd U304 ( .A(n153), .B(n156), .C(n150), .Y(N640) );
  nr2d1_hd U305 ( .A(N645), .B(N363), .Y(n150) );
  nr2d1_hd U306 ( .A(N1073), .B(N355), .Y(N645) );
  ao211d1_hd U307 ( .A(N1199), .B(N1207), .C(n128), .D(n123), .Y(n156) );
  ivd1_hd U309 ( .A(N1191), .Y(n128) );
  nr2d1_hd U310 ( .A(N355), .B(n155), .Y(n153) );
  nr2d1_hd U312 ( .A(n117), .B(n113), .Y(n106) );
  ivd1_hd U313 ( .A(N1134), .Y(n113) );
  ivd1_hd U314 ( .A(N1106), .Y(n117) );
  scg12d1_hd U315 ( .A(N1151), .B(N1142), .C(n119), .Y(n112) );
  ad2d1_hd U317 ( .A(N598), .B(n68), .Y(N638) );
  ad2d1_hd U318 ( .A(N597), .B(n68), .Y(N637) );
  ad2d1_hd U319 ( .A(N596), .B(n68), .Y(N636) );
  ivd1_hd U320 ( .A(n99), .Y(n68) );
  nr2d1_hd U321 ( .A(n408), .B(n99), .Y(N635) );
  ivd1_hd U323 ( .A(n102), .Y(N489) );
  ivd1_hd U325 ( .A(n103), .Y(N488) );
  nr2d1_hd U327 ( .A(n157), .B(n158), .Y(N487) );
  nr2d1_hd U328 ( .A(n157), .B(n159), .Y(N486) );
  nr2d1_hd U329 ( .A(n157), .B(n160), .Y(N485) );
  nr2d1_hd U330 ( .A(n157), .B(n161), .Y(N484) );
  nr2d1_hd U331 ( .A(n157), .B(n162), .Y(N483) );
  nr2d1_hd U332 ( .A(n65), .B(n157), .Y(N482) );
  ivd1_hd U333 ( .A(N481), .Y(n157) );
  ao22d1_hd U335 ( .A(n365), .B(n166), .C(N316), .D(N303), .Y(n163) );
  scg14d1_hd U337 ( .A(n168), .B(N308), .C(n911), .Y(N332) );
  ao22d1_hd U340 ( .A(n357), .B(n166), .C(N316), .D(N302), .Y(n170) );
  nr2d1_hd U342 ( .A(alt36_n298), .B(N286), .Y(n166) );
  oa211d1_hd U347 ( .A(n912), .B(n525), .C(N283), .D(n178), .Y(
        r_core_pstate[1]) );
  ao22d1_hd U351 ( .A(n168), .B(n458), .C(n563), .D(n180), .Y(n178) );
  scg14d1_hd U354 ( .A(n168), .B(N309), .C(n911), .Y(N326) );
  ivd1_hd U356 ( .A(N286), .Y(n168) );
  nr2d1_hd U358 ( .A(n447), .B(N286), .Y(N322) );
  nr2d1_hd U359 ( .A(n468), .B(N283), .Y(N319) );
  nr2d1_hd U360 ( .A(n270), .B(N286), .Y(N318) );
  nr2d1_hd U361 ( .A(N286), .B(n180), .Y(N316) );
  ivd1_hd U362 ( .A(n356), .Y(n180) );
  nr2d1_hd U364 ( .A(n457), .B(N283), .Y(N314) );
  oa211d1_hd U366 ( .A(n538), .B(n182), .C(N158), .D(n184), .Y(
        r_uart_pstate[0]) );
  oa211d1_hd U367 ( .A(n185), .B(n186), .C(n182), .D(n187), .Y(N255) );
  ivd1_hd U369 ( .A(N216), .Y(n186) );
  oa211d1_hd U370 ( .A(n9), .B(n185), .C(n182), .D(n190), .Y(N254) );
  scg6d1_hd U374 ( .A(n188), .B(N224), .C(N155), .Y(N253) );
  ivd1_hd U376 ( .A(N158), .Y(n188) );
  nr2bd1_hd U380 ( .AN(i_UART_DATA_RX_VALID), .B(n191), .Y(r_uart_pstate[1])
         );
  ad2d1_hd U381 ( .A(n536), .B(n188), .Y(N243) );
  ad2d1_hd U382 ( .A(N8), .B(i_UART_DATA_RX[15]), .Y(N241) );
  ad2d1_hd U383 ( .A(N8), .B(i_UART_DATA_RX[14]), .Y(N240) );
  ad2d1_hd U384 ( .A(N8), .B(i_UART_DATA_RX[13]), .Y(N239) );
  ad2d1_hd U385 ( .A(N8), .B(i_UART_DATA_RX[12]), .Y(N238) );
  ad2d1_hd U386 ( .A(N8), .B(i_UART_DATA_RX[11]), .Y(N237) );
  ad2d1_hd U387 ( .A(N8), .B(i_UART_DATA_RX[10]), .Y(N236) );
  ad2d1_hd U388 ( .A(N8), .B(i_UART_DATA_RX[9]), .Y(N235) );
  ad2d1_hd U389 ( .A(N8), .B(i_UART_DATA_RX[8]), .Y(N234) );
  ad2d1_hd U390 ( .A(N8), .B(i_UART_DATA_RX[7]), .Y(N233) );
  ad2d1_hd U391 ( .A(N8), .B(i_UART_DATA_RX[6]), .Y(N232) );
  ad2d1_hd U392 ( .A(N8), .B(i_UART_DATA_RX[5]), .Y(N231) );
  ad2d1_hd U393 ( .A(N8), .B(i_UART_DATA_RX[4]), .Y(N230) );
  ad2d1_hd U394 ( .A(N8), .B(i_UART_DATA_RX[3]), .Y(N229) );
  ad2d1_hd U395 ( .A(N8), .B(i_UART_DATA_RX[2]), .Y(N228) );
  ad2d1_hd U396 ( .A(N8), .B(i_UART_DATA_RX[1]), .Y(N227) );
  ad2d1_hd U397 ( .A(N8), .B(i_UART_DATA_RX[0]), .Y(N226) );
  ivd1_hd U398 ( .A(n192), .Y(N219) );
  scg5d1_hd U399 ( .A(N217), .B(n230), .C(n154), .D(n240), .E(n366), .F(N216), 
        .Y(N213) );
  scg5d1_hd U400 ( .A(N217), .B(n229), .C(n154), .D(n241), .E(n367), .F(N216), 
        .Y(N212) );
  scg5d1_hd U401 ( .A(N217), .B(n228), .C(n154), .D(n242), .E(n368), .F(N216), 
        .Y(N211) );
  scg5d1_hd U402 ( .A(N217), .B(n227), .C(n154), .D(n243), .E(n369), .F(N216), 
        .Y(N210) );
  scg5d1_hd U403 ( .A(N217), .B(n226), .C(n154), .D(n244), .E(n370), .F(N216), 
        .Y(N209) );
  scg5d1_hd U404 ( .A(N217), .B(n225), .C(n154), .D(n245), .E(n371), .F(N216), 
        .Y(N208) );
  scg5d1_hd U405 ( .A(N217), .B(n224), .C(n154), .D(n246), .E(n372), .F(N216), 
        .Y(N207) );
  scg5d1_hd U406 ( .A(N217), .B(n223), .C(n154), .D(n247), .E(n373), .F(N216), 
        .Y(N206) );
  scg5d1_hd U407 ( .A(N217), .B(n290), .C(n154), .D(n248), .E(n448), .F(N216), 
        .Y(N205) );
  scg5d1_hd U408 ( .A(N217), .B(n291), .C(n154), .D(n249), .E(n449), .F(N216), 
        .Y(N204) );
  scg5d1_hd U409 ( .A(N217), .B(n292), .C(n154), .D(n250), .E(n450), .F(N216), 
        .Y(N203) );
  scg5d1_hd U410 ( .A(N217), .B(n293), .C(n154), .D(n251), .E(n451), .F(N216), 
        .Y(N202) );
  scg5d1_hd U411 ( .A(N217), .B(n294), .C(n154), .D(n252), .E(n452), .F(N216), 
        .Y(N201) );
  scg5d1_hd U412 ( .A(N217), .B(n295), .C(n154), .D(n253), .E(n453), .F(N216), 
        .Y(N200) );
  scg5d1_hd U413 ( .A(N217), .B(n296), .C(n154), .D(n254), .E(n454), .F(N216), 
        .Y(N199) );
  scg5d1_hd U414 ( .A(N217), .B(n297), .C(n154), .D(n255), .E(n455), .F(N216), 
        .Y(N198) );
  ad2d1_hd U415 ( .A(n154), .B(n256), .Y(N197) );
  ad2d1_hd U416 ( .A(n154), .B(n257), .Y(N196) );
  ad2d1_hd U417 ( .A(n154), .B(n258), .Y(N195) );
  ad2d1_hd U418 ( .A(n154), .B(n259), .Y(N194) );
  ad2d1_hd U419 ( .A(n154), .B(n260), .Y(N193) );
  ad2d1_hd U420 ( .A(n154), .B(n261), .Y(N192) );
  ad2d1_hd U421 ( .A(n154), .B(n262), .Y(N191) );
  ad2d1_hd U422 ( .A(n154), .B(n263), .Y(N190) );
  ad2d1_hd U423 ( .A(n154), .B(n412), .Y(N185) );
  ad2d1_hd U424 ( .A(n154), .B(n413), .Y(N184) );
  ad2d1_hd U425 ( .A(n154), .B(n414), .Y(N183) );
  ad2d1_hd U426 ( .A(n154), .B(n415), .Y(N182) );
  ad2d1_hd U427 ( .A(n154), .B(n416), .Y(N181) );
  ad2d1_hd U428 ( .A(n154), .B(n417), .Y(N180) );
  ad2d1_hd U429 ( .A(n154), .B(n418), .Y(N179) );
  ad2d1_hd U430 ( .A(n154), .B(n419), .Y(N178) );
  ad2d1_hd U431 ( .A(n154), .B(n420), .Y(N177) );
  ad2d1_hd U432 ( .A(n154), .B(n421), .Y(N176) );
  ad2d1_hd U433 ( .A(n154), .B(n422), .Y(N175) );
  ad2d1_hd U434 ( .A(n154), .B(n423), .Y(N174) );
  ad2d1_hd U435 ( .A(N166), .B(n538), .Y(N170) );
  ad2d1_hd U436 ( .A(N165), .B(n538), .Y(N169) );
  ad2d1_hd U437 ( .A(N164), .B(n538), .Y(N168) );
  nr2bd1_hd U438 ( .AN(n538), .B(n352), .Y(N167) );
  nd4d1_hd U442 ( .A(n61), .B(N1111), .C(N1079), .D(n196), .Y(n195) );
  nr4d1_hd U443 ( .A(n517), .B(n551), .C(n45), .D(n60), .Y(n196) );
  scg18d1_hd U446 ( .A(N768), .B(i_ADS1292_BUSY), .C(N1282), .D(n198), .E(n44), 
        .Y(n197) );
  ao21d1_hd U449 ( .A(n491), .B(N803), .C(N1027), .Y(n200) );
  ao21d1_hd U450 ( .A(N915), .B(N768), .C(N1278), .Y(n199) );
  ivd1_hd U453 ( .A(n542), .Y(n203) );
  nd3d1_hd U454 ( .A(n204), .B(n205), .C(n206), .Y(N1022) );
  nd2bd1_hd U466 ( .AN(i_ADS1292_BUSY), .B(n527), .Y(n206) );
  nd2bd1_hd U468 ( .AN(n535), .B(n205), .Y(N1013) );
  nr2d1_hd U471 ( .A(n202), .B(n63), .Y(N1006) );
  nr2d1_hd U473 ( .A(n202), .B(n64), .Y(N1005) );
  ivd1_hd U475 ( .A(n491), .Y(n202) );
  ad2d1_hd U476 ( .A(N810), .B(n491), .Y(N1004) );
  nr2d1_hd U477 ( .A(n66), .B(n158), .Y(N810) );
  ad2d1_hd U478 ( .A(N809), .B(n491), .Y(N1003) );
  nr2d1_hd U479 ( .A(n159), .B(n66), .Y(N809) );
  scg7d1_hd U480 ( .A(n491), .B(N808), .C(N751), .D(n208), .E(n36), .Y(N1002)
         );
  oa21d1_hd U481 ( .A(n58), .B(n49), .C(N1111), .Y(n208) );
  nr2d1_hd U483 ( .A(N1172), .B(n54), .Y(n61) );
  ivd1_hd U485 ( .A(n517), .Y(n48) );
  nr2d1_hd U486 ( .A(n66), .B(n160), .Y(N808) );
  ao22d1_hd U489 ( .A(N807), .B(n491), .C(n52), .D(n54), .Y(n210) );
  ivd1_hd U490 ( .A(n55), .Y(n52) );
  nr2d1_hd U492 ( .A(n161), .B(n66), .Y(N807) );
  scg17d1_hd U493 ( .A(n491), .B(N806), .C(n36), .D(n211), .Y(N1000) );
  oa21d1_hd U494 ( .A(n212), .B(n45), .C(n39), .Y(n211) );
  ad2d1_hd U495 ( .A(N1111), .B(N751), .Y(n39) );
  ivd1_hd U496 ( .A(n209), .Y(n45) );
  nr2d1_hd U497 ( .A(n541), .B(n523), .Y(n209) );
  ao21d1_hd U498 ( .A(n42), .B(N1171), .C(n54), .Y(n212) );
  ao21d1_hd U503 ( .A(N1187), .B(n213), .C(n517), .Y(n42) );
  ivd1_hd U504 ( .A(N1195), .Y(n213) );
  nr2d1_hd U505 ( .A(N1079), .B(n193), .Y(n36) );
  nr2d1_hd U506 ( .A(n162), .B(n66), .Y(N806) );
  ivd1_hd U507 ( .A(N804), .Y(n66) );
  nr2d1_hd U771 ( .A(N773), .B(N774), .Y(n527) );
  nid1_hd U772 ( .A(n543), .Y(N8) );
  nd2d1_hd U774 ( .A(n95), .B(n73), .Y(N717) );
  ad2d1_hd U791 ( .A(N444), .B(N343), .Y(N472) );
  or2d1_hd U792 ( .A(n460), .B(N343), .Y(N426) );
  or2d1_hd U793 ( .A(n340), .B(n339), .Y(N1213) );
  ivd1_hd U794 ( .A(n406), .Y(gt_x_149_n15) );
  ivd1_hd U795 ( .A(n232), .Y(N1113) );
  or2d1_hd U796 ( .A(N470), .B(N1311), .Y(N1312) );
  ad2d1_hd U797 ( .A(N343), .B(n92), .Y(N470) );
  or2d1_hd U798 ( .A(N471), .B(N472), .Y(N1311) );
  ad2d1_hd U799 ( .A(n460), .B(n67), .Y(N471) );
  ivd1_hd U800 ( .A(n393), .Y(gt_x_61_n15) );
  or2d1_hd U801 ( .A(N429), .B(N428), .Y(N430) );
  or2d1_hd U802 ( .A(N426), .B(N427), .Y(N429) );
  or2d1_hd U803 ( .A(N395), .B(N370), .Y(N427) );
  ivd1_hd U804 ( .A(n355), .Y(N1317) );
  or2d1_hd U805 ( .A(n460), .B(N343), .Y(N396) );
  or2d1_hd U806 ( .A(n232), .B(N1097), .Y(N1098) );
  or2d1_hd U807 ( .A(N1039), .B(N1096), .Y(N1097) );
  or2d1_hd U808 ( .A(N1038), .B(n231), .Y(N1096) );
  ivd1_hd U809 ( .A(n233), .Y(N1094) );
  or2d1_hd U810 ( .A(n232), .B(N1042), .Y(N1043) );
  or2d1_hd U811 ( .A(N1039), .B(N1041), .Y(N1042) );
  or2d1_hd U812 ( .A(N1038), .B(n231), .Y(N1041) );
  or2d1_hd U814 ( .A(n460), .B(N343), .Y(N358) );
  or2d1_hd U815 ( .A(N1069), .B(n339), .Y(N1181) );
  or2d1_hd U816 ( .A(N1069), .B(n339), .Y(N1189) );
  clknd2d1_hd U817 ( .A(n112), .B(n106), .Y(n155) );
  or2d1_hd U818 ( .A(n340), .B(n339), .Y(N1209) );
  or2d1_hd U819 ( .A(n460), .B(N343), .Y(N420) );
  or2d1_hd U820 ( .A(n340), .B(N1068), .Y(N1157) );
  or2d1_hd U821 ( .A(N1131), .B(N1165), .Y(N1166) );
  or2d1_hd U822 ( .A(N1069), .B(n339), .Y(N1165) );
  clknd2d1_hd U823 ( .A(N1207), .B(N1211), .Y(n121) );
  ivd1_hd U824 ( .A(n408), .Y(N1070) );
  or2d1_hd U825 ( .A(n460), .B(N343), .Y(N351) );
  or2d1_hd U826 ( .A(N1069), .B(N1068), .Y(N1071) );
  nr2d1_hd U827 ( .A(n97), .B(N1303), .Y(n71) );
  or2d1_hd U828 ( .A(n460), .B(N343), .Y(N402) );
  or2d1_hd U829 ( .A(N765), .B(N766), .Y(N767) );
  nr2d1_hd U830 ( .A(gt_x_149_n15), .B(gt_x_149_n18), .Y(gt_x_149_n14) );
  ivd1_hd U831 ( .A(n407), .Y(gt_x_149_n18) );
  ivd1_hd U832 ( .A(n460), .Y(N444) );
  or2d1_hd U833 ( .A(N444), .B(n67), .Y(N445) );
  or2d1_hd U834 ( .A(n460), .B(N343), .Y(N371) );
  or2d1_hd U835 ( .A(N1113), .B(N1124), .Y(N1125) );
  or2d1_hd U836 ( .A(n345), .B(N1123), .Y(N1124) );
  or2d1_hd U837 ( .A(N1038), .B(n231), .Y(N1123) );
  or2d1_hd U838 ( .A(N1113), .B(N1116), .Y(N1117) );
  or2d1_hd U839 ( .A(n345), .B(N1115), .Y(N1116) );
  or2d1_hd U840 ( .A(N1038), .B(n231), .Y(N1115) );
  ivd1_hd U841 ( .A(n235), .Y(N1114) );
  ivd1_hd U842 ( .A(n347), .Y(N274) );
  ivd1_hd U843 ( .A(n78), .Y(N275) );
  or2d1_hd U844 ( .A(n460), .B(N343), .Y(N364) );
  or2d1_hd U845 ( .A(n342), .B(N1161), .Y(N1162) );
  or2d1_hd U846 ( .A(N1144), .B(n341), .Y(N1161) );
  or2d1_hd U847 ( .A(N1076), .B(N1185), .Y(N1186) );
  or2d1_hd U848 ( .A(n342), .B(N1201), .Y(N1202) );
  clknd2d1_hd U849 ( .A(n531), .B(n96), .Y(n94) );
  or2d1_hd U850 ( .A(n460), .B(N343), .Y(N438) );
  or2d1_hd U851 ( .A(n460), .B(N343), .Y(N377) );
  ivd2_hd U852 ( .A(n67), .Y(N343) );
  or2d1_hd U853 ( .A(N468), .B(N1313), .Y(N1314) );
  ad2d1_hd U854 ( .A(N343), .B(n459), .Y(N468) );
  or2d1_hd U855 ( .A(N469), .B(N1312), .Y(N1313) );
  ad2d1_hd U856 ( .A(n460), .B(n92), .Y(N469) );
  ad2d1_hd U857 ( .A(n460), .B(n459), .Y(N467) );
  clknd2d1_hd U858 ( .A(n531), .B(i_MPR121_BUSY), .Y(n84) );
  or2d1_hd U859 ( .A(n460), .B(N343), .Y(N389) );
  or2d1_hd U860 ( .A(n460), .B(N343), .Y(N414) );
  or2d1_hd U861 ( .A(n460), .B(N343), .Y(N408) );
  or2d1_hd U862 ( .A(n460), .B(N343), .Y(N344) );
  ivd1_hd U863 ( .A(N475), .Y(alt36_n129) );
  nr2d1_hd U864 ( .A(gt_x_61_n15), .B(gt_x_61_n18), .Y(gt_x_61_n14) );
  ivd1_hd U865 ( .A(n394), .Y(gt_x_61_n18) );
  or2d1_hd U866 ( .A(n460), .B(N343), .Y(N383) );
  or2d1_hd U867 ( .A(N444), .B(n67), .Y(N451) );
  ivd1_hd U868 ( .A(n459), .Y(N370) );
  or2d1_hd U869 ( .A(n460), .B(N343), .Y(N432) );
  ivd1_hd U870 ( .A(n92), .Y(N395) );
  clknd2d1_hd U871 ( .A(n519), .B(n556), .Y(n70) );
  clknd2d1_hd U872 ( .A(n7), .B(n6), .Y(n14) );
  ivd1_hd U873 ( .A(N796), .Y(alt36_n513) );
  or2d1_hd U874 ( .A(N741), .B(N742), .Y(N778) );
  ivd1_hd U875 ( .A(n238), .Y(N742) );
  ad2d1_hd U876 ( .A(i_ADS1292_FILTERED_DATA_VALID), .B(alt36_n508), .Y(N933)
         );
  ad2d1_hd U877 ( .A(n395), .B(N303), .Y(N797) );
  ad2d1_hd U878 ( .A(n349), .B(N298), .Y(N796) );
  ad2d1_hd U880 ( .A(n426), .B(n10), .Y(N798) );
  ad2d1_hd U881 ( .A(N1319), .B(n365), .Y(N929) );
  ivd1_hd U884 ( .A(n239), .Y(N764) );
  ad2d1_hd U885 ( .A(N793), .B(N742), .Y(N794) );
  ad2d1_hd U886 ( .A(N764), .B(N747), .Y(N793) );
  or2d1_hd U887 ( .A(i_ADS1292_BUSY), .B(N915), .Y(N914) );
  clknd2d1_hd U888 ( .A(n542), .B(N932), .Y(n198) );
  or2d1_hd U889 ( .A(N933), .B(n540), .Y(N932) );
  or2d1_hd U890 ( .A(N764), .B(N747), .Y(N785) );
  ad2d1_hd U891 ( .A(n355), .B(N302), .Y(N475) );
  or2d1_hd U893 ( .A(i_MPR121_BUSY), .B(N608), .Y(N626) );
  or2d1_hd U894 ( .A(N396), .B(N397), .Y(N399) );
  or2d1_hd U895 ( .A(N395), .B(n459), .Y(N397) );
  or2d1_hd U897 ( .A(n343), .B(N1064), .Y(N1065) );
  or2d1_hd U898 ( .A(N1049), .B(n435), .Y(N1064) );
  or2d1_hd U899 ( .A(N741), .B(n238), .Y(N774) );
  or2d1_hd U901 ( .A(n235), .B(N1100), .Y(N1101) );
  or2d1_hd U902 ( .A(N1095), .B(N1099), .Y(N1100) );
  ivd1_hd U903 ( .A(n234), .Y(N1095) );
  or2d1_hd U904 ( .A(N1094), .B(N1098), .Y(N1099) );
  clknd2d1_hd U905 ( .A(alt36_n329), .B(n270), .Y(n9) );
  ad2d1_hd U906 ( .A(alt36_n332), .B(n10), .Y(alt36_n329) );
  or2d1_hd U907 ( .A(n235), .B(N1045), .Y(N1046) );
  or2d1_hd U908 ( .A(n234), .B(N1044), .Y(N1045) );
  or2d1_hd U909 ( .A(n233), .B(N1043), .Y(N1044) );
  clknd2d1_hd U910 ( .A(N250), .B(i_UART_DATA_TX_READY), .Y(n185) );
  ad2d1_hd U911 ( .A(n566), .B(alt36_n509), .Y(N915) );
  ivd1_hd U912 ( .A(i_ADS1292_BUSY), .Y(alt36_n509) );
  or2d1_hd U913 ( .A(n467), .B(N1087), .Y(N1088) );
  or2d1_hd U914 ( .A(N796), .B(N1032), .Y(N803) );
  or2d1_hd U915 ( .A(N1131), .B(N1197), .Y(N1198) );
  or2d1_hd U916 ( .A(n340), .B(n339), .Y(N1197) );
  or2d1_hd U917 ( .A(N1131), .B(N1205), .Y(N1206) );
  or2d1_hd U918 ( .A(n340), .B(n339), .Y(N1205) );
  clknd2d1_hd U919 ( .A(N1175), .B(N1183), .Y(n123) );
  or2d1_hd U920 ( .A(N361), .B(N360), .Y(N362) );
  or2d1_hd U921 ( .A(N358), .B(N359), .Y(N361) );
  or2d1_hd U922 ( .A(n92), .B(n459), .Y(N359) );
  or2d1_hd U923 ( .A(N1131), .B(N1173), .Y(N1174) );
  or2d1_hd U924 ( .A(N1069), .B(n339), .Y(N1173) );
  clknd2d1_hd U925 ( .A(n109), .B(n152), .Y(n149) );
  nr2d1_hd U926 ( .A(i_UART_DATA_RX_VALID), .B(n191), .Y(N250) );
  or2d1_hd U927 ( .A(N1069), .B(N1068), .Y(N1104) );
  or2d1_hd U928 ( .A(N420), .B(N421), .Y(N423) );
  or2d1_hd U929 ( .A(N395), .B(N370), .Y(N421) );
  clknd2d1_hd U930 ( .A(N1167), .B(N1159), .Y(n119) );
  or2d1_hd U931 ( .A(n340), .B(N1068), .Y(N1149) );
  or2d1_hd U932 ( .A(N1131), .B(N1140), .Y(N1141) );
  or2d1_hd U933 ( .A(n340), .B(N1068), .Y(N1140) );
  or2d1_hd U934 ( .A(N1131), .B(N1132), .Y(N1133) );
  or2d1_hd U935 ( .A(n340), .B(N1068), .Y(N1132) );
  clknd2d1_hd U936 ( .A(n111), .B(n101), .Y(n120) );
  or2d1_hd U937 ( .A(N354), .B(N353), .Y(N355) );
  or2d1_hd U938 ( .A(N351), .B(N352), .Y(N354) );
  or2d1_hd U939 ( .A(n92), .B(n459), .Y(N352) );
  clknd2d1_hd U940 ( .A(N1073), .B(n109), .Y(n100) );
  ivd1_hd U941 ( .A(n526), .Y(n95) );
  clknd2d1_hd U942 ( .A(n70), .B(n71), .Y(N725) );
  ad2d1_hd U943 ( .A(n180), .B(alt36_n288), .Y(alt36_n287) );
  ivd1_hd U944 ( .A(n446), .Y(alt36_n288) );
  or2d1_hd U945 ( .A(N402), .B(N403), .Y(N405) );
  or2d1_hd U946 ( .A(N395), .B(n459), .Y(N403) );
  or2d1_hd U947 ( .A(N1243), .B(N1244), .Y(N709) );
  clknd2d1_hd U948 ( .A(n16), .B(n21), .Y(N1243) );
  clknd2d1_hd U949 ( .A(N481), .B(n237), .Y(n103) );
  clknd2d1_hd U950 ( .A(N481), .B(n236), .Y(n102) );
  nid1_hd U951 ( .A(n547), .Y(N68) );
  or2d1_hd U952 ( .A(N1238), .B(N1239), .Y(N1020) );
  or2d1_hd U953 ( .A(n546), .B(n527), .Y(N1239) );
  clknd2d1_hd U954 ( .A(n23), .B(N767), .Y(N1238) );
  clknd2d1_hd U955 ( .A(N63), .B(N603), .Y(n99) );
  clknd2d1_hd U956 ( .A(n530), .B(n554), .Y(n44) );
  or2d1_hd U957 ( .A(n491), .B(n530), .Y(N1019) );
  or2d1_hd U958 ( .A(n513), .B(n546), .Y(N1030) );
  or2d1_hd U959 ( .A(n92), .B(n459), .Y(N458) );
  or2d1_hd U960 ( .A(N444), .B(n67), .Y(N457) );
  clknd2d1_hd U961 ( .A(n93), .B(N68), .Y(n85) );
  or2d1_hd U962 ( .A(N445), .B(N446), .Y(N448) );
  or2d1_hd U963 ( .A(n92), .B(n459), .Y(N446) );
  or2d1_hd U964 ( .A(n526), .B(n512), .Y(N718) );
  or3d1_hd U965 ( .A(n553), .B(n514), .C(N431), .Y(N728) );
  nr2ad1_hd U966 ( .A(N760), .B(N761), .Y(n513) );
  or2d1_hd U967 ( .A(n239), .B(N747), .Y(N760) );
  or2d1_hd U968 ( .A(N741), .B(N742), .Y(N761) );
  or2d1_hd U969 ( .A(n239), .B(N747), .Y(N752) );
  or2d1_hd U970 ( .A(n239), .B(N747), .Y(N756) );
  or2d1_hd U971 ( .A(N741), .B(n238), .Y(N757) );
  nr2ad1_hd U972 ( .A(N374), .B(N373), .Y(n553) );
  or2d1_hd U973 ( .A(N371), .B(N372), .Y(N374) );
  or2d1_hd U974 ( .A(n92), .B(N370), .Y(N372) );
  or2d1_hd U975 ( .A(N1050), .B(N1055), .Y(N1056) );
  or2d1_hd U976 ( .A(N1049), .B(n435), .Y(N1055) );
  or2d1_hd U977 ( .A(N1114), .B(N1127), .Y(N1128) );
  or2d1_hd U978 ( .A(n234), .B(N1126), .Y(N1127) );
  or2d1_hd U979 ( .A(n233), .B(N1125), .Y(N1126) );
  or2d1_hd U980 ( .A(N1114), .B(N1119), .Y(N1120) );
  or2d1_hd U981 ( .A(n234), .B(N1118), .Y(N1119) );
  or2d1_hd U982 ( .A(n233), .B(N1117), .Y(N1118) );
  or2d1_hd U983 ( .A(n445), .B(alt36_n301), .Y(alt36_n298) );
  or2d1_hd U984 ( .A(n446), .B(n356), .Y(alt36_n301) );
  oa21d1_hd U985 ( .A(n462), .B(N283), .C(n911), .Y(N330) );
  or2d1_hd U986 ( .A(n347), .B(N275), .Y(N285) );
  or2d1_hd U987 ( .A(N274), .B(n78), .Y(N288) );
  ad2d1_hd U988 ( .A(N274), .B(N275), .Y(N277) );
  or2d1_hd U989 ( .A(n347), .B(n78), .Y(N279) );
  or2d1_hd U990 ( .A(N282), .B(n461), .Y(N283) );
  or2d1_hd U991 ( .A(n347), .B(N275), .Y(N282) );
  ad2d1_hd U992 ( .A(n351), .B(N1091), .Y(N1092) );
  ad2d1_hd U993 ( .A(n353), .B(n350), .Y(N1091) );
  ivd1_hd U994 ( .A(N250), .Y(n184) );
  ivd1_hd U995 ( .A(N8), .Y(n191) );
  or2d1_hd U996 ( .A(N364), .B(N365), .Y(N367) );
  or2d1_hd U997 ( .A(N357), .B(N350), .Y(N366) );
  or2d1_hd U998 ( .A(n92), .B(n459), .Y(N365) );
  or2d1_hd U999 ( .A(n526), .B(N63), .Y(N711) );
  or2d1_hd U1000 ( .A(n491), .B(N751), .Y(N1016) );
  or2d1_hd U1001 ( .A(N1076), .B(N1077), .Y(N1078) );
  or2d1_hd U1002 ( .A(N1076), .B(N1177), .Y(N1178) );
  clknd2d1_hd U1003 ( .A(N1195), .B(N1187), .Y(n60) );
  or2d1_hd U1004 ( .A(n342), .B(N1193), .Y(N1194) );
  clknd2d1_hd U1005 ( .A(N1079), .B(n39), .Y(n55) );
  clknd2d1_hd U1006 ( .A(n61), .B(n52), .Y(n46) );
  or2d1_hd U1007 ( .A(N1076), .B(N1145), .Y(N1146) );
  or2d1_hd U1008 ( .A(N1144), .B(n341), .Y(N1145) );
  or2d1_hd U1009 ( .A(N1076), .B(N1153), .Y(N1154) );
  or2d1_hd U1010 ( .A(N1144), .B(n341), .Y(N1153) );
  or2d1_hd U1011 ( .A(n342), .B(N1136), .Y(N1137) );
  or2d1_hd U1012 ( .A(n337), .B(N1170), .Y(N1171) );
  or2d1_hd U1013 ( .A(n342), .B(N1169), .Y(N1170) );
  or2d1_hd U1014 ( .A(N1144), .B(n341), .Y(N1169) );
  clknd2d1_hd U1015 ( .A(N1163), .B(N1155), .Y(n54) );
  clknd2d1_hd U1016 ( .A(n45), .B(n52), .Y(n56) );
  or2d1_hd U1017 ( .A(n239), .B(N747), .Y(N748) );
  clknd2d1_hd U1018 ( .A(n61), .B(n209), .Y(n49) );
  clknd2d1_hd U1019 ( .A(N1187), .B(n48), .Y(n58) );
  or2d1_hd U1020 ( .A(n342), .B(N1109), .Y(N1110) );
  clknd2d1_hd U1021 ( .A(N804), .B(n237), .Y(n64) );
  clknd2d1_hd U1022 ( .A(N804), .B(n236), .Y(n63) );
  ad2d1_hd U1024 ( .A(i_MPR121_FAIL), .B(alt36_n127), .Y(N608) );
  ivd1_hd U1025 ( .A(i_MPR121_BUSY), .Y(alt36_n127) );
  or2d1_hd U1026 ( .A(N438), .B(N439), .Y(N441) );
  or2d1_hd U1027 ( .A(N357), .B(N350), .Y(N440) );
  or2d1_hd U1028 ( .A(N395), .B(N370), .Y(N439) );
  clknd2d1_hd U1029 ( .A(n392), .B(N68), .Y(n73) );
  or2d1_hd U1030 ( .A(N377), .B(N378), .Y(N380) );
  or2d1_hd U1031 ( .A(n92), .B(N370), .Y(N378) );
  or2d1_hd U1032 ( .A(N466), .B(N1315), .Y(N1316) );
  or2d1_hd U1033 ( .A(N467), .B(N1314), .Y(N1315) );
  clknd2d1_hd U1034 ( .A(n84), .B(n85), .Y(n76) );
  or2d1_hd U1035 ( .A(N389), .B(N390), .Y(N392) );
  or2d1_hd U1036 ( .A(N357), .B(N350), .Y(N391) );
  or2d1_hd U1037 ( .A(n92), .B(N370), .Y(N390) );
  or2d1_hd U1038 ( .A(N414), .B(N415), .Y(N417) );
  or2d1_hd U1039 ( .A(N357), .B(N350), .Y(N416) );
  or2d1_hd U1040 ( .A(N395), .B(n459), .Y(N415) );
  or2d1_hd U1041 ( .A(N408), .B(N409), .Y(N411) );
  or2d1_hd U1042 ( .A(N395), .B(n459), .Y(N409) );
  nr2ad1_hd U1043 ( .A(N347), .B(N346), .Y(n526) );
  or2d1_hd U1044 ( .A(N344), .B(N345), .Y(N347) );
  or2d1_hd U1045 ( .A(n92), .B(n459), .Y(N345) );
  ad2d1_hd U1046 ( .A(N476), .B(alt36_n128), .Y(N481) );
  ad2d1_hd U1047 ( .A(n354), .B(N304), .Y(N476) );
  ad2d1_hd U1048 ( .A(n555), .B(alt36_n129), .Y(alt36_n128) );
  ivd1_hd U1049 ( .A(n270), .Y(N304) );
  clknd2d1_hd U1050 ( .A(n520), .B(n512), .Y(n80) );
  or2d1_hd U1051 ( .A(N383), .B(N384), .Y(N386) );
  or2d1_hd U1052 ( .A(n92), .B(N370), .Y(N384) );
  or2d1_hd U1053 ( .A(N451), .B(N452), .Y(N454) );
  or2d1_hd U1054 ( .A(n92), .B(n459), .Y(N452) );
  or2d1_hd U1055 ( .A(N432), .B(N433), .Y(N435) );
  or2d1_hd U1056 ( .A(N395), .B(N370), .Y(N433) );
  or2d1_hd U1057 ( .A(i_MPR121_BUSY), .B(n96), .Y(N607) );
  or2d1_hd U1058 ( .A(N764), .B(N747), .Y(N781) );
  ivd1_hd U1059 ( .A(alt36_n60), .Y(N802) );
  ad2d1_hd U1060 ( .A(N797), .B(alt36_n513), .Y(N1032) );
  ad2d1_hd U1061 ( .A(N798), .B(alt36_n510), .Y(N804) );
  ad2d1_hd U1062 ( .A(alt36_n513), .B(alt36_n511), .Y(alt36_n510) );
  ivd1_hd U1063 ( .A(N797), .Y(alt36_n511) );
  or2d1_hd U1064 ( .A(N741), .B(N742), .Y(N744) );
  clknd2d1_hd U1065 ( .A(n542), .B(N933), .Y(n205) );
  ivd1_hd U1066 ( .A(n62), .Y(N1027) );
  or2d1_hd U1067 ( .A(N798), .B(alt36_n63), .Y(alt36_n60) );
  or2d1_hd U1068 ( .A(N797), .B(N796), .Y(alt36_n63) );
  ivd1_hd U1069 ( .A(N929), .Y(alt36_n508) );
  or2d1_hd U1070 ( .A(N790), .B(N1318), .Y(N795) );
  ad2d1_hd U1071 ( .A(N789), .B(N741), .Y(N790) );
  or2d1_hd U1072 ( .A(N792), .B(N794), .Y(N1318) );
  ad2d1_hd U1073 ( .A(N764), .B(N747), .Y(N789) );
  clknd2d1_hd U1074 ( .A(n550), .B(n569), .Y(N1021) );
  clknd2d1_hd U1075 ( .A(N768), .B(N914), .Y(n569) );
  clknd2d1_hd U1076 ( .A(n23), .B(n193), .Y(N1240) );
  clknd2d1_hd U1077 ( .A(n198), .B(n552), .Y(N1018) );
  mx2d1_hd U1078 ( .D0(o_ADS1292_FILTERED_DATA_ACK), .D1(n542), .S(N1013), .Y(
        n619) );
  clknd2d1_hd U1079 ( .A(n572), .B(n573), .Y(r_mpr_pstate[1]) );
  ivd1_hd U1080 ( .A(n86), .Y(n572) );
  ad2d1_hd U1081 ( .A(N475), .B(n555), .Y(N480) );
  clknd2d1_hd U1082 ( .A(n88), .B(n89), .Y(r_mpr_pstate[0]) );
  clknd2d1_hd U1093 ( .A(n188), .B(n559), .Y(n190) );
  clknd2d1_hd U1095 ( .A(n188), .B(n560), .Y(n187) );
  clknd2d1_hd U1096 ( .A(n199), .B(n200), .Y(N1024) );
  mx2d1_hd U1097 ( .D0(n444), .D1(N640), .S(N712), .Y(r_mpr_second_param[0])
         );
  mx2d1_hd U1098 ( .D0(n443), .D1(N641), .S(N712), .Y(r_mpr_second_param[1])
         );
  mx2d1_hd U1099 ( .D0(n442), .D1(N642), .S(N712), .Y(r_mpr_second_param[2])
         );
  clknd2d1_hd U1100 ( .A(n150), .B(n151), .Y(N642) );
  mx2d1_hd U1101 ( .D0(n441), .D1(N643), .S(N712), .Y(r_mpr_second_param[3])
         );
  mx2d1_hd U1102 ( .D0(n440), .D1(N644), .S(N712), .Y(r_mpr_second_param[4])
         );
  mx2d1_hd U1103 ( .D0(n439), .D1(N645), .S(N712), .Y(r_mpr_second_param[6])
         );
  mx2d1_hd U1104 ( .D0(n438), .D1(N363), .S(N712), .Y(r_mpr_second_param[7])
         );
  or2d1_hd U1107 ( .A(N63), .B(n544), .Y(N700) );
  mx2d1_hd U1108 ( .D0(n435), .D1(N703), .S(n524), .Y(N1052) );
  or2d1_hd U1109 ( .A(n547), .B(N462), .Y(N703) );
  mx2d1_hd U1110 ( .D0(n434), .D1(N691), .S(N725), .Y(r_mpr_first_param[0]) );
  mx2d1_hd U1111 ( .D0(n433), .D1(N692), .S(N725), .Y(r_mpr_first_param[1]) );
  mx2d1_hd U1112 ( .D0(n432), .D1(N693), .S(N725), .Y(r_mpr_first_param[2]) );
  clknd2d1_hd U1113 ( .A(n526), .B(N484), .Y(n115) );
  mx2d1_hd U1114 ( .D0(n431), .D1(N694), .S(N725), .Y(r_mpr_first_param[3]) );
  mx2d1_hd U1115 ( .D0(n430), .D1(N695), .S(N725), .Y(r_mpr_first_param[4]) );
  clknd2d1_hd U1116 ( .A(n107), .B(n108), .Y(N695) );
  mx2d1_hd U1117 ( .D0(n429), .D1(N696), .S(N725), .Y(r_mpr_first_param[5]) );
  scg2d1_hd U1118 ( .A(n526), .B(N487), .C(n105), .D(n106), .Y(N696) );
  mx2d1_hd U1119 ( .D0(n428), .D1(N697), .S(N725), .Y(r_mpr_first_param[6]) );
  mx2d1_hd U1120 ( .D0(n427), .D1(N698), .S(N725), .Y(r_mpr_first_param[7]) );
  mx2d1_hd U1121 ( .D0(n426), .D1(N322), .S(N326), .Y(r_ads_read_reg) );
  ad2d1_hd U1122 ( .A(n445), .B(alt36_n287), .Y(N309) );
  mx2d1_hd U1123 ( .D0(o_MPR121_WRITE_ENABLE), .D1(n534), .S(N709), .Y(n597)
         );
  mx2d1_hd U1124 ( .D0(o_MPR121_READ_ENABLE), .D1(N631), .S(N709), .Y(n598) );
  or2d1_hd U1125 ( .A(n548), .B(n532), .Y(N631) );
  mx2d1_hd U1126 ( .D0(n423), .D1(N667), .S(N717), .Y(r_mpr_touch_status[0])
         );
  mx2d1_hd U1127 ( .D0(n422), .D1(N668), .S(N717), .Y(r_mpr_touch_status[1])
         );
  mx2d1_hd U1128 ( .D0(n421), .D1(N669), .S(N717), .Y(r_mpr_touch_status[2])
         );
  mx2d1_hd U1129 ( .D0(n420), .D1(N670), .S(N717), .Y(r_mpr_touch_status[3])
         );
  mx2d1_hd U1130 ( .D0(n419), .D1(N671), .S(N717), .Y(r_mpr_touch_status[4])
         );
  mx2d1_hd U1131 ( .D0(n418), .D1(N672), .S(N717), .Y(r_mpr_touch_status[5])
         );
  mx2d1_hd U1132 ( .D0(n417), .D1(N673), .S(N717), .Y(r_mpr_touch_status[6])
         );
  mx2d1_hd U1133 ( .D0(n416), .D1(N674), .S(N717), .Y(r_mpr_touch_status[7])
         );
  mx2d1_hd U1134 ( .D0(n415), .D1(N675), .S(N717), .Y(r_mpr_touch_status[8])
         );
  mx2d1_hd U1135 ( .D0(n414), .D1(N676), .S(N717), .Y(r_mpr_touch_status[9])
         );
  mx2d1_hd U1136 ( .D0(n413), .D1(N677), .S(N717), .Y(r_mpr_touch_status[10])
         );
  mx2d1_hd U1137 ( .D0(n412), .D1(N678), .S(N717), .Y(r_mpr_touch_status[11])
         );
  mx2d1_hd U1138 ( .D0(o_ADS1292_CONTROL[0]), .D1(N990), .S(N1020), .Y(n602)
         );
  clknd2d1_hd U1139 ( .A(n4), .B(n6), .Y(N990) );
  mx2d1_hd U1140 ( .D0(o_ADS1292_CONTROL[1]), .D1(N991), .S(N1020), .Y(n601)
         );
  mx2d1_hd U1141 ( .D0(o_ADS1292_CONTROL[2]), .D1(N992), .S(N1020), .Y(n600)
         );
  mx2d1_hd U1142 ( .D0(n408), .D1(N635), .S(N711), .Y(r_mpr_set_counter[0]) );
  mx2d1_hd U1143 ( .D0(n407), .D1(N986), .S(N1019), .Y(gt_x_149_n17) );
  mx2d1_hd U1144 ( .D0(n406), .D1(N987), .S(N1019), .Y(r_ads_clk_counter[2])
         );
  mx2d1_hd U1145 ( .D0(n405), .D1(N988), .S(N1019), .Y(gt_x_149_n9) );
  xo2d1_hd U1146 ( .A(add_x_150_n1), .B(n405), .Y(N923) );
  mx2d1_hd U1147 ( .D0(n404), .D1(N985), .S(N1019), .Y(r_ads_clk_counter[0])
         );
  mx2d1_hd U1148 ( .D0(o_ADS1292_REG_ADDR[0]), .D1(n317), .S(N1030), .Y(n610)
         );
  mx2d1_hd U1149 ( .D0(o_ADS1292_REG_ADDR[1]), .D1(n316), .S(N1030), .Y(n609)
         );
  mx2d1_hd U1150 ( .D0(o_ADS1292_REG_ADDR[2]), .D1(n315), .S(N1030), .Y(n608)
         );
  mx2d1_hd U1151 ( .D0(o_ADS1292_REG_ADDR[3]), .D1(n314), .S(N1030), .Y(n607)
         );
  mx2d1_hd U1152 ( .D0(o_ADS1292_REG_ADDR[4]), .D1(n313), .S(N1030), .Y(n606)
         );
  mx2d1_hd U1153 ( .D0(o_ADS1292_REG_ADDR[5]), .D1(n312), .S(N1030), .Y(n605)
         );
  mx2d1_hd U1154 ( .D0(o_ADS1292_REG_ADDR[6]), .D1(n311), .S(N1030), .Y(n604)
         );
  mx2d1_hd U1155 ( .D0(o_ADS1292_REG_ADDR[7]), .D1(n310), .S(N1030), .Y(n603)
         );
  nr3d1_hd U1156 ( .A(n193), .B(gt_x_147_n12), .C(N1075), .Y(n3) );
  clknd2d1_hd U1158 ( .A(n163), .B(n911), .Y(N333) );
  mx2d1_hd U1159 ( .D0(n394), .D1(N681), .S(N718), .Y(gt_x_61_n17) );
  mx2d1_hd U1160 ( .D0(n393), .D1(N682), .S(N718), .Y(r_mpr_clk_counter[2]) );
  or2d1_hd U1162 ( .A(n526), .B(n547), .Y(N714) );
  xo2d1_hd U1164 ( .A(add_x_62_n1), .B(n391), .Y(N618) );
  mx2d1_hd U1165 ( .D0(n390), .D1(N680), .S(N718), .Y(r_mpr_clk_counter[0]) );
  mx2d1_hd U1166 ( .D0(o_MPR121_REG_ADDR[0]), .D1(n434), .S(N728), .Y(n589) );
  mx2d1_hd U1167 ( .D0(o_MPR121_REG_ADDR[1]), .D1(n433), .S(N728), .Y(n588) );
  mx2d1_hd U1168 ( .D0(o_MPR121_REG_ADDR[2]), .D1(n432), .S(N728), .Y(n587) );
  mx2d1_hd U1169 ( .D0(o_MPR121_REG_ADDR[3]), .D1(n431), .S(N728), .Y(n586) );
  mx2d1_hd U1170 ( .D0(o_MPR121_REG_ADDR[4]), .D1(n430), .S(N728), .Y(n585) );
  mx2d1_hd U1171 ( .D0(o_MPR121_REG_ADDR[5]), .D1(n429), .S(N728), .Y(n584) );
  mx2d1_hd U1172 ( .D0(o_MPR121_REG_ADDR[6]), .D1(n428), .S(N728), .Y(n583) );
  mx2d1_hd U1173 ( .D0(o_MPR121_REG_ADDR[7]), .D1(n427), .S(N728), .Y(n582) );
  mx2d1_hd U1174 ( .D0(o_ADS1292_DATA_IN[0]), .D1(n201), .S(n513), .Y(n618) );
  mx2d1_hd U1175 ( .D0(o_ADS1292_DATA_IN[1]), .D1(n194), .S(n513), .Y(n617) );
  mx2d1_hd U1176 ( .D0(o_ADS1292_DATA_IN[2]), .D1(n189), .S(n513), .Y(n616) );
  mx2d1_hd U1177 ( .D0(o_ADS1292_DATA_IN[3]), .D1(n183), .S(n513), .Y(n615) );
  mx2d1_hd U1178 ( .D0(o_ADS1292_DATA_IN[4]), .D1(n177), .S(n513), .Y(n614) );
  mx2d1_hd U1179 ( .D0(o_ADS1292_DATA_IN[5]), .D1(n175), .S(n513), .Y(n613) );
  mx2d1_hd U1180 ( .D0(o_ADS1292_DATA_IN[6]), .D1(n319), .S(n513), .Y(n612) );
  mx2d1_hd U1181 ( .D0(o_ADS1292_DATA_IN[7]), .D1(n318), .S(n513), .Y(n611) );
  mx2d1_hd U1182 ( .D0(n373), .D1(N805), .S(n491), .Y(r_ads_reg_addr[0]) );
  mx2d1_hd U1183 ( .D0(n372), .D1(N806), .S(n491), .Y(r_ads_reg_addr[1]) );
  mx2d1_hd U1184 ( .D0(n371), .D1(N807), .S(n491), .Y(r_ads_reg_addr[2]) );
  mx2d1_hd U1185 ( .D0(n370), .D1(N808), .S(n491), .Y(r_ads_reg_addr[3]) );
  mx2d1_hd U1186 ( .D0(n369), .D1(N809), .S(n491), .Y(r_ads_reg_addr[4]) );
  mx2d1_hd U1187 ( .D0(n368), .D1(N810), .S(n491), .Y(r_ads_reg_addr[5]) );
  mx2d1_hd U1188 ( .D0(n367), .D1(N811), .S(n491), .Y(r_ads_reg_addr[6]) );
  mx2d1_hd U1189 ( .D0(n366), .D1(N812), .S(n491), .Y(r_ads_reg_addr[7]) );
  mx2d1_hd U1190 ( .D0(n365), .D1(n516), .S(N1029), .Y(r_ads_run_set_done) );
  or2d1_hd U1191 ( .A(n516), .B(n545), .Y(N1029) );
  mx2d1_hd U1192 ( .D0(o_MPR121_DATA_IN[0]), .D1(n444), .S(n553), .Y(n596) );
  mx2d1_hd U1193 ( .D0(o_MPR121_DATA_IN[1]), .D1(n443), .S(n553), .Y(n595) );
  mx2d1_hd U1194 ( .D0(o_MPR121_DATA_IN[2]), .D1(n442), .S(n553), .Y(n594) );
  mx2d1_hd U1195 ( .D0(o_MPR121_DATA_IN[3]), .D1(n441), .S(n553), .Y(n593) );
  mx2d1_hd U1196 ( .D0(o_MPR121_DATA_IN[4]), .D1(n440), .S(n553), .Y(n592) );
  mx2d1_hd U1197 ( .D0(o_MPR121_DATA_IN[6]), .D1(n439), .S(n553), .Y(n591) );
  mx2d1_hd U1198 ( .D0(o_MPR121_DATA_IN[7]), .D1(n438), .S(n553), .Y(n590) );
  mx2d1_hd U1199 ( .D0(n357), .D1(n533), .S(N707), .Y(r_mpr_run_set_done) );
  nr2d1_hd U1200 ( .A(n574), .B(n539), .Y(N707) );
  ivd1_hd U1201 ( .A(n521), .Y(n574) );
  mx2d1_hd U1202 ( .D0(n356), .D1(N243), .S(N253), .Y(r_run_mode) );
  or2d1_hd U1203 ( .A(n536), .B(n557), .Y(N224) );
  mx2d1_hd U1204 ( .D0(n355), .D1(N316), .S(N331), .Y(r_mpr_run_set) );
  clknd2d1_hd U1205 ( .A(n170), .B(n911), .Y(N331) );
  mx2d1_hd U1206 ( .D0(n354), .D1(N318), .S(N332), .Y(r_mpr_read_reg) );
  ad2d1_hd U1207 ( .A(n446), .B(n180), .Y(N308) );
  mx2d1_hd U1208 ( .D0(n353), .D1(N169), .S(N155), .Y(r_uart_clk_counter[2])
         );
  mx2d1_hd U1209 ( .D0(n352), .D1(N167), .S(N155), .Y(r_uart_clk_counter[0])
         );
  mx2d1_hd U1210 ( .D0(n351), .D1(N168), .S(N155), .Y(r_uart_clk_counter[1])
         );
  mx2d1_hd U1211 ( .D0(n350), .D1(N170), .S(N155), .Y(r_uart_clk_counter[3])
         );
  xo2d1_hd U1212 ( .A(add_x_1_n1), .B(n350), .Y(N166) );
  mx2d1_hd U1213 ( .D0(n349), .D1(N319), .S(N330), .Y(r_ads_chip_set) );
  mx2d1_hd U1214 ( .D0(n348), .D1(N314), .S(N330), .Y(r_mpr_chip_set) );
  oa21d1_hd U1215 ( .A(n458), .B(N286), .C(n174), .Y(r_core_pstate[2]) );
  clknd2d1_hd U1216 ( .A(n356), .B(n563), .Y(n174) );
  ad2d1_hd U1217 ( .A(n457), .B(n468), .Y(r_chip_set) );
  ad2d1_hd U1218 ( .A(n357), .B(n365), .Y(r_run_set) );
  mx2d1_hd U1224 ( .D0(n343), .D1(N701), .S(n524), .Y(r_mpr_lstate_1_) );
  mx2d1_hd U1225 ( .D0(n342), .D1(N946), .S(N1016), .Y(r_ads_set_counter[1])
         );
  mx2d1_hd U1226 ( .D0(n341), .D1(N948), .S(N1016), .Y(r_ads_set_counter[3])
         );
  xo2d1_hd U1227 ( .A(add_x_148_n1), .B(n341), .Y(N907) );
  mx2d1_hd U1228 ( .D0(n340), .D1(N637), .S(N711), .Y(r_mpr_set_counter[2]) );
  mx2d1_hd U1229 ( .D0(n339), .D1(N638), .S(N711), .Y(r_mpr_set_counter[3]) );
  xo2d1_hd U1230 ( .A(add_x_60_n1), .B(n339), .Y(N598) );
  or3d1_hd U1232 ( .A(N63), .B(N363), .C(n544), .Y(N702) );
  mx2d1_hd U1233 ( .D0(n337), .D1(N945), .S(N1016), .Y(r_ads_set_counter[0])
         );
  mx2d1_hd U1251 ( .D0(n319), .D1(N955), .S(N1026), .Y(r_ads_second_param[6])
         );
  clknd2d1_hd U1252 ( .A(n523), .B(n52), .Y(n51) );
  mx2d1_hd U1253 ( .D0(n318), .D1(N956), .S(N1026), .Y(r_ads_second_param[7])
         );
  mx2d1_hd U1254 ( .D0(n317), .D1(N999), .S(N1026), .Y(r_ads_first_param[0])
         );
  mx2d1_hd U1255 ( .D0(n316), .D1(N1000), .S(N1026), .Y(r_ads_first_param[1])
         );
  mx2d1_hd U1256 ( .D0(n315), .D1(N1001), .S(N1026), .Y(r_ads_first_param[2])
         );
  clknd2d1_hd U1257 ( .A(n210), .B(n56), .Y(N1001) );
  mx2d1_hd U1258 ( .D0(n314), .D1(N1002), .S(N1026), .Y(r_ads_first_param[3])
         );
  mx2d1_hd U1259 ( .D0(n313), .D1(N1003), .S(N1026), .Y(r_ads_first_param[4])
         );
  mx2d1_hd U1260 ( .D0(n312), .D1(N1004), .S(N1026), .Y(r_ads_first_param[5])
         );
  mx2d1_hd U1261 ( .D0(n311), .D1(N1005), .S(N1026), .Y(r_ads_first_param[6])
         );
  mx2d1_hd U1262 ( .D0(n310), .D1(N1006), .S(N1026), .Y(r_ads_first_param[7])
         );
  or2d1_hd U1294 ( .A(n154), .B(N217), .Y(N215) );
  clknd2d1_hd U1310 ( .A(n72), .B(n73), .Y(r_mpr_pstate[5]) );
  or2d1_hd U1311 ( .A(N608), .B(n96), .Y(N627) );
  or2d1_hd U1312 ( .A(N464), .B(N1316), .Y(N473) );
  clknd2d1_hd U1313 ( .A(n82), .B(n81), .Y(r_mpr_pstate[2]) );
  or2d1_hd U1314 ( .A(n532), .B(n549), .Y(N1290) );
  clknd2d1_hd U1341 ( .A(n570), .B(n571), .Y(N1025) );
  clknd2d1_hd U1342 ( .A(N804), .B(n491), .Y(n571) );
  ivd1_hd U1343 ( .A(n197), .Y(n570) );
  oa22d1_hd U1345 ( .A(n491), .B(N1273), .C(N801), .D(N1273), .Y(n204) );
  or3d1_hd U1346 ( .A(N1032), .B(N804), .C(N802), .Y(N801) );
  clknd2d1_hd U1347 ( .A(n492), .B(n528), .Y(N1023) );
  ivd1_hd U1356 ( .A(n464), .Y(N357) );
  nr2d1_hd U1357 ( .A(N1275), .B(N795), .Y(n492) );
  clknd2d1_hd U1358 ( .A(N713), .B(N480), .Y(n573) );
  mx2d1_hd U1359 ( .D0(n230), .D1(N489), .S(N713), .Y(r_mpr_reg_addr[7]) );
  mx2d1_hd U1360 ( .D0(n229), .D1(N488), .S(N713), .Y(r_mpr_reg_addr[6]) );
  mx2d1_hd U1361 ( .D0(n228), .D1(N487), .S(N713), .Y(r_mpr_reg_addr[5]) );
  mx2d1_hd U1362 ( .D0(n227), .D1(N486), .S(N713), .Y(r_mpr_reg_addr[4]) );
  mx2d1_hd U1363 ( .D0(n226), .D1(N485), .S(N713), .Y(r_mpr_reg_addr[3]) );
  mx2d1_hd U1364 ( .D0(n225), .D1(N484), .S(N713), .Y(r_mpr_reg_addr[2]) );
  mx2d1_hd U1365 ( .D0(n224), .D1(N483), .S(N713), .Y(r_mpr_reg_addr[1]) );
  mx2d1_hd U1366 ( .D0(n223), .D1(N482), .S(N713), .Y(r_mpr_reg_addr[0]) );
  ad2d1_hd U1370 ( .A(n239), .B(n222), .Y(N791) );
  or2d1_hd U1372 ( .A(N764), .B(n222), .Y(N765) );
  or2d1_hd U1373 ( .A(N764), .B(n222), .Y(N777) );
  or2d1_hd U1374 ( .A(N764), .B(n222), .Y(N769) );
  or2d1_hd U1375 ( .A(n239), .B(n222), .Y(N743) );
  or2d1_hd U1376 ( .A(N764), .B(n222), .Y(N773) );
  or2d1_hd U1378 ( .A(n221), .B(n238), .Y(N766) );
  or2d1_hd U1379 ( .A(n221), .B(N742), .Y(N786) );
  ad2d1_hd U1380 ( .A(N791), .B(n221), .Y(N792) );
  or2d1_hd U1381 ( .A(n221), .B(n238), .Y(N782) );
  or2d1_hd U1382 ( .A(n221), .B(N742), .Y(N753) );
  or2d1_hd U1383 ( .A(n221), .B(N742), .Y(N770) );
  ivd1_hd U1384 ( .A(n221), .Y(N741) );
  or2d1_hd U1385 ( .A(n221), .B(n238), .Y(N749) );
  mx2d1_hd U1393 ( .D0(n214), .D1(N636), .S(N711), .Y(r_mpr_set_counter[1]) );
  or2d1_hd U1394 ( .A(n214), .B(N1213), .Y(N1214) );
  or2d1_hd U1395 ( .A(n214), .B(N1071), .Y(N1072) );
  or2d1_hd U1396 ( .A(n214), .B(N1209), .Y(N1210) );
  or2d1_hd U1397 ( .A(n214), .B(N1189), .Y(N1190) );
  or2d1_hd U1398 ( .A(n214), .B(N1181), .Y(N1182) );
  or2d1_hd U1399 ( .A(n214), .B(N1149), .Y(N1150) );
  or2d1_hd U1400 ( .A(n214), .B(N1157), .Y(N1158) );
  or2d1_hd U1401 ( .A(n214), .B(N1104), .Y(N1105) );
  mx2d1_hd U1402 ( .D0(n207), .D1(N947), .S(N1016), .Y(gt_x_147_n15) );
  or2d1_hd U1403 ( .A(n207), .B(N1075), .Y(N1109) );
  or2d1_hd U1404 ( .A(n207), .B(n341), .Y(N1201) );
  or2d1_hd U1405 ( .A(n207), .B(N1075), .Y(N1077) );
  or2d1_hd U1406 ( .A(n207), .B(n341), .Y(N1177) );
  or2d1_hd U1407 ( .A(n207), .B(n341), .Y(N1193) );
  or2d1_hd U1408 ( .A(n207), .B(n341), .Y(N1185) );
  or2d1_hd U1409 ( .A(n207), .B(N1075), .Y(N1136) );
  mx2d1_hd U1410 ( .D0(n201), .D1(N949), .S(N1026), .Y(r_ads_second_param[0])
         );
  mx2d1_hd U1411 ( .D0(n194), .D1(N950), .S(N1026), .Y(r_ads_second_param[1])
         );
  mx2d1_hd U1412 ( .D0(n189), .D1(N951), .S(N1026), .Y(r_ads_second_param[2])
         );
  mx2d1_hd U1413 ( .D0(n183), .D1(N952), .S(N1026), .Y(r_ads_second_param[3])
         );
  mx2d1_hd U1414 ( .D0(n177), .D1(N953), .S(N1026), .Y(r_ads_second_param[4])
         );
  mx2d1_hd U1415 ( .D0(n175), .D1(N954), .S(N1026), .Y(r_ads_second_param[5])
         );
  scg6d2_hd U1416 ( .A(N1027), .B(n195), .C(n491), .Y(N1026) );
  ad2d1_hd U1424 ( .A(N463), .B(n463), .Y(N464) );
  ad2d1_hd U1425 ( .A(N465), .B(n463), .Y(N466) );
  or2d1_hd U1426 ( .A(N357), .B(n463), .Y(N385) );
  or2d1_hd U1427 ( .A(N357), .B(n463), .Y(N434) );
  or2d1_hd U1428 ( .A(N357), .B(n463), .Y(N410) );
  or2d1_hd U1429 ( .A(N357), .B(n463), .Y(N360) );
  ivd1_hd U1430 ( .A(n463), .Y(N350) );
  ad2d1_hd U1431 ( .A(n460), .B(n464), .Y(N463) );
  ad2d1_hd U1432 ( .A(N343), .B(n464), .Y(N465) );
  or2d1_hd U1433 ( .A(n464), .B(N350), .Y(N453) );
  or2d1_hd U1434 ( .A(n464), .B(n463), .Y(N373) );
  or2d1_hd U1435 ( .A(n464), .B(N350), .Y(N428) );
  or2d1_hd U1436 ( .A(n464), .B(N350), .Y(N379) );
  or2d1_hd U1437 ( .A(n464), .B(n463), .Y(N398) );
  or2d1_hd U1438 ( .A(n464), .B(N350), .Y(N404) );
  or2d1_hd U1439 ( .A(n464), .B(n463), .Y(N422) );
  or2d1_hd U1440 ( .A(n464), .B(n463), .Y(N447) );
  or2d1_hd U1441 ( .A(n464), .B(n463), .Y(N346) );
  or2d1_hd U1442 ( .A(n464), .B(N350), .Y(N353) );
  nr2ad1_hd U1444 ( .A(n154), .B(n10), .Y(N216) );
  mx2d1_hd U1445 ( .D0(n154), .D1(N1013), .S(N1018), .Y(r_ads_data_send_ready)
         );
  ivd1_hd U1446 ( .A(n154), .Y(alt36_n332) );
  ivd1_hd U1460 ( .A(n346), .Y(N1040) );
  ivd1_hd U1462 ( .A(n345), .Y(N1039) );
  ivd1_hd U1466 ( .A(n461), .Y(N276) );
  ivd1_hd U1468 ( .A(n75), .Y(N154) );
  ivd1_hd U1470 ( .A(n465), .Y(N153) );
  ivd1_hd U1472 ( .A(n343), .Y(N1050) );
  ivd1_hd U1474 ( .A(n342), .Y(N1076) );
  ivd1_hd U1476 ( .A(n341), .Y(N1075) );
  ivd1_hd U1478 ( .A(n340), .Y(N1069) );
  ivd1_hd U1479 ( .A(n339), .Y(N1068) );
  nr2d1_hd U1482 ( .A(N417), .B(N416), .Y(n512) );
  nr2d1_hd U1483 ( .A(N399), .B(N398), .Y(n514) );
  scg6d1_hd U1484 ( .A(n526), .B(N481), .C(n79), .Y(r_mpr_pstate[3]) );
  or2d1_hd U1485 ( .A(N1070), .B(N1133), .Y(N1134) );
  or2d1_hd U1486 ( .A(n408), .B(N1105), .Y(N1106) );
  or2d1_hd U1487 ( .A(N1070), .B(N1198), .Y(N1199) );
  nr2d1_hd U1488 ( .A(N752), .B(N753), .Y(n516) );
  nr2d1_hd U1489 ( .A(N1108), .B(N1178), .Y(n517) );
  nr2d1_hd U1490 ( .A(N386), .B(N385), .Y(n518) );
  nr2d1_hd U1491 ( .A(N423), .B(N422), .Y(n519) );
  ad2d1_hd U1492 ( .A(N153), .B(N154), .Y(N155) );
  scg9d1_hd U1493 ( .A(gt_x_61_n12), .B(n391), .C(gt_x_61_n7), .Y(n520) );
  nr2d1_hd U1494 ( .A(N392), .B(N391), .Y(n521) );
  or2d1_hd U1495 ( .A(N285), .B(N276), .Y(N286) );
  scg8d1_hd U1496 ( .A(N607), .B(n74), .C(N1259), .D(n76), .Y(r_mpr_pstate[4])
         );
  nr2d1_hd U1497 ( .A(N1108), .B(N1146), .Y(n523) );
  or3d1_hd U1498 ( .A(N701), .B(n68), .C(n69), .Y(n524) );
  clknd2d1_hd U1499 ( .A(i_MPR121_INIT_SET), .B(i_ADS1292_INIT_SET), .Y(n525)
         );
  or2d1_hd U1500 ( .A(N1108), .B(N1162), .Y(N1163) );
  scg10d1_hd U1501 ( .A(alt36_n60), .B(n202), .C(alt36_n508), .D(n203), .Y(
        n528) );
  nr2d1_hd U1502 ( .A(N411), .B(N410), .Y(n529) );
  nr2d1_hd U1503 ( .A(N777), .B(N778), .Y(n530) );
  nr2d1_hd U1504 ( .A(N441), .B(N440), .Y(n531) );
  or2d1_hd U1505 ( .A(N1070), .B(N1150), .Y(N1151) );
  or2d1_hd U1506 ( .A(N1108), .B(N1110), .Y(N1111) );
  or2d1_hd U1507 ( .A(n408), .B(N1206), .Y(N1207) );
  or2d1_hd U1508 ( .A(n337), .B(N1186), .Y(N1187) );
  or2d1_hd U1509 ( .A(n408), .B(N1174), .Y(N1175) );
  or2d1_hd U1510 ( .A(n408), .B(N1158), .Y(N1159) );
  nr2d1_hd U1511 ( .A(N435), .B(N434), .Y(n532) );
  ivd1_hd U1512 ( .A(n214), .Y(N1131) );
  nr2d1_hd U1513 ( .A(n436), .B(N1056), .Y(n533) );
  nr2d1_hd U1514 ( .A(N380), .B(N379), .Y(n534) );
  nr2d1_hd U1515 ( .A(N785), .B(N786), .Y(n535) );
  ivd1_hd U1516 ( .A(n405), .Y(gt_x_149_n10) );
  nr2d1_hd U1517 ( .A(n346), .B(N1128), .Y(n536) );
  or2d1_hd U1518 ( .A(N153), .B(n75), .Y(N158) );
  clknd2d1_hd U1520 ( .A(r_run_mode), .B(r_run_set), .Y(n537) );
  clknd2d1_hd U1521 ( .A(n352), .B(N1092), .Y(n538) );
  nr2d1_hd U1522 ( .A(n533), .B(n565), .Y(n539) );
  or2d1_hd U1523 ( .A(i_MPR121_FAIL), .B(i_MPR121_BUSY), .Y(alt36_n159) );
  ivd1_hd U1524 ( .A(alt36_n159), .Y(n96) );
  nr2d1_hd U1525 ( .A(i_ADS1292_FILTERED_DATA_VALID), .B(N929), .Y(n540) );
  ivd1_hd U1526 ( .A(n207), .Y(N1144) );
  nr2d1_hd U1527 ( .A(n337), .B(N1137), .Y(n541) );
  or2d1_hd U1528 ( .A(n337), .B(N1154), .Y(N1155) );
  nr2d4_hd U1529 ( .A(N781), .B(N782), .Y(n542) );
  nr2d1_hd U1530 ( .A(n465), .B(N154), .Y(n543) );
  nr2d1_hd U1531 ( .A(N367), .B(N366), .Y(n544) );
  ivd1_hd U1532 ( .A(N430), .Y(N431) );
  nr2d1_hd U1533 ( .A(N756), .B(N757), .Y(n545) );
  nr2d1_hd U1534 ( .A(N769), .B(N770), .Y(n546) );
  or4d1_hd U1535 ( .A(N751), .B(n545), .C(n530), .D(N795), .Y(N1273) );
  nr2d1_hd U1536 ( .A(N448), .B(N447), .Y(n547) );
  nr2d1_hd U1537 ( .A(N405), .B(N404), .Y(n548) );
  or2d1_hd U1538 ( .A(N1070), .B(N1072), .Y(N1073) );
  or2d1_hd U1539 ( .A(n408), .B(N1141), .Y(N1142) );
  or2d1_hd U1540 ( .A(n337), .B(N1078), .Y(N1079) );
  nr2d1_hd U1541 ( .A(N454), .B(N453), .Y(n549) );
  or2d1_hd U1542 ( .A(N1108), .B(N1194), .Y(N1195) );
  or3d1_hd U1543 ( .A(n526), .B(N363), .C(n544), .Y(N1303) );
  nr3d1_hd U1544 ( .A(N1240), .B(N1229), .C(N795), .Y(n550) );
  ivd1_hd U1545 ( .A(N362), .Y(N363) );
  or2d1_hd U1546 ( .A(N1070), .B(N1210), .Y(N1211) );
  ivd1_hd U1547 ( .A(n337), .Y(N1108) );
  or2d1_hd U1548 ( .A(N1070), .B(N1182), .Y(N1183) );
  or2d1_hd U1549 ( .A(N1070), .B(N1166), .Y(N1167) );
  or2d1_hd U1550 ( .A(n408), .B(N1190), .Y(N1191) );
  clknd2d1_hd U1551 ( .A(n11), .B(n12), .Y(N1294) );
  nr2d1_hd U1552 ( .A(n337), .B(N1202), .Y(n551) );
  or3d1_hd U1553 ( .A(N363), .B(n544), .C(N462), .Y(N701) );
  or4d1_hd U1554 ( .A(N1256), .B(N1257), .C(N1258), .D(N473), .Y(N1259) );
  or2d1_hd U1555 ( .A(N1289), .B(N1290), .Y(N1291) );
  or2d1_hd U1556 ( .A(N1270), .B(n532), .Y(N1271) );
  nr2d1_hd U1557 ( .A(n491), .B(n535), .Y(n552) );
  ivd1_hd U1558 ( .A(N1171), .Y(N1172) );
  ivd1_hd U1559 ( .A(N767), .Y(N768) );
  scg9d1_hd U1560 ( .A(gt_x_149_n12), .B(n405), .C(gt_x_149_n10), .Y(n554) );
  clknd2d1_hd U1561 ( .A(n348), .B(N297), .Y(n555) );
  or2d1_hd U1562 ( .A(N363), .B(n544), .Y(N1299) );
  clknd2d1_hd U1563 ( .A(N1317), .B(n357), .Y(n556) );
  nr2d1_hd U1564 ( .A(N1040), .B(N1120), .Y(n557) );
  nr2d1_hd U1565 ( .A(n408), .B(N1214), .Y(n558) );
  nr2d1_hd U1566 ( .A(N1040), .B(N1101), .Y(n559) );
  nr2d1_hd U1567 ( .A(N1040), .B(N1046), .Y(n560) );
  or2d1_hd U1568 ( .A(N1069), .B(N1131), .Y(n561) );
  or4d1_hd U1569 ( .A(n553), .B(n514), .C(n519), .D(n532), .Y(N1286) );
  or3d1_hd U1570 ( .A(n516), .B(n542), .C(n535), .Y(N1278) );
  ivd1_hd U1571 ( .A(N155), .Y(n182) );
  ivd1_hd U1572 ( .A(n365), .Y(N303) );
  ivd1_hd U1573 ( .A(n357), .Y(N302) );
  nr2d1_hd U1576 ( .A(N1059), .B(N1065), .Y(n562) );
  nr2d1_hd U1577 ( .A(N288), .B(n461), .Y(n563) );
  nr2d1_hd U1579 ( .A(n533), .B(n562), .Y(n565) );
  nr2d1_hd U1580 ( .A(n466), .B(N1088), .Y(n566) );
  fd3qd1_hd clk_r_REG250_S4 ( .D(1'b0), .CK(n932), .SN(n767), .Q(n467) );
  fd3qd1_hd clk_r_REG251_S4 ( .D(1'b0), .CK(n932), .SN(n767), .Q(n466) );
  fd3qd1_hd clk_r_REG155_S7 ( .D(n537), .CK(i_CLK), .SN(n767), .Q(n458) );
  fd3qd1_hd clk_r_REG82_S4 ( .D(N1022), .CK(n930), .SN(n767), .Q(n238) );
  fd3qd1_hd clk_r_REG77_S4 ( .D(N1023), .CK(n930), .SN(n767), .Q(n221) );
  fd3qd1_hd clk_r_REG136_S4 ( .D(r_mpr_pstate[4]), .CK(i_CLK), .SN(n767), .Q(
        n67) );
  fd4qd1_hd clk_r_REG273_S2 ( .D(r_uart_clk_counter[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n350) );
  fd4qd1_hd clk_r_REG109_S2 ( .D(r_mpr_read_reg), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n354) );
  fd4qd1_hd clk_r_REG51_S2 ( .D(r_ads_read_reg), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n426) );
  fd4qd1_hd clk_r_REG275_S2 ( .D(r_uart_clk_counter[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n352) );
  fd4qd1_hd clk_r_REG274_S2 ( .D(r_uart_clk_counter[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n351) );
  fd4qd1_hd clk_r_REG162_S9 ( .D(r_mpr_chip_set), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n348) );
  fd4qd1_hd clk_r_REG161_S9 ( .D(r_ads_chip_set), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n349) );
  fd4qd1_hd clk_r_REG160_S7 ( .D(r_mpr_run_set), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n355) );
  fd4qd1_hd clk_r_REG182_S6 ( .D(n590), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_DATA_IN[7]) );
  fd4qd1_hd clk_r_REG180_S6 ( .D(n591), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_MPR121_DATA_IN[6]) );
  fd4qd1_hd clk_r_REG176_S6 ( .D(n593), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_MPR121_DATA_IN[3]) );
  fd4qd1_hd clk_r_REG174_S6 ( .D(n594), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_DATA_IN[2]) );
  fd4qd1_hd clk_r_REG248_S4 ( .D(r_ads_set_counter[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n337) );
  fd4qd1_hd clk_r_REG218_S5 ( .D(r_ads_clk_counter[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n404) );
  fd4qd1_hd clk_r_REG217_S5 ( .D(gt_x_149_n17), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n407) );
  fd4qd1_hd clk_r_REG216_S5 ( .D(r_ads_clk_counter[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n406) );
  fd4qd1_hd clk_r_REG215_S5 ( .D(gt_x_149_n9), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(n405) );
  fd4qd1_hd clk_r_REG247_S4 ( .D(gt_x_147_n15), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n207) );
  fd4qd1_hd clk_r_REG245_S4 ( .D(r_ads_set_counter[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n341) );
  fd4qd1_hd clk_r_REG236_S4 ( .D(r_ads_set_counter[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n342) );
  fd4qd1_hd clk_r_REG185_S7 ( .D(r_chip_set), .CK(i_CLK), .SN(1'b1), .RN(n636), 
        .Q(n462) );
  fd4qd1_hd clk_r_REG156_S8 ( .D(r_core_pstate[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n347) );
  fd4qd1_hd clk_r_REG154_S6 ( .D(r_mpr_run_set_done), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n357) );
  fd4qd1_hd clk_r_REG152_S6 ( .D(n599), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_ERROR) );
  fd4qd1_hd clk_r_REG271_S2 ( .D(r_uart_clk_counter[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n353) );
  fd4qd1_hd clk_r_REG252_S5 ( .D(r_ads_run_set_done), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n365) );
  fd4qd1_hd clk_r_REG226_S5 ( .D(n611), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[7]) );
  fd4qd1_hd clk_r_REG225_S5 ( .D(n612), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[6]) );
  fd4qd1_hd clk_r_REG224_S5 ( .D(n613), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[5]) );
  fd4qd1_hd clk_r_REG223_S5 ( .D(n614), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[4]) );
  fd4qd1_hd clk_r_REG222_S5 ( .D(n615), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[3]) );
  fd4qd1_hd clk_r_REG221_S5 ( .D(n616), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[2]) );
  fd4qd1_hd clk_r_REG220_S5 ( .D(n617), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[1]) );
  fd4qd1_hd clk_r_REG219_S5 ( .D(n618), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_DATA_IN[0]) );
  fd4qd1_hd clk_r_REG214_S5 ( .D(r_mpr_clk_counter[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n390) );
  fd4qd1_hd clk_r_REG213_S5 ( .D(r_mpr_clk_counter[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n393) );
  fd4qd1_hd clk_r_REG211_S5 ( .D(gt_x_61_n17), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(n394) );
  fd4qd1_hd clk_r_REG178_S6 ( .D(n592), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_DATA_IN[4]) );
  fd4qd1_hd clk_r_REG172_S6 ( .D(n595), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_MPR121_DATA_IN[1]) );
  fd4qd1_hd clk_r_REG170_S6 ( .D(n596), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_DATA_IN[0]) );
  fd4qd1_hd clk_r_REG73_S3 ( .D(r_ads_reg_addr[7]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n366) );
  fd4qd1_hd clk_r_REG70_S3 ( .D(r_ads_reg_addr[6]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n367) );
  fd4qd1_hd clk_r_REG69_S3 ( .D(r_ads_reg_addr[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n372) );
  fd4qd1_hd clk_r_REG66_S3 ( .D(r_ads_reg_addr[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n371) );
  fd4qd1_hd clk_r_REG63_S3 ( .D(r_ads_reg_addr[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n370) );
  fd4qd1_hd clk_r_REG60_S3 ( .D(r_ads_reg_addr[4]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n369) );
  fd4qd1_hd clk_r_REG57_S3 ( .D(r_ads_reg_addr[5]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n368) );
  fd4qd1_hd clk_r_REG54_S3 ( .D(r_ads_reg_addr[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n373) );
  fd4qd1_hd clk_r_REG254_S2 ( .D(r_run_mode), .CK(i_CLK), .SN(1'b1), .RN(n768), 
        .Q(n356) );
  fd4qd1_hd clk_r_REG75_S4 ( .D(n603), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_REG_ADDR[7]) );
  fd4qd1_hd clk_r_REG72_S4 ( .D(n604), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_ADS1292_REG_ADDR[6]) );
  fd4qd1_hd clk_r_REG68_S4 ( .D(n609), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_REG_ADDR[1]) );
  fd4qd1_hd clk_r_REG65_S4 ( .D(n608), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_ADS1292_REG_ADDR[2]) );
  fd4qd1_hd clk_r_REG62_S4 ( .D(n607), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_REG_ADDR[3]) );
  fd4qd1_hd clk_r_REG59_S4 ( .D(n606), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_ADS1292_REG_ADDR[4]) );
  fd4qd1_hd clk_r_REG56_S4 ( .D(n605), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_REG_ADDR[5]) );
  fd4qd1_hd clk_r_REG53_S4 ( .D(n610), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_ADS1292_REG_ADDR[0]) );
  fd4qd1_hd clk_r_REG132_S4 ( .D(n582), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[7]) );
  fd4qd1_hd clk_r_REG129_S4 ( .D(n583), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[6]) );
  fd4qd1_hd clk_r_REG126_S4 ( .D(n589), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[0]) );
  fd4qd1_hd clk_r_REG123_S4 ( .D(n588), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[1]) );
  fd4qd1_hd clk_r_REG120_S4 ( .D(n587), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[2]) );
  fd4qd1_hd clk_r_REG117_S4 ( .D(n586), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[3]) );
  fd4qd1_hd clk_r_REG114_S4 ( .D(n585), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[4]) );
  fd4qd1_hd clk_r_REG111_S4 ( .D(n584), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_REG_ADDR[5]) );
  fd4qd1_hd clk_r_REG78_S5 ( .D(n601), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_ADS1292_CONTROL[1]) );
  fd4qd1_hd clk_r_REG80_S5 ( .D(n602), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_ADS1292_CONTROL[0]) );
  fd4qd1_hd clk_r_REG79_S5 ( .D(n600), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_ADS1292_CONTROL[2]) );
  fd4qd1_hd clk_r_REG189_S6 ( .D(r_mpr_set_counter[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n408) );
  fd4qd1_hd clk_r_REG168_S4 ( .D(n598), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_READ_ENABLE) );
  fd4qd1_hd clk_r_REG167_S4 ( .D(n597), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        o_MPR121_WRITE_ENABLE) );
  fd4qd1_hd clk_r_REG133_S3 ( .D(r_mpr_reg_addr[7]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n230) );
  fd4qd1_hd clk_r_REG130_S3 ( .D(r_mpr_reg_addr[6]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n229) );
  fd4qd1_hd clk_r_REG127_S3 ( .D(r_mpr_reg_addr[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n223) );
  fd4qd1_hd clk_r_REG124_S3 ( .D(r_mpr_reg_addr[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n224) );
  fd4qd1_hd clk_r_REG121_S3 ( .D(r_mpr_reg_addr[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n225) );
  fd4qd1_hd clk_r_REG118_S3 ( .D(r_mpr_reg_addr[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n226) );
  fd4qd1_hd clk_r_REG115_S3 ( .D(r_mpr_reg_addr[4]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n227) );
  fd4qd1_hd clk_r_REG112_S3 ( .D(r_mpr_reg_addr[5]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n228) );
  fd4qd1_hd clk_r_REG243_S5 ( .D(r_ads_second_param[4]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n177) );
  fd4qd1_hd clk_r_REG242_S5 ( .D(r_ads_second_param[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n183) );
  fd4qd1_hd clk_r_REG240_S5 ( .D(r_ads_second_param[6]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n319) );
  fd4qd1_hd clk_r_REG239_S5 ( .D(r_ads_second_param[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n201) );
  fd4qd1_hd clk_r_REG238_S5 ( .D(r_ads_second_param[7]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n318) );
  fd4qd1_hd clk_r_REG74_S3 ( .D(r_ads_first_param[7]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n310) );
  fd4qd1_hd clk_r_REG71_S3 ( .D(r_ads_first_param[6]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n311) );
  fd4qd1_hd clk_r_REG67_S3 ( .D(r_ads_first_param[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n316) );
  fd4qd1_hd clk_r_REG64_S3 ( .D(r_ads_first_param[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n315) );
  fd4qd1_hd clk_r_REG61_S3 ( .D(r_ads_first_param[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n314) );
  fd4qd1_hd clk_r_REG58_S3 ( .D(r_ads_first_param[4]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n313) );
  fd4qd1_hd clk_r_REG55_S3 ( .D(r_ads_first_param[5]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n312) );
  fd4qd1_hd clk_r_REG52_S3 ( .D(r_ads_first_param[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n317) );
  fd4qd1_hd clk_r_REG237_S5 ( .D(r_ads_second_param[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n189) );
  fd4qd1_hd clk_r_REG241_S5 ( .D(r_ads_second_param[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n194) );
  fd4qd1_hd clk_r_REG244_S5 ( .D(r_ads_second_param[5]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n175) );
  fd4qd1_hd clk_r_REG188_S6 ( .D(r_mpr_set_counter[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n214) );
  fd4qd1_hd clk_r_REG187_S6 ( .D(r_mpr_set_counter[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n340) );
  fd4qd1_hd clk_r_REG186_S6 ( .D(r_mpr_set_counter[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n339) );
  fd4qd1_hd clk_r_REG148_S5 ( .D(r_mpr_touch_status[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n423) );
  fd4qd1_hd clk_r_REG147_S5 ( .D(r_mpr_touch_status[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n422) );
  fd4qd1_hd clk_r_REG146_S5 ( .D(r_mpr_touch_status[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n421) );
  fd4qd1_hd clk_r_REG145_S5 ( .D(r_mpr_touch_status[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n420) );
  fd4qd1_hd clk_r_REG144_S5 ( .D(r_mpr_touch_status[4]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n419) );
  fd4qd1_hd clk_r_REG143_S5 ( .D(r_mpr_touch_status[5]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n418) );
  fd4qd1_hd clk_r_REG142_S5 ( .D(r_mpr_touch_status[6]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n417) );
  fd4qd1_hd clk_r_REG141_S5 ( .D(r_mpr_touch_status[7]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n416) );
  fd4qd1_hd clk_r_REG140_S5 ( .D(r_mpr_touch_status[8]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n415) );
  fd4qd1_hd clk_r_REG139_S5 ( .D(r_mpr_touch_status[9]), .CK(i_CLK), .SN(1'b1), 
        .RN(n636), .Q(n414) );
  fd4qd1_hd clk_r_REG138_S5 ( .D(r_mpr_touch_status[10]), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(n413) );
  fd4qd1_hd clk_r_REG137_S5 ( .D(r_mpr_touch_status[11]), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(n412) );
  fd4qd1_hd clk_r_REG164_S6 ( .D(r_mpr_lstate_1_), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n343) );
  fd4qd1_hd clk_r_REG153_S5 ( .D(N1052), .CK(i_CLK), .SN(1'b1), .RN(n767), .Q(
        n435) );
  fd4qd1_hd clk_r_REG181_S5 ( .D(r_mpr_second_param[7]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n438) );
  fd4qd1_hd clk_r_REG179_S5 ( .D(r_mpr_second_param[6]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n439) );
  fd4qd1_hd clk_r_REG177_S5 ( .D(r_mpr_second_param[4]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n440) );
  fd4qd1_hd clk_r_REG175_S5 ( .D(r_mpr_second_param[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n441) );
  fd4qd1_hd clk_r_REG173_S5 ( .D(r_mpr_second_param[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n442) );
  fd4qd1_hd clk_r_REG171_S5 ( .D(r_mpr_second_param[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n443) );
  fd4qd1_hd clk_r_REG169_S5 ( .D(r_mpr_second_param[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n444) );
  fd4qd1_hd clk_r_REG131_S3 ( .D(r_mpr_first_param[7]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n427) );
  fd4qd1_hd clk_r_REG128_S3 ( .D(r_mpr_first_param[6]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n428) );
  fd4qd1_hd clk_r_REG125_S3 ( .D(r_mpr_first_param[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n434) );
  fd4qd1_hd clk_r_REG122_S3 ( .D(r_mpr_first_param[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n433) );
  fd4qd1_hd clk_r_REG119_S3 ( .D(r_mpr_first_param[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n432) );
  fd4qd1_hd clk_r_REG116_S3 ( .D(r_mpr_first_param[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n431) );
  fd4qd1_hd clk_r_REG113_S3 ( .D(r_mpr_first_param[4]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n430) );
  fd4qd1_hd clk_r_REG110_S3 ( .D(r_mpr_first_param[5]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n429) );
  fd4qd1_hd clk_r_REG270_S1 ( .D(r_uart_pstate[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n767), .Q(n465) );
  fd4qd1_hd clk_r_REG157_S8 ( .D(r_core_pstate[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n78) );
  fd2qd1_hd clk_r_REG1_S1 ( .D(1'b1), .CK(n924), .RN(n768), .Q(
        o_UART_DATA_TX[53]) );
  fd2d1_hd clk_r_REG255_S1 ( .D(N240), .CK(n926), .RN(n767), .QN(N1038) );
  fd2d1_hd clk_r_REG81_S5 ( .D(N1024), .CK(n930), .RN(n767), .Q(n222), .QN(
        N747) );
  fd2d1_hd clk_r_REG268_S1 ( .D(N227), .CK(n926), .RN(n767), .QN(n162) );
  fd2d1_hd clk_r_REG267_S1 ( .D(N228), .CK(n926), .RN(n767), .QN(n161) );
  fd2d1_hd clk_r_REG266_S1 ( .D(N229), .CK(n926), .RN(n767), .QN(n160) );
  fd2d1_hd clk_r_REG265_S1 ( .D(N230), .CK(n926), .RN(n767), .QN(n159) );
  fd2d1_hd clk_r_REG264_S1 ( .D(N231), .CK(n926), .RN(n767), .QN(n158) );
  nr2d2_hd U2 ( .A(N743), .B(N744), .Y(n491) );
  ivd1_hd U52 ( .A(n9), .Y(N217) );
  clknd2d1_hd U53 ( .A(n202), .B(n206), .Y(N1014) );
  nid4_hd U464 ( .A(n767), .Y(n768) );
  nid2_hd U465 ( .A(n636), .Y(n767) );
  fd3qd1_hd clk_r_REG166_S5 ( .D(n933), .CK(i_CLK), .SN(n767), .Q(n338) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_18 clk_gate_clk_r_REG249_S4_0 ( .CLK(i_CLK), 
        .EN(N1027), .ENCLK(n932), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_19 clk_gate_clk_r_REG202_S6_0 ( .CLK(i_CLK), 
        .EN(N716), .ENCLK(n931), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_20 clk_gate_clk_r_REG81_S5_0 ( .CLK(i_CLK), 
        .EN(N1021), .ENCLK(n930), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_21 clk_gate_clk_r_REG210_S6_0 ( .CLK(i_CLK), 
        .EN(N715), .ENCLK(n929), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_22 clk_gate_clk_r_REG198_S6_0 ( .CLK(i_CLK), 
        .EN(N710), .ENCLK(n928), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_23 clk_gate_clk_r_REG235_S5_0 ( .CLK(i_CLK), 
        .EN(N1014), .ENCLK(n927), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_24 clk_gate_clk_r_REG264_S1_0 ( .CLK(i_CLK), 
        .EN(N252), .ENCLK(n926), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_25 clk_gate_clk_r_REG83_S5_0 ( .CLK(i_CLK), 
        .EN(N1017), .ENCLK(n925), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_sensor_core_26 clk_gate_clk_r_REG49_S1_0 ( .CLK(i_CLK), 
        .EN(N251), .ENCLK(n924), .TE(1'b0) );
  fd2qd1_hd R_2_clk_r_REG31_S1 ( .D(n154), .CK(n924), .RN(n636), .Q(
        o_UART_DATA_TX[49]) );
  fd2qd1_hd R_3_clk_r_REG39_S1 ( .D(n961), .CK(n924), .RN(n768), .Q(
        o_UART_DATA_TX[48]) );
  fd4qd1_hd clk_r_REG249_S4 ( .D(n908), .CK(n932), .SN(1'b1), .RN(n636), .Q(
        n909) );
  fd4qd1_hd clk_r_REG269_S1 ( .D(N226), .CK(n926), .SN(1'b1), .RN(n636), .Q(
        n906) );
  fd4qd1_hd clk_r_REG246_S5 ( .D(r_ads_chip_set_done), .CK(n930), .SN(1'b1), 
        .RN(n636), .Q(n468) );
  fd4qd2_hd clk_r_REG183_S5 ( .D(r_mpr_pstate[5]), .CK(i_CLK), .SN(1'b1), .RN(
        n636), .Q(n460) );
  fd4qd1_hd clk_r_REG30_S1 ( .D(N185), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[19]) );
  fd4qd1_hd clk_r_REG29_S1 ( .D(N184), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[18]) );
  fd4qd1_hd clk_r_REG28_S1 ( .D(N183), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[17]) );
  fd4qd1_hd clk_r_REG27_S1 ( .D(N182), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[16]) );
  fd4qd1_hd clk_r_REG26_S1 ( .D(N181), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[15]) );
  fd4qd1_hd clk_r_REG25_S1 ( .D(N180), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[14]) );
  fd4qd1_hd clk_r_REG24_S1 ( .D(N179), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[13]) );
  fd4qd1_hd clk_r_REG23_S1 ( .D(N178), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[12]) );
  fd4qd1_hd clk_r_REG22_S1 ( .D(N177), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[11]) );
  fd4qd1_hd clk_r_REG21_S1 ( .D(N176), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[10]) );
  fd4qd1_hd clk_r_REG20_S1 ( .D(N175), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[9]) );
  fd4qd1_hd clk_r_REG19_S1 ( .D(N174), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[8]) );
  fd4qd1_hd clk_r_REG2_S1 ( .D(N217), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[50]) );
  fd4qd1_hd clk_r_REG235_S5 ( .D(n527), .CK(n927), .SN(1'b1), .RN(n636), .Q(
        n447) );
  fd4qd1_hd clk_r_REG18_S1 ( .D(N213), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[47]) );
  fd4qd1_hd clk_r_REG16_S1 ( .D(N211), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[45]) );
  fd4qd1_hd clk_r_REG15_S1 ( .D(N210), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[44]) );
  fd4qd1_hd clk_r_REG14_S1 ( .D(N209), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[43]) );
  fd4qd1_hd clk_r_REG13_S1 ( .D(N208), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[42]) );
  fd4qd1_hd clk_r_REG12_S1 ( .D(N207), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[41]) );
  fd4qd1_hd clk_r_REG11_S1 ( .D(N206), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[40]) );
  fd4qd1_hd clk_r_REG10_S1 ( .D(N205), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[39]) );
  fd4qd1_hd clk_r_REG9_S1 ( .D(N204), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[38]) );
  fd4qd1_hd clk_r_REG8_S1 ( .D(N203), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[37]) );
  fd4qd1_hd clk_r_REG7_S1 ( .D(N202), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[36]) );
  fd4qd1_hd clk_r_REG6_S1 ( .D(N201), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[35]) );
  fd4qd1_hd clk_r_REG5_S1 ( .D(N200), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[34]) );
  fd4qd1_hd clk_r_REG4_S1 ( .D(N199), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[33]) );
  fd4qd1_hd clk_r_REG3_S1 ( .D(N198), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[32]) );
  fd4qd1_hd clk_r_REG158_S9 ( .D(n939), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        n395) );
  fd4qd1_hd clk_r_REG198_S6 ( .D(n529), .CK(n928), .SN(1'b1), .RN(n636), .Q(
        n270) );
  fd4qd1_hd clk_r_REG49_S1 ( .D(N197), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[31]) );
  fd4qd1_hd clk_r_REG48_S1 ( .D(N196), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[30]) );
  fd4qd1_hd clk_r_REG47_S1 ( .D(N195), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[29]) );
  fd4qd1_hd clk_r_REG46_S1 ( .D(N194), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[28]) );
  fd4qd1_hd clk_r_REG45_S1 ( .D(N193), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[27]) );
  fd4qd1_hd clk_r_REG44_S1 ( .D(N192), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[26]) );
  fd4qd1_hd clk_r_REG43_S1 ( .D(N191), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[25]) );
  fd4qd1_hd clk_r_REG42_S1 ( .D(N190), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[24]) );
  fd4qd1_hd clk_r_REG41_S1 ( .D(N215), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[51]) );
  fd4qd1_hd clk_r_REG17_S1 ( .D(N212), .CK(n924), .SN(1'b1), .RN(n636), .Q(
        o_UART_DATA_TX[46]) );
  fd4qd1_hd clk_r_REG149_S5 ( .D(n940), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        n392) );
  fd4qd1_hd clk_r_REG184_S6 ( .D(n937), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        n457) );
  fd4qd1_hd clk_r_REG212_S5 ( .D(n936), .CK(i_CLK), .SN(1'b1), .RN(n636), .Q(
        n391) );
  fd4qd1_hd clk_r_REG234_S5 ( .D(N943), .CK(n927), .SN(1'b1), .RN(n636), .Q(
        n448) );
  fd4qd1_hd clk_r_REG233_S5 ( .D(N942), .CK(n927), .SN(1'b1), .RN(n636), .Q(
        n449) );
  fd4qd1_hd clk_r_REG232_S5 ( .D(N941), .CK(n927), .SN(1'b1), .RN(n636), .Q(
        n450) );
  fd4qd1_hd clk_r_REG231_S5 ( .D(N940), .CK(n927), .SN(1'b1), .RN(n636), .Q(
        n451) );
  fd4qd1_hd clk_r_REG230_S5 ( .D(N939), .CK(n927), .SN(1'b1), .RN(n636), .Q(
        n452) );
  fd4qd1_hd clk_r_REG229_S5 ( .D(N938), .CK(n927), .SN(1'b1), .RN(n768), .Q(
        n453) );
  fd4qd1_hd clk_r_REG228_S5 ( .D(N937), .CK(n927), .SN(1'b1), .RN(n768), .Q(
        n454) );
  fd4qd1_hd clk_r_REG227_S5 ( .D(N936), .CK(n927), .SN(1'b1), .RN(n768), .Q(
        n455) );
  fd4qd1_hd clk_r_REG106_S5 ( .D(N958), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n263) );
  fd4qd1_hd clk_r_REG105_S5 ( .D(N959), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n262) );
  fd4qd1_hd clk_r_REG104_S5 ( .D(N960), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n261) );
  fd4qd1_hd clk_r_REG103_S5 ( .D(N961), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n260) );
  fd4qd1_hd clk_r_REG102_S5 ( .D(N962), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n259) );
  fd4qd1_hd clk_r_REG101_S5 ( .D(N963), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n258) );
  fd4qd1_hd clk_r_REG100_S5 ( .D(N964), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n257) );
  fd4qd1_hd clk_r_REG99_S5 ( .D(N965), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n256) );
  fd4qd1_hd clk_r_REG98_S5 ( .D(N966), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n255) );
  fd4qd1_hd clk_r_REG97_S5 ( .D(N967), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n254) );
  fd4qd1_hd clk_r_REG96_S5 ( .D(N968), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n253) );
  fd4qd1_hd clk_r_REG95_S5 ( .D(N969), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n252) );
  fd4qd1_hd clk_r_REG94_S5 ( .D(N970), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n251) );
  fd4qd1_hd clk_r_REG93_S5 ( .D(N971), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n250) );
  fd4qd1_hd clk_r_REG92_S5 ( .D(N972), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n249) );
  fd4qd1_hd clk_r_REG91_S5 ( .D(N973), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n248) );
  fd4qd1_hd clk_r_REG90_S5 ( .D(N974), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n247) );
  fd4qd1_hd clk_r_REG89_S5 ( .D(N975), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n246) );
  fd4qd1_hd clk_r_REG88_S5 ( .D(N976), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n245) );
  fd4qd1_hd clk_r_REG87_S5 ( .D(N977), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n244) );
  fd4qd1_hd clk_r_REG86_S5 ( .D(N978), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n243) );
  fd4qd1_hd clk_r_REG85_S5 ( .D(N979), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n242) );
  fd4qd1_hd clk_r_REG84_S5 ( .D(N980), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n241) );
  fd4qd1_hd clk_r_REG83_S5 ( .D(N981), .CK(n925), .SN(1'b1), .RN(n768), .Q(
        n240) );
  fd4qd1_hd clk_r_REG263_S1 ( .D(N232), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n237) );
  fd4qd1_hd clk_r_REG262_S1 ( .D(N233), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n236) );
  fd4qd1_hd clk_r_REG261_S1 ( .D(N234), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n346) );
  fd4qd1_hd clk_r_REG260_S1 ( .D(N235), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n235) );
  fd4qd1_hd clk_r_REG259_S1 ( .D(N236), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n234) );
  fd4qd1_hd clk_r_REG258_S1 ( .D(N237), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n233) );
  fd4qd1_hd clk_r_REG257_S1 ( .D(N238), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n232) );
  fd4qd1_hd clk_r_REG256_S1 ( .D(N239), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n345) );
  fd4qd1_hd clk_r_REG253_S1 ( .D(N241), .CK(n926), .SN(1'b1), .RN(n768), .Q(
        n231) );
  fd4qd1_hd clk_r_REG210_S6 ( .D(N662), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n215) );
  fd4qd1_hd clk_r_REG209_S6 ( .D(N661), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n216) );
  fd4qd1_hd clk_r_REG204_S6 ( .D(N664), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n268) );
  fd4qd1_hd clk_r_REG203_S6 ( .D(N663), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n269) );
  fd4qd1_hd clk_r_REG197_S6 ( .D(N653), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n290) );
  fd4qd1_hd clk_r_REG196_S6 ( .D(N652), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n291) );
  fd4qd1_hd clk_r_REG195_S6 ( .D(N651), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n292) );
  fd4qd1_hd clk_r_REG194_S6 ( .D(N650), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n293) );
  fd4qd1_hd clk_r_REG193_S6 ( .D(N649), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n294) );
  fd4qd1_hd clk_r_REG192_S6 ( .D(N648), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n295) );
  fd4qd1_hd clk_r_REG191_S6 ( .D(N647), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n296) );
  fd4qd1_hd clk_r_REG190_S6 ( .D(N646), .CK(n928), .SN(1'b1), .RN(n768), .Q(
        n297) );
  fd4qd1_hd clk_r_REG208_S6 ( .D(N660), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n217) );
  fd4qd1_hd clk_r_REG207_S6 ( .D(N659), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n218) );
  fd4qd1_hd clk_r_REG206_S6 ( .D(N658), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n219) );
  fd4qd1_hd clk_r_REG205_S6 ( .D(N657), .CK(n929), .SN(1'b1), .RN(n768), .Q(
        n220) );
  fd4qd1_hd clk_r_REG202_S6 ( .D(N660), .CK(n931), .SN(1'b1), .RN(n768), .Q(
        n264) );
  fd4qd1_hd clk_r_REG201_S6 ( .D(N659), .CK(n931), .SN(1'b1), .RN(n768), .Q(
        n265) );
  fd4qd1_hd clk_r_REG200_S6 ( .D(N658), .CK(n931), .SN(1'b1), .RN(n768), .Q(
        n266) );
  fd4qd1_hd clk_r_REG199_S6 ( .D(N657), .CK(n931), .SN(1'b1), .RN(n768), .Q(
        n267) );
  fd4qd1_hd clk_r_REG165_S5 ( .D(n934), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        n436) );
  fd4qd1_hd clk_r_REG0_S1 ( .D(n942), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        o_UART_DATA_TX_VALID) );
  fd4qd1_hd clk_r_REG272_S3 ( .D(r_uart_pstate[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n768), .Q(n75) );
  fd4qd1_hd clk_r_REG163_S8 ( .D(n938), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        n461) );
  fd4qd1_hd clk_r_REG150_S5 ( .D(r_mpr_pstate[0]), .CK(i_CLK), .SN(1'b1), .RN(
        n768), .Q(n463) );
  fd4qd1_hd clk_r_REG76_S3 ( .D(N1025), .CK(n930), .SN(1'b1), .RN(n768), .Q(
        n239) );
  fd4qd1_hd clk_r_REG108_S1 ( .D(n941), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        n446) );
  fd4qd1_hd clk_r_REG50_S1 ( .D(n935), .CK(i_CLK), .SN(1'b1), .RN(n768), .Q(
        n445) );
  fd4qd1_hd clk_r_REG159_S5 ( .D(n619), .CK(n930), .SN(1'b1), .RN(n768), .Q(
        o_ADS1292_FILTERED_DATA_ACK) );
  fd4qd1_hd clk_r_REG135_S4 ( .D(r_mpr_pstate[2]), .CK(i_CLK), .SN(1'b1), .RN(
        n768), .Q(n459) );
  fd4qd1_hd clk_r_REG151_S4 ( .D(r_mpr_pstate[1]), .CK(i_CLK), .SN(1'b1), .RN(
        n768), .Q(n464) );
  fd4qd1_hd clk_r_REG134_S3 ( .D(r_mpr_pstate[3]), .CK(i_CLK), .SN(1'b1), .RN(
        n768), .Q(n92) );
  fd4qd2_hd clk_r_REG107_S5 ( .D(r_ads_data_send_ready), .CK(n930), .SN(1'b1), 
        .RN(n636), .Q(n154) );
  ivd1_hd U1 ( .A(1'b1), .Y(o_MPR121_DATA_IN[5]) );
  ivd1_hd U4 ( .A(1'b1), .Y(o_UART_DATA_TX[2]) );
  ivd1_hd U8 ( .A(1'b1), .Y(o_UART_DATA_TX[6]) );
  ivd1_hd U10 ( .A(1'b1), .Y(o_UART_DATA_TX[20]) );
  ivd1_hd U14 ( .A(1'b1), .Y(o_UART_DATA_TX[21]) );
  ivd1_hd U21 ( .A(1'b1), .Y(o_UART_DATA_TX[22]) );
  ivd1_hd U24 ( .A(1'b1), .Y(o_UART_DATA_TX[23]) );
  ivd1_hd U26 ( .A(1'b1), .Y(o_UART_DATA_TX[52]) );
  ivd1_hd U29 ( .A(n338), .Y(N1049) );
  ivd1_hd U35 ( .A(n395), .Y(N1319) );
  ivd1_hd U39 ( .A(o_UART_DATA_TX[49]), .Y(n914) );
  ivd1_hd U46 ( .A(n392), .Y(n93) );
  ivd1_hd U50 ( .A(n436), .Y(N1059) );
  ivd1_hd U55 ( .A(n391), .Y(gt_x_61_n7) );
  nr2d1_hd U58 ( .A(n192), .B(n184), .Y(N251) );
  clknd2d1_hd U339 ( .A(n202), .B(n205), .Y(N1017) );
  nd2bd1_hd U348 ( .AN(r_uart_pstate[1]), .B(n182), .Y(N252) );
  oa21d1_hd U352 ( .A(n392), .B(n94), .C(n95), .Y(N715) );
  mx2d1_hd U467 ( .D0(n445), .D1(n188), .S(N255), .Y(n935) );
  mx2d1_hd U469 ( .D0(n446), .D1(n188), .S(N254), .Y(n941) );
  mx2d1_hd U470 ( .D0(n461), .D1(n948), .S(n949), .Y(n938) );
  mx2d1_hd U472 ( .D0(o_UART_DATA_TX_VALID), .D1(N219), .S(N250), .Y(n942) );
  mx2d1_hd U474 ( .D0(n436), .D1(N700), .S(n524), .Y(n934) );
  mx2d1_hd U482 ( .D0(n391), .D1(N683), .S(N718), .Y(n936) );
  clknd2d1_hd U484 ( .A(n910), .B(N297), .Y(n937) );
  mx2d1_hd U487 ( .D0(n392), .D1(N654), .S(N714), .Y(n940) );
  mx2d1_hd U488 ( .D0(n395), .D1(N316), .S(N333), .Y(n939) );
  mx2d1_hd U491 ( .D0(n338), .D1(N702), .S(n524), .Y(n933) );
  ivd6_hd U499 ( .A(w_rst), .Y(n636) );
  ivd1_hd U624 ( .A(n468), .Y(N298) );
  ivd1_hd U626 ( .A(n906), .Y(n65) );
  ivd1_hd U628 ( .A(n909), .Y(N1087) );
  nd2bd1_hd U630 ( .AN(n909), .B(n62), .Y(n908) );
  clknd2d1_hd U631 ( .A(n2), .B(N63), .Y(n910) );
  clknd2d1_hd U632 ( .A(N277), .B(N276), .Y(n911) );
  ivd1_hd U633 ( .A(n457), .Y(N297) );
  or2d1_hd U634 ( .A(N279), .B(N276), .Y(n912) );
  ivd1_hd U635 ( .A(n914), .Y(o_UART_DATA_TX[7]) );
  ivd1_hd U636 ( .A(n914), .Y(o_UART_DATA_TX[5]) );
  ivd1_hd U637 ( .A(n914), .Y(o_UART_DATA_TX[4]) );
  ivd1_hd U638 ( .A(n914), .Y(o_UART_DATA_TX[3]) );
  ivd1_hd U639 ( .A(n914), .Y(o_UART_DATA_TX[1]) );
  ivd1_hd U640 ( .A(n914), .Y(o_UART_DATA_TX[0]) );
  ivd1_hd U641 ( .A(n914), .Y(o_UART_DATA_TX[55]) );
  nid1_hd U642 ( .A(o_UART_DATA_TX[48]), .Y(o_UART_DATA_TX[54]) );
  or2d1_hd U643 ( .A(n943), .B(n944), .Y(n948) );
  ao211d1_hd U644 ( .A(n78), .B(n945), .C(n347), .D(n946), .Y(n944) );
  ao21d1_hd U645 ( .A(n525), .B(n461), .C(n78), .Y(n946) );
  scg16d1_hd U646 ( .A(n461), .B(n458), .C(n462), .Y(n945) );
  scg21d1_hd U647 ( .A(N274), .B(n180), .C(n461), .D(n78), .Y(n943) );
  nd3d1_hd U648 ( .A(n458), .B(n78), .C(n947), .Y(n949) );
  nr2d1_hd U649 ( .A(n347), .B(n462), .Y(n947) );
  nd2bd1_hd U650 ( .AN(N217), .B(n154), .Y(n961) );
endmodule


module i2c_master_DW01_dec_0 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97;

  xo2d1_hd U35 ( .A(A[16]), .B(n79), .Y(SUM[16]) );
  clknd2d1_hd U36 ( .A(n57), .B(n59), .Y(n55) );
  clknd2d1_hd U37 ( .A(n95), .B(n96), .Y(n92) );
  clknd2d1_hd U38 ( .A(n89), .B(n90), .Y(n86) );
  clknd2d1_hd U39 ( .A(n83), .B(n84), .Y(n80) );
  clknd2d1_hd U40 ( .A(n75), .B(n77), .Y(n73) );
  clknd2d1_hd U41 ( .A(n69), .B(n71), .Y(n67) );
  clknd2d1_hd U42 ( .A(n63), .B(n65), .Y(n61) );
  ao22d1_hd U43 ( .A(A[9]), .B(n54), .C(n55), .D(n56), .Y(SUM[9]) );
  ivd1_hd U44 ( .A(A[9]), .Y(n56) );
  ivd1_hd U45 ( .A(n55), .Y(n54) );
  ao22d1_hd U46 ( .A(A[8]), .B(n57), .C(n58), .D(n59), .Y(SUM[8]) );
  ivd1_hd U47 ( .A(n57), .Y(n58) );
  ao22d1_hd U48 ( .A(A[7]), .B(n60), .C(n61), .D(n62), .Y(SUM[7]) );
  ivd1_hd U49 ( .A(A[7]), .Y(n62) );
  ivd1_hd U50 ( .A(n61), .Y(n60) );
  ao22d1_hd U51 ( .A(A[6]), .B(n63), .C(n64), .D(n65), .Y(SUM[6]) );
  ivd1_hd U52 ( .A(n63), .Y(n64) );
  ao22d1_hd U53 ( .A(A[5]), .B(n66), .C(n67), .D(n68), .Y(SUM[5]) );
  ivd1_hd U54 ( .A(A[5]), .Y(n68) );
  ivd1_hd U55 ( .A(n67), .Y(n66) );
  ao22d1_hd U56 ( .A(A[4]), .B(n69), .C(n70), .D(n71), .Y(SUM[4]) );
  ivd1_hd U57 ( .A(n69), .Y(n70) );
  ao22d1_hd U58 ( .A(A[3]), .B(n72), .C(n73), .D(n74), .Y(SUM[3]) );
  ivd1_hd U59 ( .A(A[3]), .Y(n74) );
  ivd1_hd U60 ( .A(n73), .Y(n72) );
  ao22d1_hd U61 ( .A(A[2]), .B(n75), .C(n76), .D(n77), .Y(SUM[2]) );
  ivd1_hd U62 ( .A(n75), .Y(n76) );
  ao22d1_hd U63 ( .A(A[1]), .B(SUM[0]), .C(A[0]), .D(n78), .Y(SUM[1]) );
  ivd1_hd U64 ( .A(A[1]), .Y(n78) );
  nr2d1_hd U65 ( .A(A[15]), .B(n80), .Y(n79) );
  ao22d1_hd U66 ( .A(A[15]), .B(n81), .C(n80), .D(n82), .Y(SUM[15]) );
  ivd1_hd U67 ( .A(A[15]), .Y(n82) );
  ivd1_hd U68 ( .A(n80), .Y(n81) );
  ao22d1_hd U69 ( .A(A[14]), .B(n83), .C(n85), .D(n84), .Y(SUM[14]) );
  ivd1_hd U70 ( .A(A[14]), .Y(n84) );
  ivd1_hd U71 ( .A(n83), .Y(n85) );
  nr2d1_hd U72 ( .A(A[13]), .B(n86), .Y(n83) );
  ao22d1_hd U73 ( .A(A[13]), .B(n87), .C(n86), .D(n88), .Y(SUM[13]) );
  ivd1_hd U74 ( .A(A[13]), .Y(n88) );
  ivd1_hd U75 ( .A(n86), .Y(n87) );
  ao22d1_hd U76 ( .A(A[12]), .B(n89), .C(n91), .D(n90), .Y(SUM[12]) );
  ivd1_hd U77 ( .A(A[12]), .Y(n90) );
  ivd1_hd U78 ( .A(n89), .Y(n91) );
  nr2d1_hd U79 ( .A(A[11]), .B(n92), .Y(n89) );
  ao22d1_hd U80 ( .A(A[11]), .B(n93), .C(n92), .D(n94), .Y(SUM[11]) );
  ivd1_hd U81 ( .A(A[11]), .Y(n94) );
  ivd1_hd U82 ( .A(n92), .Y(n93) );
  ao22d1_hd U83 ( .A(A[10]), .B(n95), .C(n97), .D(n96), .Y(SUM[10]) );
  ivd1_hd U84 ( .A(A[10]), .Y(n96) );
  ivd1_hd U85 ( .A(n95), .Y(n97) );
  nr2d1_hd U86 ( .A(A[9]), .B(n55), .Y(n95) );
  ivd1_hd U87 ( .A(A[8]), .Y(n59) );
  nr2d1_hd U88 ( .A(A[7]), .B(n61), .Y(n57) );
  ivd1_hd U89 ( .A(A[6]), .Y(n65) );
  nr2d1_hd U90 ( .A(A[5]), .B(n67), .Y(n63) );
  ivd1_hd U91 ( .A(A[4]), .Y(n71) );
  nr2d1_hd U92 ( .A(A[3]), .B(n73), .Y(n69) );
  ivd1_hd U93 ( .A(A[2]), .Y(n77) );
  nr2d1_hd U94 ( .A(A[1]), .B(A[0]), .Y(n75) );
  ivd1_hd U95 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_master_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_master_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_master_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_master_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_master_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module i2c_master ( i_CLK, i_RSTN, cmd_start, cmd_read, cmd_write, 
        cmd_write_multiple, cmd_stop, cmd_valid, cmd_ready, data_in, 
        data_in_valid, data_in_ready, data_in_last, data_out, data_out_valid, 
        data_out_ready, data_out_last, scl_i, scl_o, scl_t, sda_i, sda_o, 
        sda_t, busy, bus_control, bus_active, missed_ack );
  input [7:0] data_in;
  output [7:0] data_out;
  input i_CLK, i_RSTN, cmd_start, cmd_read, cmd_write, cmd_write_multiple,
         cmd_stop, cmd_valid, data_in_valid, data_in_last, data_out_ready,
         scl_i, sda_i;
  output cmd_ready, data_in_ready, data_out_valid, data_out_last, scl_o, scl_t,
         sda_o, sda_t, busy, bus_control, bus_active, missed_ack;
  wire   n271, n272, n281, n283, n284, n285, n287, sda_posedge, sda_negedge,
         last_reg, bit_count_reg_0_, N127, N128, N129, N130, phy_start_bit,
         phy_stop_bit, phy_write_bit, phy_read_bit, N131, N132, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N150, N151,
         N154, N155, N158, N159, N162, N163, N166, N167, N170, N171, N172,
         N173, N174, N175, N178, N179, N182, N183, N229, N232, N249, N255,
         N278, N312, N354, N355, N356, N357, N358, N361, N377, N402, N405,
         N407, N497, N498, N503, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N524,
         N525, N526, N527, N528, N529, N530, N531, N534, N535, N536, N537,
         N538, N539, N542, N543, N546, N547, N550, N551, N552, N553, N554,
         N555, N558, N559, N562, N563, N566, N567, N570, N571, N574, N575,
         N578, N579, N582, N583, N586, N587, N588, N610, N629, N630, N631,
         N632, N693, N696, N699, w_rstn, N701, N907, N908, N911, N913, N914,
         N917, N919, N920, N924, N925, N928, N930, N931, N939, N941, N943,
         N944, N945, N947, N949, N951, N952, N953, N955, N956, N957, N958,
         N960, N961, N962, N963, N965, N966, N967, N968, N969, N970, N971,
         N972, N973, N975, N976, N977, N978, N979, N983, N995, N998, N999,
         N1000, N1001, N1005, N1007, N1013, N1014, N1016, N1017, N1018, N1019,
         N1020, N1021, N1022, N1023, N1024, N1027, N1028, N1029, N1033, N1034,
         N1038, N1039, N1041, N1042, N1043, N1044, N1045, N1046, N1049, N1050,
         N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062,
         N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072,
         N1073, N1074, N1077, N1078, N1079, N1080, N1081, N1082, N1083,
         alt5_n94, alt5_n96, alt5_n97, alt5_n98, alt5_n99, alt5_n100,
         alt5_n101, alt5_n102, alt5_n103, alt5_n104, alt5_n105, alt5_n110,
         alt5_n111, alt5_n112, alt5_n113, alt5_n114, alt5_n115, alt5_n116,
         alt5_n118, alt5_n119, alt5_n120, alt5_n121, alt5_n125, alt5_n126,
         alt5_n127, alt5_n129, alt5_n130, alt5_n131, alt5_n132, alt5_n133,
         alt5_n137, alt5_n138, alt5_n140, alt5_n141, alt5_n142, alt5_n143,
         alt5_n144, alt5_n145, alt5_n146, alt5_n151, alt5_n152, alt5_n153,
         alt5_n154, alt5_n155, alt5_n156, alt5_n157, alt5_n158, alt5_n159,
         alt5_n165, alt5_n166, alt5_n167, alt5_n168, alt5_n169, alt5_n170,
         alt5_n171, alt5_n173, alt5_n174, alt5_n175, alt5_n176, alt5_n177,
         alt5_n178, alt5_n179, alt5_n180, alt5_n181, alt5_n182, alt5_n184,
         alt5_n185, alt5_n186, alt5_n187, alt5_n188, alt5_n189, alt5_n190,
         alt5_n191, alt5_n192, alt5_n193, alt5_n195, alt5_n196, alt5_n197,
         alt5_n198, alt5_n200, alt5_n204, alt5_n207, alt5_n209, alt5_n211,
         alt5_n213, alt5_n215, alt5_n218, alt5_n220, alt5_n221, alt5_n225,
         alt5_n231, alt5_n232, alt5_n233, alt5_n234, alt5_n235, alt5_n236,
         alt5_n237, alt5_n239, alt5_n240, alt5_n241, alt5_n242, alt5_n243,
         alt5_n244, alt5_n245, alt5_n246, alt5_n247, alt5_n248, alt5_n250,
         alt5_n251, alt5_n252, alt5_n253, alt5_n254, alt5_n266, alt5_n267,
         alt5_n269, alt5_n270, alt5_n272, alt5_n278, alt5_n292, alt5_n293,
         alt5_n294, alt5_n370, alt5_n376, alt5_n416, alt5_n417, alt5_n418,
         alt5_n419, alt5_n420, alt5_n421, alt5_n422, alt5_n424, alt5_n425,
         alt5_n426, alt5_n427, alt5_n446, alt5_n492, alt5_n562, gt_x_195_n22,
         gt_x_195_n18, gt_x_195_n17, gt_x_195_n16, gt_x_195_n14, gt_x_195_n13,
         gt_x_195_n12, gt_x_195_n7, gt_x_2_n15, gt_x_2_n9, sub_x_1_n2,
         sub_x_1_n1, n1, n2, n3, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n18, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n41, n43, n45, n46, n47, n48, n49, n50, n51, n53, n54,
         n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n83, n84, n85,
         n86, n87, n88, n90, n91, n94, n95, n98, n100, n103, n106, n109, n112,
         n115, n118, n121, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n139, n142, n144, n145,
         n146, n147, n148, n149, n150, n151, n153, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n181,
         n182, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n223, n227, n228, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n328, n332, n334, n336, n337, n340, n342, n344,
         n347, n348, n349, n350, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n22, n23, n44, n82,
         n89, n92, n107, n108, n110, n113, n114, n116, n117, n119, n120, n122,
         n138, n224, n225, n226, n229, n230, n231, n232, n233, n234, n235,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n266, n267, n268, n269, n270, n404,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n476, n477, n478, n480, n481, n482, n483, n484,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n496, n497,
         n498, n499, n500, n502;
  wire   [7:0] data_reg;
  wire   [3:1] phy_state_reg;
  wire   [16:0] delay_reg;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  oa21d1_hd gt_x_195_U18 ( .A(n117), .B(gt_x_195_n18), .C(gt_x_195_n16), .Y(
        gt_x_195_n14) );
  nr2d1_hd gt_x_195_U17 ( .A(n116), .B(n117), .Y(gt_x_195_n13) );
  ao21d1_hd gt_x_195_U16 ( .A(gt_x_195_n13), .B(n119), .C(gt_x_195_n14), .Y(
        gt_x_195_n12) );
  ivd1_hd gt_x_195_U11 ( .A(n224), .Y(gt_x_195_n7) );
  oa21d1_hd gt_x_195_U4 ( .A(gt_x_195_n12), .B(n224), .C(gt_x_195_n7), .Y(N358) );
  oa21d1_hd gt_x_2_U4 ( .A(n325), .B(n224), .C(gt_x_195_n7), .Y(N357) );
  nd3d1_hd U3 ( .A(n172), .B(N172), .C(n1), .Y(N999) );
  nr3d1_hd U4 ( .A(n310), .B(n332), .C(n318), .Y(n1) );
  nd3d1_hd U5 ( .A(n26), .B(N144), .C(n2), .Y(N995) );
  nr3d1_hd U6 ( .A(n326), .B(N141), .C(n313), .Y(n2) );
  nd3d1_hd U7 ( .A(n3), .B(N552), .C(n5), .Y(N971) );
  scg13d1_hd U9 ( .A(n311), .B(n336), .C(n8), .Y(N966) );
  nd2bd1_hd U10 ( .AN(n315), .B(n6), .Y(N965) );
  scg12d1_hd U11 ( .A(n9), .B(n145), .C(N529), .Y(n6) );
  nr4d1_hd U13 ( .A(n311), .B(n315), .C(n342), .D(n319), .Y(n10) );
  scg13d1_hd U14 ( .A(N529), .B(n334), .C(n11), .Y(N960) );
  nr2bd1_hd U16 ( .AN(n13), .B(n336), .Y(n3) );
  nd3d1_hd U17 ( .A(n9), .B(n12), .C(N552), .Y(N1033) );
  nr2d1_hd U19 ( .A(n228), .B(n314), .Y(n12) );
  ivd1_hd U21 ( .A(n342), .Y(n5) );
  nd4d1_hd U22 ( .A(n9), .B(n15), .C(N536), .D(n16), .Y(N1021) );
  ivd1_hd U24 ( .A(n334), .Y(n15) );
  nr2d1_hd U25 ( .A(n337), .B(n319), .Y(n9) );
  nr3d1_hd U27 ( .A(n342), .B(n320), .C(n314), .Y(n8) );
  ivd1_hd U29 ( .A(n336), .Y(n16) );
  nr4d1_hd U30 ( .A(N553), .B(N537), .C(n337), .D(n315), .Y(n14) );
  nr3d1_hd U32 ( .A(N553), .B(N537), .C(n228), .Y(n11) );
  nr2d1_hd U33 ( .A(n334), .B(n311), .Y(n13) );
  ivd1_hd U35 ( .A(N975), .Y(n18) );
  nr2bd1_hd U57 ( .AN(n24), .B(N132), .Y(phy_write_bit) );
  oa211d1_hd U58 ( .A(n26), .B(n27), .C(n28), .D(n29), .Y(n24) );
  ao21d1_hd U59 ( .A(N312), .B(N128), .C(N130), .Y(n27) );
  scg20d1_hd U60 ( .A(n317), .B(n30), .C(N132), .Y(phy_stop_bit) );
  nr2d1_hd U62 ( .A(n32), .B(N132), .Y(phy_read_bit) );
  nr3d1_hd U63 ( .A(n33), .B(n34), .C(n35), .Y(n32) );
  scg12d1_hd U64 ( .A(N998), .B(n266), .C(n36), .Y(n287) );
  ao22d1_hd U67 ( .A(w_rstn), .B(N977), .C(n41), .D(N973), .Y(n39) );
  oa21d1_hd U70 ( .A(n45), .B(n46), .C(n47), .Y(n284) );
  scg20d1_hd U71 ( .A(sda_t), .B(n48), .C(n43), .Y(n47) );
  ao21d1_hd U72 ( .A(N1020), .B(n41), .C(n49), .Y(n48) );
  ao211d1_hd U73 ( .A(n340), .B(n50), .C(n51), .D(n227), .Y(n46) );
  oa211d1_hd U74 ( .A(sda_t), .B(alt5_n292), .C(n324), .D(n53), .Y(n50) );
  oa211d1_hd U75 ( .A(n54), .B(n55), .C(N693), .D(alt5_n133), .Y(n53) );
  nd4d1_hd U76 ( .A(n57), .B(n58), .C(n59), .D(n60), .Y(n55) );
  nd3d1_hd U77 ( .A(n110), .B(N497), .C(n316), .Y(n58) );
  oa22d1_hd U78 ( .A(alt5_n376), .B(n61), .C(n62), .D(n28), .Y(n54) );
  nr2d1_hd U80 ( .A(n63), .B(n64), .Y(n62) );
  scg4d1_hd U81 ( .A(N1056), .B(n233), .C(N1070), .D(n234), .E(N1060), .F(n231), .G(N1058), .H(n232), .Y(n64) );
  scg4d1_hd U82 ( .A(N1064), .B(n229), .C(N1062), .D(n230), .E(N1068), .F(n225), .G(N1066), .H(n226), .Y(n63) );
  scg7d1_hd U88 ( .A(n37), .B(N960), .C(scl_o), .D(n68), .E(n43), .Y(n283) );
  scg6d1_hd U89 ( .A(N963), .B(n41), .C(n49), .Y(n68) );
  scg14d1_hd U91 ( .A(n70), .B(n71), .C(n72), .Y(n281) );
  oa211d1_hd U92 ( .A(N1001), .B(n73), .C(N131), .D(w_rstn), .Y(n72) );
  ao21d1_hd U94 ( .A(n75), .B(n76), .C(n36), .Y(n272) );
  ivd1_hd U95 ( .A(n77), .Y(n76) );
  ao21d1_hd U96 ( .A(n78), .B(n79), .C(n36), .Y(n271) );
  oa21d1_hd U97 ( .A(N145), .B(n80), .C(n81), .Y(n79) );
  nr2d1_hd U98 ( .A(n26), .B(data_out_valid), .Y(n80) );
  scg22d1_hd U100 ( .A(n120), .B(N503), .C(n43), .D(n83), .Y(alt5_n200) );
  ao22d1_hd U101 ( .A(n37), .B(N969), .C(n120), .D(n84), .Y(n83) );
  ao22d1_hd U104 ( .A(w_rstn), .B(N976), .C(n41), .D(N968), .Y(n85) );
  nr2d1_hd U107 ( .A(n384), .B(n91), .Y(n87) );
  oa21d1_hd U108 ( .A(n359), .B(n91), .C(n94), .Y(delay_reg[15]) );
  ao22d1_hd U109 ( .A(n86), .B(n252), .C(n88), .D(N521), .Y(n94) );
  oa21d1_hd U112 ( .A(n360), .B(n91), .C(n100), .Y(delay_reg[14]) );
  ao22d1_hd U113 ( .A(n86), .B(n251), .C(n88), .D(N520), .Y(n100) );
  oa21d1_hd U116 ( .A(n361), .B(n91), .C(n103), .Y(delay_reg[13]) );
  ao22d1_hd U117 ( .A(n86), .B(n250), .C(n88), .D(N519), .Y(n103) );
  oa21d1_hd U120 ( .A(n362), .B(n91), .C(n106), .Y(delay_reg[12]) );
  ao22d1_hd U121 ( .A(n86), .B(n249), .C(n88), .D(N518), .Y(n106) );
  oa21d1_hd U124 ( .A(n363), .B(n91), .C(n109), .Y(delay_reg[11]) );
  ao22d1_hd U125 ( .A(n86), .B(n248), .C(n88), .D(N517), .Y(n109) );
  oa21d1_hd U128 ( .A(n364), .B(n91), .C(n112), .Y(delay_reg[10]) );
  ao22d1_hd U129 ( .A(n86), .B(n247), .C(n88), .D(N516), .Y(n112) );
  oa21d1_hd U132 ( .A(n365), .B(n91), .C(n115), .Y(delay_reg[9]) );
  ao22d1_hd U133 ( .A(n86), .B(n246), .C(n88), .D(N515), .Y(n115) );
  oa21d1_hd U136 ( .A(n366), .B(n91), .C(n118), .Y(delay_reg[8]) );
  ao22d1_hd U137 ( .A(n86), .B(n245), .C(n88), .D(N514), .Y(n118) );
  oa21d1_hd U140 ( .A(n367), .B(n91), .C(n121), .Y(delay_reg[7]) );
  ao22d1_hd U141 ( .A(n86), .B(n244), .C(n88), .D(N513), .Y(n121) );
  oa21d1_hd U144 ( .A(n123), .B(n91), .C(n124), .Y(delay_reg[6]) );
  ao22d1_hd U145 ( .A(n86), .B(n243), .C(n88), .D(N512), .Y(n124) );
  oa21d1_hd U148 ( .A(n126), .B(n91), .C(n127), .Y(delay_reg[5]) );
  ao22d1_hd U149 ( .A(n86), .B(n242), .C(n88), .D(N511), .Y(n127) );
  oa21d1_hd U152 ( .A(n129), .B(n91), .C(n130), .Y(delay_reg[4]) );
  ao22d1_hd U153 ( .A(n86), .B(n241), .C(n88), .D(N510), .Y(n130) );
  oa21d1_hd U156 ( .A(n132), .B(n91), .C(n133), .Y(delay_reg[3]) );
  ao22d1_hd U157 ( .A(n86), .B(n240), .C(n88), .D(N509), .Y(n133) );
  oa21d1_hd U160 ( .A(n135), .B(n91), .C(n136), .Y(delay_reg[2]) );
  ao22d1_hd U161 ( .A(n86), .B(n239), .C(n88), .D(N508), .Y(n136) );
  oa21d1_hd U164 ( .A(n368), .B(n91), .C(n139), .Y(delay_reg[1]) );
  ao22d1_hd U165 ( .A(n238), .B(n86), .C(n88), .D(N507), .Y(n139) );
  ao21d1_hd U172 ( .A(n138), .B(n237), .C(n270), .Y(delay_reg[0]) );
  nr2d1_hd U174 ( .A(alt5_n370), .B(n384), .Y(n144) );
  nr2d1_hd U177 ( .A(n51), .B(N1024), .Y(n146) );
  ad2d1_hd U178 ( .A(N529), .B(alt5_n272), .Y(n51) );
  nr2bd1_hd U180 ( .AN(n95), .B(alt5_n370), .Y(n147) );
  ao211d1_hd U182 ( .A(N1016), .B(n340), .C(N1023), .D(n149), .Y(n148) );
  nr2bd1_hd U183 ( .AN(N529), .B(alt5_n272), .Y(n149) );
  scg5d1_hd U185 ( .A(n37), .B(N1039), .C(n150), .D(N632), .E(n151), .F(n44), 
        .Y(phy_state_reg[3]) );
  scg5d1_hd U190 ( .A(n37), .B(N1014), .C(n150), .D(N630), .E(n151), .F(n23), 
        .Y(phy_state_reg[1]) );
  nr2d1_hd U192 ( .A(n45), .B(n145), .Y(n150) );
  ivd1_hd U193 ( .A(n340), .Y(n145) );
  ivd1_hd U194 ( .A(n37), .Y(n45) );
  nr2d1_hd U197 ( .A(alt5_n370), .B(n43), .Y(n41) );
  ivd1_hd U198 ( .A(n69), .Y(n151) );
  nd3d1_hd U201 ( .A(n156), .B(n157), .C(n60), .Y(n155) );
  ao211d1_hd U202 ( .A(n312), .B(n108), .C(N173), .D(n33), .Y(n157) );
  ivd1_hd U203 ( .A(n158), .Y(n33) );
  nr4d1_hd U206 ( .A(n162), .B(n163), .C(N983), .D(n164), .Y(n160) );
  oa211d1_hd U208 ( .A(n166), .B(n26), .C(n167), .D(n168), .Y(n165) );
  ao21d1_hd U209 ( .A(bus_active), .B(n169), .C(n77), .Y(n168) );
  ivd1_hd U210 ( .A(n170), .Y(n169) );
  nr4d1_hd U211 ( .A(n171), .B(n35), .C(n163), .D(N1007), .Y(n167) );
  nr2bd1_hd U212 ( .AN(n318), .B(alt5_n446), .Y(n163) );
  nr2d1_hd U213 ( .A(alt5_n492), .B(n172), .Y(n35) );
  ivd1_hd U214 ( .A(n328), .Y(n26) );
  ao211d1_hd U215 ( .A(N128), .B(N978), .C(N979), .D(n173), .Y(n166) );
  nr2d1_hd U216 ( .A(N278), .B(n174), .Y(n173) );
  nd4d1_hd U218 ( .A(n75), .B(n176), .C(n60), .D(n177), .Y(n175) );
  scg6d1_hd U220 ( .A(N128), .B(N129), .C(N130), .Y(n31) );
  nr4d1_hd U221 ( .A(n34), .B(N1005), .C(n178), .D(n179), .Y(n176) );
  oa211d1_hd U222 ( .A(alt5_n562), .B(N144), .C(n29), .D(n181), .Y(n179) );
  ao21d1_hd U224 ( .A(n316), .B(N361), .C(n182), .Y(n29) );
  scg12d1_hd U225 ( .A(N128), .B(N255), .C(N144), .Y(n178) );
  nr2d1_hd U226 ( .A(N358), .B(N172), .Y(n34) );
  ivd1_hd U227 ( .A(n36), .Y(n71) );
  ivd1_hd U231 ( .A(w_rstn), .Y(n43) );
  ivd1_hd U241 ( .A(n57), .Y(n182) );
  nr2d1_hd U243 ( .A(N358), .B(n74), .Y(n70) );
  scg14d1_hd U246 ( .A(n185), .B(data_in_last), .C(n186), .Y(last_reg) );
  oa21d1_hd U247 ( .A(n171), .B(n187), .C(n235), .Y(n186) );
  oa21d1_hd U248 ( .A(n188), .B(n74), .C(n189), .Y(data_reg[7]) );
  ao22d1_hd U249 ( .A(n234), .B(n190), .C(n185), .D(data_in[7]), .Y(n189) );
  oa21d1_hd U250 ( .A(n191), .B(n188), .C(n192), .Y(data_reg[6]) );
  ao22d1_hd U251 ( .A(n232), .B(n312), .C(n185), .D(data_in[6]), .Y(n192) );
  ivd1_hd U252 ( .A(n233), .Y(n188) );
  oa21d1_hd U253 ( .A(n193), .B(n74), .C(n194), .Y(data_reg[5]) );
  ao22d1_hd U254 ( .A(n232), .B(n190), .C(n185), .D(data_in[5]), .Y(n194) );
  oa21d1_hd U255 ( .A(n191), .B(n193), .C(n195), .Y(data_reg[4]) );
  ao22d1_hd U256 ( .A(n230), .B(n312), .C(n185), .D(data_in[4]), .Y(n195) );
  ivd1_hd U257 ( .A(n231), .Y(n193) );
  oa21d1_hd U258 ( .A(n196), .B(n74), .C(n197), .Y(data_reg[3]) );
  ao22d1_hd U259 ( .A(n230), .B(n190), .C(n185), .D(data_in[3]), .Y(n197) );
  oa21d1_hd U260 ( .A(n191), .B(n196), .C(n198), .Y(data_reg[2]) );
  ao22d1_hd U261 ( .A(n226), .B(n312), .C(n185), .D(data_in[2]), .Y(n198) );
  ivd1_hd U262 ( .A(n229), .Y(n196) );
  oa21d1_hd U263 ( .A(n199), .B(n74), .C(n200), .Y(data_reg[1]) );
  ao22d1_hd U264 ( .A(n226), .B(n190), .C(n185), .D(data_in[1]), .Y(n200) );
  ivd1_hd U265 ( .A(n191), .Y(n190) );
  oa21d1_hd U266 ( .A(n191), .B(n199), .C(n201), .Y(data_reg[0]) );
  ao22d1_hd U267 ( .A(n312), .B(n266), .C(n185), .D(data_in[0]), .Y(n201) );
  ivd1_hd U268 ( .A(n225), .Y(n199) );
  ao211d1_hd U269 ( .A(n328), .B(n81), .C(n164), .D(n187), .Y(n191) );
  ivd1_hd U270 ( .A(alt5_n416), .Y(n187) );
  ivd1_hd U271 ( .A(n202), .Y(n81) );
  nd3d1_hd U272 ( .A(n153), .B(n156), .C(n203), .Y(gt_x_2_n9) );
  ao22d1_hd U273 ( .A(n224), .B(n204), .C(N356), .D(n205), .Y(n203) );
  nr4d1_hd U275 ( .A(n326), .B(n332), .C(n310), .D(n208), .Y(n207) );
  ao211d1_hd U276 ( .A(n332), .B(n110), .C(n209), .D(n185), .Y(n156) );
  ad2d1_hd U277 ( .A(N377), .B(n310), .Y(n185) );
  nr2d1_hd U278 ( .A(n210), .B(N278), .Y(n209) );
  ao211d1_hd U279 ( .A(n211), .B(N232), .C(n162), .D(n313), .Y(n153) );
  nr2d1_hd U280 ( .A(bus_active), .B(n170), .Y(n162) );
  nr2d1_hd U281 ( .A(n212), .B(n326), .Y(n170) );
  ivd1_hd U284 ( .A(n214), .Y(n213) );
  ao22ad1_hd U285 ( .A(n119), .B(n214), .C(n205), .D(n119), .Y(
        bit_count_reg_0_) );
  nd3d1_hd U286 ( .A(n172), .B(N172), .C(n74), .Y(n205) );
  ivd1_hd U287 ( .A(n312), .Y(n74) );
  ivd1_hd U289 ( .A(n316), .Y(n172) );
  nr4d1_hd U290 ( .A(n77), .B(n164), .C(n215), .D(n216), .Y(n214) );
  oa21d1_hd U292 ( .A(n326), .B(N141), .C(bus_active), .Y(n217) );
  nd2bd1_hd U294 ( .AN(n210), .B(N278), .Y(n59) );
  ao21d1_hd U296 ( .A(n332), .B(n219), .C(n171), .Y(n75) );
  nr2bd1_hd U297 ( .AN(n310), .B(N377), .Y(n171) );
  ivd1_hd U298 ( .A(n110), .Y(n219) );
  nr2d1_hd U299 ( .A(N232), .B(n161), .Y(n77) );
  ivd1_hd U300 ( .A(n211), .Y(n161) );
  nr2d1_hd U301 ( .A(n174), .B(N144), .Y(n211) );
  nr2d1_hd U314 ( .A(n223), .B(n174), .Y(n208) );
  ivd1_hd U315 ( .A(n177), .Y(n212) );
  nr2d1_hd U318 ( .A(N141), .B(n215), .Y(n206) );
  nd2bd1_hd U320 ( .AN(n215), .B(n78), .Y(n220) );
  oa21d1_hd U323 ( .A(n202), .B(n223), .C(alt5_n416), .Y(n215) );
  nr2d1_hd U324 ( .A(n328), .B(N145), .Y(n223) );
  ao21d1_hd U325 ( .A(N249), .B(N128), .C(N958), .Y(n202) );
  ad2d1_hd U333 ( .A(N953), .B(N957), .Y(N132) );
  nr2d1_hd U335 ( .A(N154), .B(N155), .Y(n313) );
  nr2d1_hd U336 ( .A(N158), .B(N159), .Y(n316) );
  nr2d1_hd U338 ( .A(N582), .B(N583), .Y(n227) );
  nr2d1_hd U339 ( .A(N162), .B(N163), .Y(n332) );
  or2d1_hd U340 ( .A(N127), .B(N129), .Y(N312) );
  or2d1_hd U341 ( .A(phy_stop_bit), .B(alt5_n293), .Y(alt5_n292) );
  or2d1_hd U342 ( .A(phy_read_bit), .B(alt5_n294), .Y(alt5_n293) );
  or2d1_hd U343 ( .A(phy_write_bit), .B(phy_start_bit), .Y(alt5_n294) );
  or2d1_hd U344 ( .A(cmd_read), .B(cmd_write), .Y(N1074) );
  or2d1_hd U345 ( .A(cmd_write), .B(cmd_write_multiple), .Y(N1073) );
  scg2d1_hd U347 ( .A(N407), .B(n318), .C(N145), .D(n31), .Y(n30) );
  ad2d1_hd U348 ( .A(n108), .B(alt5_n446), .Y(N407) );
  ad2d1_hd U349 ( .A(alt5_n272), .B(alt5_n270), .Y(alt5_n269) );
  ivd1_hd U350 ( .A(phy_write_bit), .Y(alt5_n270) );
  ivd1_hd U351 ( .A(phy_start_bit), .Y(alt5_n272) );
  ivd1_hd U352 ( .A(cmd_valid), .Y(N1077) );
  or2d1_hd U353 ( .A(N357), .B(N497), .Y(N361) );
  clknd2d1_hd U354 ( .A(N128), .B(N127), .Y(n174) );
  or2d1_hd U355 ( .A(cmd_start), .B(N949), .Y(N1079) );
  or2d1_hd U357 ( .A(N944), .B(N947), .Y(N949) );
  ad2d1_hd U358 ( .A(N137), .B(N138), .Y(N139) );
  ad2d1_hd U359 ( .A(N917), .B(N911), .Y(N140) );
  clknd2d1_hd U360 ( .A(n238), .B(n98), .Y(n369) );
  ivd1_hd U361 ( .A(alt5_n292), .Y(N610) );
  ad2d1_hd U362 ( .A(phy_stop_bit), .B(alt5_n266), .Y(N699) );
  ad2d1_hd U363 ( .A(alt5_n269), .B(alt5_n267), .Y(alt5_n266) );
  ivd1_hd U364 ( .A(phy_read_bit), .Y(alt5_n267) );
  ad2d1_hd U365 ( .A(phy_read_bit), .B(alt5_n269), .Y(N696) );
  ad2d1_hd U366 ( .A(phy_write_bit), .B(alt5_n272), .Y(N693) );
  clknd2d1_hd U367 ( .A(n75), .B(n59), .Y(n164) );
  or2d1_hd U368 ( .A(N358), .B(N357), .Y(alt5_n492) );
  clknd2d1_hd U369 ( .A(n218), .B(N141), .Y(n177) );
  or2d1_hd U370 ( .A(N127), .B(n358), .Y(N255) );
  clknd2d1_hd U371 ( .A(n328), .B(n31), .Y(n60) );
  clknd2d1_hd U372 ( .A(N141), .B(n174), .Y(n78) );
  or2d1_hd U373 ( .A(N917), .B(n113), .Y(N179) );
  ao21d1_hd U374 ( .A(N976), .B(N506), .C(n147), .Y(n142) );
  or2d1_hd U375 ( .A(n120), .B(N976), .Y(alt5_n198) );
  or2d1_hd U376 ( .A(alt5_n195), .B(alt5_n193), .Y(alt5_n192) );
  ad2d1_hd U377 ( .A(n340), .B(alt5_n197), .Y(alt5_n193) );
  or2d1_hd U378 ( .A(alt5_n198), .B(alt5_n196), .Y(alt5_n195) );
  ad2d1_hd U379 ( .A(N529), .B(alt5_n197), .Y(alt5_n196) );
  or2d1_hd U380 ( .A(alt5_n190), .B(alt5_n189), .Y(alt5_n188) );
  ad2d1_hd U381 ( .A(n319), .B(alt5_n197), .Y(alt5_n189) );
  or2d1_hd U382 ( .A(alt5_n192), .B(alt5_n191), .Y(alt5_n190) );
  ad2d1_hd U383 ( .A(N537), .B(alt5_n197), .Y(alt5_n191) );
  or2d1_hd U384 ( .A(alt5_n186), .B(alt5_n185), .Y(alt5_n184) );
  ad2d1_hd U385 ( .A(n315), .B(alt5_n197), .Y(alt5_n185) );
  or2d1_hd U386 ( .A(alt5_n188), .B(alt5_n187), .Y(alt5_n186) );
  ad2d1_hd U387 ( .A(n337), .B(alt5_n197), .Y(alt5_n187) );
  ad2d1_hd U388 ( .A(gt_x_195_n22), .B(gt_x_195_n18), .Y(N1053) );
  ivd1_hd U389 ( .A(n436), .Y(N944) );
  or2d1_hd U392 ( .A(alt5_n181), .B(alt5_n180), .Y(alt5_n179) );
  ad2d1_hd U393 ( .A(n336), .B(alt5_n197), .Y(alt5_n180) );
  or2d1_hd U394 ( .A(alt5_n184), .B(alt5_n182), .Y(alt5_n181) );
  ad2d1_hd U395 ( .A(N553), .B(alt5_n197), .Y(alt5_n182) );
  or2d1_hd U396 ( .A(N132), .B(alt5_n253), .Y(alt5_n252) );
  ad2d1_hd U397 ( .A(N141), .B(alt5_n254), .Y(alt5_n253) );
  or2d1_hd U398 ( .A(n326), .B(alt5_n426), .Y(alt5_n425) );
  or2d1_hd U399 ( .A(n328), .B(alt5_n427), .Y(alt5_n426) );
  or2d1_hd U400 ( .A(N145), .B(N141), .Y(alt5_n427) );
  ad2d1_hd U403 ( .A(gt_x_195_n22), .B(gt_x_195_n18), .Y(N1069) );
  ad2d1_hd U404 ( .A(gt_x_195_n22), .B(n116), .Y(N1057) );
  ad2d1_hd U405 ( .A(gt_x_195_n22), .B(gt_x_195_n18), .Y(N1061) );
  ad2d1_hd U406 ( .A(gt_x_195_n22), .B(n116), .Y(N1065) );
  ad2d1_hd U407 ( .A(N358), .B(alt5_n376), .Y(N497) );
  or2d1_hd U408 ( .A(N132), .B(alt5_n146), .Y(alt5_n145) );
  ad2d1_hd U409 ( .A(N141), .B(alt5_n221), .Y(alt5_n146) );
  or2d1_hd U411 ( .A(N944), .B(N945), .Y(N947) );
  or2d1_hd U412 ( .A(N944), .B(N944), .Y(N945) );
  or2d1_hd U416 ( .A(N944), .B(N939), .Y(N941) );
  or2d1_hd U417 ( .A(N944), .B(N944), .Y(N939) );
  or2d1_hd U419 ( .A(N917), .B(n113), .Y(N147) );
  or2d1_hd U420 ( .A(alt5_n247), .B(alt5_n246), .Y(alt5_n245) );
  ad2d1_hd U421 ( .A(n326), .B(alt5_n254), .Y(alt5_n246) );
  or2d1_hd U422 ( .A(alt5_n177), .B(alt5_n176), .Y(alt5_n175) );
  ad2d1_hd U423 ( .A(n334), .B(alt5_n197), .Y(alt5_n176) );
  or2d1_hd U424 ( .A(alt5_n179), .B(alt5_n178), .Y(alt5_n177) );
  ad2d1_hd U425 ( .A(n342), .B(alt5_n197), .Y(alt5_n178) );
  ad2d1_hd U426 ( .A(n326), .B(alt5_n221), .Y(alt5_n220) );
  or2d1_hd U427 ( .A(alt5_n250), .B(alt5_n248), .Y(alt5_n247) );
  ad2d1_hd U428 ( .A(n328), .B(alt5_n254), .Y(alt5_n248) );
  or2d1_hd U429 ( .A(alt5_n252), .B(alt5_n251), .Y(alt5_n250) );
  ad2d1_hd U430 ( .A(N145), .B(alt5_n254), .Y(alt5_n251) );
  or2d1_hd U431 ( .A(n310), .B(alt5_n421), .Y(alt5_n420) );
  or2d1_hd U432 ( .A(n332), .B(alt5_n422), .Y(alt5_n421) );
  or2d1_hd U433 ( .A(n316), .B(alt5_n424), .Y(alt5_n422) );
  or2d1_hd U434 ( .A(n313), .B(alt5_n425), .Y(alt5_n424) );
  or4d1_hd U435 ( .A(n311), .B(n314), .C(n228), .D(n227), .Y(N1022) );
  ivd1_hd U436 ( .A(N357), .Y(alt5_n376) );
  clknd2d1_hd U437 ( .A(N358), .B(N173), .Y(n28) );
  clknd2d1_hd U438 ( .A(n316), .B(n65), .Y(n61) );
  or2d1_hd U439 ( .A(N526), .B(N928), .Y(N555) );
  ivd1_hd U440 ( .A(N402), .Y(alt5_n446) );
  ad2d1_hd U441 ( .A(n107), .B(N1081), .Y(N402) );
  ivd1_hd U442 ( .A(n235), .Y(N1081) );
  or2d1_hd U443 ( .A(N130), .B(N128), .Y(alt5_n562) );
  ivd1_hd U444 ( .A(N128), .Y(N958) );
  or2d1_hd U445 ( .A(N142), .B(N143), .Y(N144) );
  or2d1_hd U446 ( .A(n114), .B(N911), .Y(N143) );
  or2d1_hd U447 ( .A(n227), .B(N588), .Y(N967) );
  or2d1_hd U448 ( .A(N526), .B(N928), .Y(N539) );
  clknd2d1_hd U449 ( .A(w_rstn), .B(N975), .Y(n69) );
  or2d1_hd U450 ( .A(N534), .B(N535), .Y(N536) );
  or2d1_hd U451 ( .A(N526), .B(n22), .Y(N535) );
  or2d1_hd U452 ( .A(N526), .B(N928), .Y(N571) );
  or2d1_hd U453 ( .A(N550), .B(N551), .Y(N552) );
  or2d1_hd U454 ( .A(N526), .B(n22), .Y(N551) );
  or2d1_hd U455 ( .A(alt5_n120), .B(alt5_n119), .Y(alt5_n118) );
  ad2d1_hd U456 ( .A(N145), .B(alt5_n133), .Y(alt5_n119) );
  or2d1_hd U457 ( .A(N132), .B(alt5_n121), .Y(alt5_n120) );
  ad2d1_hd U458 ( .A(N141), .B(alt5_n133), .Y(alt5_n121) );
  ad2d1_hd U459 ( .A(n326), .B(alt5_n133), .Y(alt5_n116) );
  or2d1_hd U460 ( .A(alt5_n142), .B(alt5_n218), .Y(alt5_n141) );
  or2d1_hd U461 ( .A(alt5_n143), .B(alt5_n220), .Y(alt5_n142) );
  or2d1_hd U462 ( .A(alt5_n145), .B(alt5_n144), .Y(alt5_n143) );
  ad2d1_hd U463 ( .A(N145), .B(alt5_n221), .Y(alt5_n144) );
  clknd2d1_hd U467 ( .A(n328), .B(n218), .Y(n210) );
  or2d1_hd U468 ( .A(cmd_start), .B(N943), .Y(N1080) );
  or2d1_hd U470 ( .A(N944), .B(N941), .Y(N943) );
  or2d1_hd U471 ( .A(N170), .B(N171), .Y(N172) );
  or2d1_hd U472 ( .A(n114), .B(n113), .Y(N171) );
  or2d1_hd U474 ( .A(alt5_n158), .B(alt5_n215), .Y(alt5_n157) );
  or2d1_hd U475 ( .A(alt5_n159), .B(alt5_n218), .Y(alt5_n158) );
  or2d1_hd U476 ( .A(N132), .B(alt5_n220), .Y(alt5_n159) );
  or2d1_hd U477 ( .A(alt5_n104), .B(alt5_n116), .Y(alt5_n103) );
  or2d1_hd U478 ( .A(alt5_n118), .B(alt5_n105), .Y(alt5_n104) );
  ad2d1_hd U479 ( .A(n328), .B(alt5_n133), .Y(alt5_n105) );
  ad2d1_hd U480 ( .A(n313), .B(alt5_n133), .Y(alt5_n114) );
  ad2d1_hd U481 ( .A(n332), .B(alt5_n133), .Y(alt5_n100) );
  ad2d1_hd U482 ( .A(n316), .B(alt5_n133), .Y(alt5_n132) );
  clknd2d1_hd U483 ( .A(n70), .B(n108), .Y(n57) );
  or2d1_hd U484 ( .A(alt5_n243), .B(alt5_n242), .Y(alt5_n241) );
  ad2d1_hd U485 ( .A(n316), .B(alt5_n254), .Y(alt5_n242) );
  or2d1_hd U486 ( .A(alt5_n245), .B(alt5_n244), .Y(alt5_n243) );
  ad2d1_hd U487 ( .A(n313), .B(alt5_n254), .Y(alt5_n244) );
  nr2d1_hd U488 ( .A(N166), .B(N167), .Y(n310) );
  or2d1_hd U489 ( .A(N917), .B(N911), .Y(N167) );
  or2d1_hd U490 ( .A(alt5_n173), .B(alt5_n171), .Y(alt5_n170) );
  ad2d1_hd U491 ( .A(n320), .B(alt5_n197), .Y(alt5_n171) );
  or2d1_hd U492 ( .A(alt5_n175), .B(alt5_n174), .Y(alt5_n173) );
  ad2d1_hd U493 ( .A(n314), .B(alt5_n197), .Y(alt5_n174) );
  ad2d1_hd U494 ( .A(n316), .B(alt5_n221), .Y(alt5_n215) );
  ad2d1_hd U495 ( .A(n313), .B(alt5_n221), .Y(alt5_n218) );
  ad2d1_hd U497 ( .A(n332), .B(alt5_n221), .Y(alt5_n213) );
  ad2d1_hd U498 ( .A(n310), .B(alt5_n221), .Y(alt5_n211) );
  or2d1_hd U499 ( .A(N917), .B(N911), .Y(N183) );
  ivd1_hd U500 ( .A(N132), .Y(alt5_n133) );
  clknd2d1_hd U501 ( .A(N358), .B(n312), .Y(n158) );
  or2d1_hd U502 ( .A(n312), .B(alt5_n418), .Y(alt5_n417) );
  or2d1_hd U503 ( .A(n318), .B(alt5_n419), .Y(alt5_n418) );
  or2d1_hd U504 ( .A(N173), .B(alt5_n420), .Y(alt5_n419) );
  or2d1_hd U505 ( .A(n114), .B(N913), .Y(N914) );
  or2d1_hd U507 ( .A(N498), .B(n120), .Y(alt5_n370) );
  nr2d1_hd U508 ( .A(n384), .B(n377), .Y(n137) );
  clknd2d1_hd U509 ( .A(n90), .B(n370), .Y(n134) );
  clknd2d1_hd U510 ( .A(n240), .B(n98), .Y(n370) );
  clknd2d1_hd U511 ( .A(n90), .B(n371), .Y(n131) );
  clknd2d1_hd U512 ( .A(n241), .B(n98), .Y(n371) );
  clknd2d1_hd U513 ( .A(n90), .B(n372), .Y(n128) );
  clknd2d1_hd U514 ( .A(n242), .B(n98), .Y(n372) );
  clknd2d1_hd U515 ( .A(n90), .B(n373), .Y(n125) );
  clknd2d1_hd U516 ( .A(n243), .B(n98), .Y(n373) );
  clknd2d1_hd U517 ( .A(n244), .B(n98), .Y(n374) );
  or2d1_hd U519 ( .A(n228), .B(N588), .Y(N1019) );
  clknd2d1_hd U520 ( .A(n14), .B(n16), .Y(N1017) );
  clknd2d1_hd U521 ( .A(n13), .B(n8), .Y(N1018) );
  nr2d1_hd U522 ( .A(N574), .B(N575), .Y(n320) );
  or2d1_hd U523 ( .A(N524), .B(N525), .Y(N574) );
  or2d1_hd U524 ( .A(N526), .B(n22), .Y(N567) );
  clknd2d1_hd U525 ( .A(n14), .B(n5), .Y(N1027) );
  or2d1_hd U526 ( .A(N524), .B(N525), .Y(N582) );
  or2d1_hd U527 ( .A(N526), .B(n22), .Y(N583) );
  or2d1_hd U528 ( .A(n114), .B(N911), .Y(N159) );
  or2d1_hd U529 ( .A(N129), .B(n358), .Y(N978) );
  or2d1_hd U530 ( .A(N130), .B(N229), .Y(N979) );
  ivd1_hd U531 ( .A(alt5_n562), .Y(N229) );
  or2d1_hd U532 ( .A(N917), .B(N911), .Y(N151) );
  or2d1_hd U533 ( .A(n114), .B(n113), .Y(N155) );
  clknd2d1_hd U534 ( .A(n318), .B(N405), .Y(n181) );
  or2d1_hd U535 ( .A(N402), .B(n344), .Y(N405) );
  ivd1_hd U536 ( .A(data_out_ready), .Y(N1078) );
  or2d1_hd U537 ( .A(n317), .B(n187), .Y(N1000) );
  nr2d1_hd U538 ( .A(N578), .B(N579), .Y(n228) );
  or2d1_hd U539 ( .A(N524), .B(N525), .Y(N578) );
  or3d1_hd U542 ( .A(N965), .B(N966), .C(N967), .Y(N968) );
  ad2d1_hd U543 ( .A(N524), .B(N525), .Y(N527) );
  ad2d1_hd U544 ( .A(N526), .B(N928), .Y(N528) );
  clknd2d1_hd U545 ( .A(n145), .B(n10), .Y(N961) );
  or3d1_hd U546 ( .A(n320), .B(n227), .C(N588), .Y(N962) );
  ivd1_hd U548 ( .A(N976), .Y(n376) );
  or3d1_hd U551 ( .A(N970), .B(N971), .C(N972), .Y(N973) );
  or4d1_hd U552 ( .A(n314), .B(n320), .C(n228), .D(n227), .Y(N972) );
  clknd2d1_hd U553 ( .A(n6), .B(N536), .Y(N970) );
  nr2d1_hd U554 ( .A(N174), .B(N175), .Y(n318) );
  or2d1_hd U555 ( .A(n114), .B(N911), .Y(N175) );
  or2d1_hd U556 ( .A(N917), .B(n113), .Y(N163) );
  clknd2d1_hd U557 ( .A(w_rstn), .B(alt5_n133), .Y(n36) );
  or2d1_hd U558 ( .A(alt5_n113), .B(alt5_n132), .Y(alt5_n112) );
  or2d1_hd U559 ( .A(alt5_n115), .B(alt5_n114), .Y(alt5_n113) );
  or2d1_hd U560 ( .A(alt5_n118), .B(alt5_n116), .Y(alt5_n115) );
  or2d1_hd U561 ( .A(alt5_n141), .B(alt5_n132), .Y(alt5_n131) );
  ad2d1_hd U562 ( .A(N173), .B(alt5_n133), .Y(alt5_n130) );
  or2d1_hd U563 ( .A(alt5_n141), .B(alt5_n215), .Y(alt5_n140) );
  or2d1_hd U568 ( .A(sub_x_1_n2), .B(n117), .Y(sub_x_1_n1) );
  clknd2d1_hd U569 ( .A(n78), .B(n217), .Y(n216) );
  or2d1_hd U570 ( .A(alt5_n154), .B(alt5_n207), .Y(alt5_n153) );
  or2d1_hd U571 ( .A(alt5_n155), .B(alt5_n209), .Y(alt5_n154) );
  or2d1_hd U572 ( .A(alt5_n156), .B(alt5_n211), .Y(alt5_n155) );
  or2d1_hd U573 ( .A(alt5_n157), .B(alt5_n213), .Y(alt5_n156) );
  or2d1_hd U574 ( .A(alt5_n99), .B(alt5_n130), .Y(alt5_n98) );
  or2d1_hd U575 ( .A(alt5_n101), .B(alt5_n100), .Y(alt5_n99) );
  or2d1_hd U576 ( .A(alt5_n102), .B(alt5_n132), .Y(alt5_n101) );
  or2d1_hd U577 ( .A(alt5_n103), .B(alt5_n114), .Y(alt5_n102) );
  ad2d1_hd U578 ( .A(n318), .B(alt5_n133), .Y(alt5_n127) );
  ad2d1_hd U579 ( .A(n312), .B(alt5_n133), .Y(alt5_n96) );
  ad2d1_hd U580 ( .A(n317), .B(alt5_n133), .Y(alt5_n125) );
  or2d1_hd U581 ( .A(alt5_n239), .B(alt5_n237), .Y(alt5_n236) );
  ad2d1_hd U582 ( .A(n310), .B(alt5_n254), .Y(alt5_n237) );
  or2d1_hd U583 ( .A(alt5_n241), .B(alt5_n240), .Y(alt5_n239) );
  ad2d1_hd U584 ( .A(n332), .B(alt5_n254), .Y(alt5_n240) );
  ad2d1_hd U585 ( .A(N173), .B(alt5_n254), .Y(alt5_n235) );
  ad2d1_hd U586 ( .A(n318), .B(alt5_n254), .Y(alt5_n233) );
  ad2d1_hd U587 ( .A(n317), .B(alt5_n254), .Y(alt5_n231) );
  ivd1_hd U588 ( .A(alt5_n370), .Y(alt5_n197) );
  ad2d1_hd U589 ( .A(N586), .B(N587), .Y(N588) );
  or2d1_hd U590 ( .A(alt5_n168), .B(alt5_n167), .Y(alt5_n166) );
  ad2d1_hd U591 ( .A(n227), .B(alt5_n197), .Y(alt5_n167) );
  or2d1_hd U592 ( .A(alt5_n170), .B(alt5_n169), .Y(alt5_n168) );
  ad2d1_hd U593 ( .A(n228), .B(alt5_n197), .Y(alt5_n169) );
  ad2d1_hd U598 ( .A(N173), .B(alt5_n221), .Y(alt5_n209) );
  ad2d1_hd U599 ( .A(n318), .B(alt5_n221), .Y(alt5_n207) );
  ad2d1_hd U600 ( .A(n317), .B(alt5_n221), .Y(alt5_n204) );
  clknd2d1_hd U602 ( .A(alt5_n416), .B(n158), .Y(n184) );
  or2d1_hd U604 ( .A(n349), .B(n323), .Y(N1083) );
  or2d1_hd U605 ( .A(n114), .B(N907), .Y(N908) );
  or2d1_hd U606 ( .A(N917), .B(N919), .Y(N920) );
  or2d1_hd U608 ( .A(n22), .B(N952), .Y(N953) );
  or2d1_hd U609 ( .A(N928), .B(N956), .Y(N957) );
  ad2d1_hd U610 ( .A(n268), .B(N1071), .Y(sda_posedge) );
  ad2d1_hd U612 ( .A(N1072), .B(n267), .Y(sda_negedge) );
  scg2d1_hd U613 ( .A(N355), .B(n205), .C(n117), .D(n213), .Y(gt_x_2_n15) );
  xn2d1_hd U614 ( .A(sub_x_1_n2), .B(n117), .Y(N355) );
  scg2d1_hd U615 ( .A(N354), .B(n205), .C(n116), .D(n213), .Y(gt_x_195_n17) );
  nd3d1_hd U616 ( .A(n387), .B(n388), .C(n389), .Y(delay_reg[16]) );
  clknd2d1_hd U617 ( .A(n86), .B(n122), .Y(n389) );
  clknd2d1_hd U618 ( .A(n88), .B(N522), .Y(n388) );
  clknd2d1_hd U619 ( .A(n122), .B(n87), .Y(n387) );
  ad2d1_hd U620 ( .A(n90), .B(n369), .Y(n368) );
  or2d1_hd U621 ( .A(N693), .B(N699), .Y(N631) );
  or2d1_hd U622 ( .A(N1027), .B(N1028), .Y(N1029) );
  or3d1_hd U623 ( .A(N696), .B(N699), .C(N610), .Y(N629) );
  or3d1_hd U624 ( .A(n311), .B(n320), .C(n227), .Y(N1028) );
  or2d1_hd U625 ( .A(N696), .B(N699), .Y(N632) );
  clknd2d1_hd U626 ( .A(n12), .B(n3), .Y(N1038) );
  or2d1_hd U627 ( .A(phy_start_bit), .B(N693), .Y(N630) );
  clknd2d1_hd U628 ( .A(n13), .B(n11), .Y(N1013) );
  clknd2d1_hd U629 ( .A(n160), .B(n161), .Y(n159) );
  or2d1_hd U630 ( .A(n313), .B(n316), .Y(N983) );
  clknd2d1_hd U633 ( .A(alt5_n133), .B(n74), .Y(n73) );
  ad2d1_hd U634 ( .A(data_out_valid), .B(N1078), .Y(N131) );
  ad2d1_hd U635 ( .A(scl_o), .B(N1082), .Y(N503) );
  or4d1_hd U636 ( .A(N537), .B(N553), .C(n334), .D(n228), .Y(N969) );
  scg2d1_hd U637 ( .A(n37), .B(n315), .C(bus_control), .D(n38), .Y(n285) );
  or2d1_hd U640 ( .A(n332), .B(n318), .Y(N998) );
  or2d1_hd U642 ( .A(alt5_n111), .B(alt5_n127), .Y(alt5_n110) );
  or2d1_hd U643 ( .A(alt5_n112), .B(alt5_n130), .Y(alt5_n111) );
  or2d1_hd U645 ( .A(alt5_n129), .B(alt5_n127), .Y(alt5_n126) );
  or2d1_hd U646 ( .A(alt5_n131), .B(alt5_n130), .Y(alt5_n129) );
  or2d1_hd U648 ( .A(alt5_n138), .B(alt5_n207), .Y(alt5_n137) );
  or2d1_hd U649 ( .A(alt5_n140), .B(alt5_n209), .Y(alt5_n138) );
  xn2d1_hd U656 ( .A(sub_x_1_n1), .B(n224), .Y(N356) );
  clknd2d1_hd U657 ( .A(n206), .B(n207), .Y(n204) );
  or2d1_hd U659 ( .A(N132), .B(alt5_n233), .Y(alt5_n225) );
  or2d1_hd U661 ( .A(alt5_n153), .B(alt5_n152), .Y(alt5_n151) );
  ad2d1_hd U662 ( .A(n312), .B(alt5_n221), .Y(alt5_n152) );
  or2d1_hd U664 ( .A(alt5_n97), .B(alt5_n96), .Y(alt5_n94) );
  or2d1_hd U665 ( .A(alt5_n98), .B(alt5_n127), .Y(alt5_n97) );
  or2d1_hd U674 ( .A(alt5_n234), .B(alt5_n233), .Y(alt5_n232) );
  or2d1_hd U675 ( .A(alt5_n236), .B(alt5_n235), .Y(alt5_n234) );
  ad2d1_hd U679 ( .A(N588), .B(alt5_n197), .Y(alt5_n165) );
  or2d1_hd U686 ( .A(n350), .B(n322), .Y(N701) );
  xn2d1_hd U689 ( .A(n119), .B(n116), .Y(N354) );
  or2d1_hd U690 ( .A(n119), .B(n116), .Y(sub_x_1_n2) );
  ad2d1_hd U691 ( .A(n119), .B(n116), .Y(N1049) );
  ad2d1_hd U692 ( .A(n119), .B(gt_x_195_n18), .Y(N1067) );
  ad2d1_hd U693 ( .A(n119), .B(n116), .Y(N1063) );
  ad2d1_hd U694 ( .A(n119), .B(gt_x_195_n18), .Y(N1059) );
  ad2d1_hd U695 ( .A(n119), .B(n116), .Y(N1055) );
  ad2d1_hd U696 ( .A(n119), .B(gt_x_195_n18), .Y(N1045) );
  ivd1_hd U697 ( .A(n119), .Y(gt_x_195_n22) );
  nr2bd2_hd U698 ( .AN(n120), .B(n43), .Y(n86) );
  ivd1_hd U699 ( .A(n117), .Y(gt_x_195_n16) );
  ivd2_hd U700 ( .A(n41), .Y(n91) );
  or2d1_hd U705 ( .A(n92), .B(N138), .Y(N166) );
  or2d1_hd U706 ( .A(n92), .B(N138), .Y(N162) );
  or2d1_hd U707 ( .A(n92), .B(N138), .Y(N154) );
  or2d1_hd U708 ( .A(n92), .B(N138), .Y(N158) );
  or2d1_hd U710 ( .A(n89), .B(n92), .Y(N919) );
  or2d1_hd U711 ( .A(n89), .B(n92), .Y(N907) );
  or2d1_hd U712 ( .A(n89), .B(n92), .Y(N913) );
  or2d1_hd U713 ( .A(N137), .B(n89), .Y(N182) );
  or2d1_hd U714 ( .A(N137), .B(n89), .Y(N174) );
  or2d1_hd U715 ( .A(n92), .B(n89), .Y(N142) );
  or2d1_hd U716 ( .A(N137), .B(n89), .Y(N170) );
  or2d1_hd U717 ( .A(n92), .B(n89), .Y(N146) );
  or2d1_hd U718 ( .A(n92), .B(n89), .Y(N150) );
  or2d1_hd U719 ( .A(N137), .B(n89), .Y(N178) );
  nr2d1_hd U720 ( .A(n95), .B(n125), .Y(n123) );
  nr2d1_hd U721 ( .A(n95), .B(n128), .Y(n126) );
  nr2d1_hd U722 ( .A(n95), .B(n131), .Y(n129) );
  nr2d1_hd U723 ( .A(n95), .B(n134), .Y(n132) );
  nr2d1_hd U724 ( .A(n95), .B(n137), .Y(n135) );
  or2d1_hd U725 ( .A(n23), .B(N930), .Y(N931) );
  or2d1_hd U726 ( .A(n23), .B(N924), .Y(N925) );
  ad2d1_hd U727 ( .A(n23), .B(n22), .Y(N587) );
  or2d1_hd U728 ( .A(n23), .B(n22), .Y(N559) );
  or2d1_hd U729 ( .A(n23), .B(N928), .Y(N579) );
  or2d1_hd U730 ( .A(n23), .B(N928), .Y(N547) );
  or2d1_hd U731 ( .A(n23), .B(n22), .Y(N575) );
  or2d1_hd U732 ( .A(n23), .B(n22), .Y(N543) );
  or2d1_hd U733 ( .A(n23), .B(N928), .Y(N531) );
  or2d1_hd U734 ( .A(n23), .B(N928), .Y(N563) );
  or2d1_hd U735 ( .A(n23), .B(N951), .Y(N952) );
  or2d1_hd U736 ( .A(n23), .B(N955), .Y(N956) );
  or2d1_hd U741 ( .A(n44), .B(N525), .Y(N550) );
  or2d1_hd U742 ( .A(n44), .B(N525), .Y(N546) );
  or2d1_hd U743 ( .A(n44), .B(N525), .Y(N542) );
  or2d1_hd U744 ( .A(n44), .B(N525), .Y(N554) );
  or2d1_hd U746 ( .A(n82), .B(n44), .Y(N930) );
  or2d1_hd U747 ( .A(n82), .B(n44), .Y(N924) );
  ad2d1_hd U748 ( .A(n44), .B(n82), .Y(N586) );
  or2d1_hd U749 ( .A(N524), .B(n82), .Y(N558) );
  or2d1_hd U750 ( .A(n44), .B(n82), .Y(N538) );
  or2d1_hd U751 ( .A(N524), .B(n82), .Y(N566) );
  or2d1_hd U752 ( .A(n44), .B(n82), .Y(N534) );
  or2d1_hd U753 ( .A(N524), .B(n82), .Y(N562) );
  or2d1_hd U754 ( .A(n44), .B(n82), .Y(N530) );
  or2d1_hd U755 ( .A(N524), .B(n82), .Y(N570) );
  or2d1_hd U756 ( .A(n82), .B(n44), .Y(N951) );
  or2d1_hd U757 ( .A(n82), .B(n44), .Y(N955) );
  nr2bd2_hd U758 ( .AN(N976), .B(n43), .Y(n88) );
  ad2d1_hd U759 ( .A(N498), .B(alt5_n278), .Y(N976) );
  ivd1_hd U760 ( .A(n116), .Y(gt_x_195_n18) );
  ad2d1_hd U761 ( .A(gt_x_195_n22), .B(n116), .Y(N1043) );
  ad2d1_hd U762 ( .A(n119), .B(n116), .Y(N1041) );
  nr2d1_hd U841 ( .A(N566), .B(N567), .Y(n311) );
  ad2d1_hd U842 ( .A(N1043), .B(n117), .Y(N1044) );
  ad2d1_hd U843 ( .A(N1057), .B(n117), .Y(N1058) );
  ad2d1_hd U844 ( .A(N1061), .B(n117), .Y(N1062) );
  nr2d1_hd U846 ( .A(N570), .B(N571), .Y(n314) );
  nr2d1_hd U847 ( .A(N546), .B(N547), .Y(n315) );
  ad2d1_hd U848 ( .A(N1041), .B(n117), .Y(N1042) );
  ad2d1_hd U849 ( .A(N1059), .B(n117), .Y(N1060) );
  ad2d1_hd U850 ( .A(N1065), .B(gt_x_195_n16), .Y(N1066) );
  or2d1_hd U851 ( .A(N1079), .B(cmd_read), .Y(N232) );
  ad2d1_hd U852 ( .A(cmd_ready), .B(N1077), .Y(N130) );
  ad2d1_hd U853 ( .A(data_in_ready), .B(data_in_valid), .Y(N377) );
  ad2d1_hd U854 ( .A(N139), .B(N140), .Y(N141) );
  nr2d1_hd U855 ( .A(N182), .B(N183), .Y(n317) );
  ad2d1_hd U856 ( .A(N527), .B(N528), .Y(N529) );
  nr2d1_hd U857 ( .A(N538), .B(N539), .Y(n319) );
  ad2d1_hd U858 ( .A(N1045), .B(n117), .Y(N1046) );
  ad2d1_hd U859 ( .A(N1069), .B(gt_x_195_n16), .Y(N1070) );
  ad2d1_hd U861 ( .A(N1063), .B(gt_x_195_n16), .Y(N1064) );
  nr2d1_hd U862 ( .A(N928), .B(N931), .Y(n321) );
  nr2d1_hd U863 ( .A(n348), .B(n321), .Y(n322) );
  nr2d1_hd U864 ( .A(N911), .B(N914), .Y(n323) );
  nr2d1_hd U865 ( .A(phy_start_bit), .B(N696), .Y(n324) );
  scg9d1_hd U866 ( .A(n117), .B(gt_x_195_n18), .C(gt_x_195_n16), .Y(n325) );
  or2d1_hd U867 ( .A(N1080), .B(cmd_write), .Y(N278) );
  ad2d1_hd U868 ( .A(cmd_ready), .B(cmd_valid), .Y(N128) );
  nr2d1_hd U869 ( .A(N150), .B(N151), .Y(n326) );
  ivd1_hd U870 ( .A(N144), .Y(N145) );
  ivd1_hd U871 ( .A(N172), .Y(N173) );
  nr2d1_hd U872 ( .A(N146), .B(N147), .Y(n328) );
  ivd1_hd U876 ( .A(N536), .Y(N537) );
  nr2d1_hd U878 ( .A(N562), .B(N563), .Y(n334) );
  nr2d1_hd U880 ( .A(N554), .B(N555), .Y(n336) );
  nr2d1_hd U881 ( .A(N542), .B(N543), .Y(n337) );
  nr2d1_hd U884 ( .A(N530), .B(N531), .Y(n340) );
  or2d1_hd U885 ( .A(n317), .B(alt5_n417), .Y(alt5_n416) );
  or3d1_hd U887 ( .A(N995), .B(N999), .C(N1000), .Y(N1001) );
  or2d1_hd U888 ( .A(N1021), .B(N1022), .Y(N1023) );
  ad2d1_hd U889 ( .A(N1053), .B(gt_x_195_n16), .Y(N1054) );
  ivd1_hd U891 ( .A(N552), .Y(N553) );
  nr2d1_hd U892 ( .A(N558), .B(N559), .Y(n342) );
  nr2d1_hd U894 ( .A(n108), .B(N402), .Y(n344) );
  or2d1_hd U895 ( .A(n332), .B(n312), .Y(N1007) );
  or2d1_hd U896 ( .A(n326), .B(n313), .Y(N1005) );
  or3d1_hd U897 ( .A(N1017), .B(N1018), .C(N1019), .Y(N1020) );
  or4d1_hd U898 ( .A(n315), .B(n342), .C(n320), .D(N588), .Y(N1024) );
  ad2d1_hd U900 ( .A(N1055), .B(n117), .Y(N1056) );
  or2d1_hd U901 ( .A(N1033), .B(n227), .Y(N1034) );
  or2d1_hd U902 ( .A(N961), .B(N962), .Y(N963) );
  ad2d1_hd U903 ( .A(N1049), .B(gt_x_195_n16), .Y(N1050) );
  or2d1_hd U904 ( .A(N1013), .B(n227), .Y(N1014) );
  or2d1_hd U905 ( .A(N1038), .B(n227), .Y(N1039) );
  ad2d1_hd U906 ( .A(N1067), .B(gt_x_195_n16), .Y(N1068) );
  nr2d1_hd U909 ( .A(n113), .B(N920), .Y(n347) );
  nr2d1_hd U910 ( .A(n22), .B(N925), .Y(n348) );
  nr2d1_hd U911 ( .A(n113), .B(N908), .Y(n349) );
  nr2d1_hd U913 ( .A(N1083), .B(n347), .Y(n350) );
  nid1_hd U914 ( .A(scl_o), .Y(scl_t) );
  nr4d1_hd U915 ( .A(n245), .B(n243), .C(n242), .D(n241), .Y(n356) );
  nr4d1_hd U916 ( .A(n240), .B(n239), .C(n238), .D(n122), .Y(n355) );
  nr4d1_hd U917 ( .A(n252), .B(n251), .C(n250), .D(n249), .Y(n354) );
  or4d1_hd U918 ( .A(n247), .B(delay_reg[0]), .C(n244), .D(n246), .Y(n352) );
  nr2d1_hd U919 ( .A(n248), .B(n352), .Y(n353) );
  nd4d1_hd U920 ( .A(n356), .B(n355), .C(n354), .D(n353), .Y(N498) );
  nr2d1_hd U921 ( .A(N1074), .B(cmd_write_multiple), .Y(n357) );
  ad2d1_hd U922 ( .A(cmd_stop), .B(n357), .Y(N129) );
  nr2d1_hd U923 ( .A(N129), .B(N127), .Y(n358) );
  ivd1_hd U924 ( .A(N127), .Y(N249) );
  xo2d1_hd U925 ( .A(cmd_read), .B(N1073), .Y(N127) );
  or4d1_hd U926 ( .A(phy_start_bit), .B(N693), .C(N696), .D(N699), .Y(N1016)
         );
  or2d1_hd U927 ( .A(n384), .B(n386), .Y(n359) );
  or2d1_hd U928 ( .A(n384), .B(n385), .Y(n360) );
  or2d1_hd U929 ( .A(n384), .B(n383), .Y(n361) );
  ivd1_hd U930 ( .A(n98), .Y(n384) );
  or2d1_hd U931 ( .A(n384), .B(n382), .Y(n362) );
  or2d1_hd U932 ( .A(n384), .B(n381), .Y(n363) );
  or2d1_hd U933 ( .A(n384), .B(n380), .Y(n364) );
  or2d1_hd U934 ( .A(n384), .B(n379), .Y(n365) );
  or2d1_hd U935 ( .A(n384), .B(n378), .Y(n366) );
  ad2d1_hd U936 ( .A(n90), .B(n374), .Y(n367) );
  ad2d1_hd u_cell_6241 ( .A(N701), .B(w_rstn), .Y(n404) );
  fd3qd1_hd clk_r_REG28_S5 ( .D(n404), .CK(i_CLK), .SN(1'b1), .Q(busy) );
  fd1eqd1_hd clk_r_REG31_S6 ( .D(last_reg), .E(n430), .CK(n439), .Q(n235) );
  fd1eqd1_hd clk_r_REG73_S2 ( .D(n268), .E(n431), .CK(n440), .Q(n266) );
  fd1eqd1_hd clk_r_REG57_S8 ( .D(bit_count_reg_0_), .E(n435), .CK(n439), .Q(
        n119) );
  fd1eqd1_hd clk_r_REG52_S1 ( .D(gt_x_2_n9), .E(n435), .CK(n439), .Q(n224) );
  fd1eqd1_hd clk_r_REG49_S8 ( .D(data_reg[0]), .E(n434), .CK(n439), .Q(n225)
         );
  fd1eqd1_hd clk_r_REG43_S8 ( .D(data_reg[2]), .E(n434), .CK(n439), .Q(n229)
         );
  fd1eqd1_hd clk_r_REG39_S8 ( .D(data_reg[4]), .E(n429), .CK(n439), .Q(n231)
         );
  fd1eqd1_hd clk_r_REG36_S8 ( .D(data_reg[6]), .E(n428), .CK(n439), .Q(n233)
         );
  fd1eqd1_hd clk_r_REG58_S8 ( .D(gt_x_195_n17), .E(n435), .CK(n439), .Q(n116)
         );
  fd1eqd1_hd clk_r_REG51_S8 ( .D(gt_x_2_n15), .E(n435), .CK(n439), .Q(n117) );
  fd1eqd1_hd clk_r_REG47_S6 ( .D(data_reg[1]), .E(n434), .CK(n439), .Q(n226)
         );
  fd1eqd1_hd clk_r_REG44_S9 ( .D(data_reg[3]), .E(n434), .CK(n439), .Q(n230)
         );
  fd1eqd1_hd clk_r_REG40_S9 ( .D(data_reg[5]), .E(n428), .CK(n439), .Q(n232)
         );
  fd1eqd1_hd clk_r_REG37_S9 ( .D(data_reg[7]), .E(n428), .CK(n439), .Q(n234)
         );
  fd3d1_hd clk_r_REG1_S2 ( .D(alt5_n200), .CK(n441), .SN(1'b1), .Q(n120), .QN(
        alt5_n278) );
  fd3d1_hd clk_r_REG72_S1 ( .D(sda_i), .CK(i_CLK), .SN(1'b1), .Q(n268), .QN(
        N1072) );
  fd3d1_hd clk_r_REG70_S1 ( .D(scl_i), .CK(i_CLK), .SN(1'b1), .Q(n269), .QN(
        N1082) );
  fd3d1_hd clk_r_REG53_S6 ( .D(n481), .CK(n439), .SN(1'b1), .Q(n113), .QN(N911) );
  fd3d1_hd clk_r_REG35_S6 ( .D(n482), .CK(n439), .SN(1'b1), .Q(n92), .QN(N137)
         );
  fd3d1_hd clk_r_REG54_S1 ( .D(n483), .CK(n439), .SN(1'b1), .Q(n114), .QN(N917) );
  fd3d1_hd clk_r_REG32_S7 ( .D(n484), .CK(n439), .SN(1'b1), .Q(n89), .QN(N138)
         );
  fd3d1_hd clk_r_REG27_S4 ( .D(phy_state_reg[1]), .CK(n440), .SN(1'b1), .Q(n23), .QN(N526) );
  fd3d1_hd clk_r_REG24_S4 ( .D(phy_state_reg[3]), .CK(n440), .SN(1'b1), .Q(n44), .QN(N524) );
  fd3d1_hd clk_r_REG5_S4 ( .D(n284), .CK(n440), .SN(1'b1), .Q(sda_o), .QN(
        sda_t) );
  fd3d1_hd clk_r_REG25_S4 ( .D(n477), .CK(n440), .SN(1'b1), .Q(n22), .QN(N928)
         );
  fd3d1_hd clk_r_REG0_S1 ( .D(n478), .CK(n440), .SN(1'b1), .Q(n82), .QN(N525)
         );
  fd3d1_hd clk_r_REG18_S5 ( .D(delay_reg[8]), .CK(n441), .SN(1'b1), .Q(n245), 
        .QN(n378) );
  fd3d1_hd clk_r_REG17_S5 ( .D(delay_reg[10]), .CK(n441), .SN(1'b1), .Q(n247), 
        .QN(n380) );
  fd3d1_hd clk_r_REG16_S5 ( .D(delay_reg[11]), .CK(n441), .SN(1'b1), .Q(n248), 
        .QN(n381) );
  fd3d1_hd clk_r_REG15_S5 ( .D(delay_reg[12]), .CK(n441), .SN(1'b1), .Q(n249), 
        .QN(n382) );
  fd3d1_hd clk_r_REG14_S5 ( .D(delay_reg[13]), .CK(n441), .SN(1'b1), .Q(n250), 
        .QN(n383) );
  fd3d1_hd clk_r_REG13_S5 ( .D(delay_reg[14]), .CK(n441), .SN(1'b1), .Q(n251), 
        .QN(n385) );
  fd3d1_hd clk_r_REG12_S5 ( .D(delay_reg[15]), .CK(n441), .SN(1'b1), .Q(n252), 
        .QN(n386) );
  fd3d1_hd clk_r_REG10_S5 ( .D(delay_reg[9]), .CK(n441), .SN(1'b1), .Q(n246), 
        .QN(n379) );
  fd3d1_hd clk_r_REG22_S4 ( .D(delay_reg[2]), .CK(n441), .SN(1'b1), .Q(n239), 
        .QN(n377) );
  fd1qd1_hd clk_r_REG59_S7 ( .D(n500), .CK(n437), .Q(n110) );
  fd1qd1_hd clk_r_REG60_S7 ( .D(n499), .CK(n437), .Q(n108) );
  fd1qd1_hd clk_r_REG61_S7 ( .D(n498), .CK(n437), .Q(n107) );
  fd1qd1_hd clk_r_REG38_S9 ( .D(n494), .CK(n438), .Q(data_out[7]) );
  fd1qd1_hd clk_r_REG41_S10 ( .D(n493), .CK(n438), .Q(data_out[6]) );
  fd1qd1_hd clk_r_REG42_S9 ( .D(n492), .CK(n438), .Q(data_out[5]) );
  fd1qd1_hd clk_r_REG45_S10 ( .D(n491), .CK(n438), .Q(data_out[4]) );
  fd1qd1_hd clk_r_REG46_S9 ( .D(n490), .CK(n438), .Q(data_out[3]) );
  fd1qd1_hd clk_r_REG48_S7 ( .D(n489), .CK(n438), .Q(data_out[2]) );
  fd1qd1_hd clk_r_REG50_S9 ( .D(n488), .CK(n438), .Q(data_out[1]) );
  fd1qd1_hd clk_r_REG55_S2 ( .D(n182), .CK(n438), .Q(data_out_last) );
  fd1qd1_hd clk_r_REG56_S2 ( .D(n487), .CK(n438), .Q(data_out[0]) );
  i2c_master_DW01_dec_0 sub_x_144 ( .A({n122, n252, n251, n250, n249, n248, 
        n247, n246, n245, n244, n243, n242, n241, n240, n239, n238, 
        delay_reg[0]}), .SUM({N522, N521, N520, N519, N518, N517, N516, N515, 
        N514, N513, N512, N511, N510, N509, N508, N507, N506}) );
  SNPS_CLOCK_GATE_HIGH_i2c_master_8 clk_gate_clk_r_REG9_S5_0 ( .CLK(i_CLK), 
        .EN(n476), .ENCLK(n441), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_master_9 clk_gate_clk_r_REG0_S1_0 ( .CLK(i_CLK), 
        .EN(n480), .ENCLK(n440), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_master_10 clk_gate_clk_r_REG32_S7_0 ( .CLK(i_CLK), 
        .EN(n486), .ENCLK(n439), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_master_11 clk_gate_clk_r_REG38_S9_0 ( .CLK(i_CLK), 
        .EN(n496), .ENCLK(n438), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_master_12 clk_gate_clk_r_REG59_S7_0 ( .CLK(i_CLK), 
        .EN(n502), .ENCLK(n437), .TE(1'b0) );
  fd1qd1_hd R_0_clk_r_REG65_S7 ( .D(n497), .CK(n437), .Q(n436) );
  fd3qd1_hd clk_r_REG74_S2 ( .D(n268), .CK(i_CLK), .SN(1'b1), .Q(n267) );
  fd3qd1_hd clk_r_REG29_S5 ( .D(n287), .CK(i_CLK), .SN(1'b1), .Q(missed_ack)
         );
  fd3qd1_hd clk_r_REG23_S4 ( .D(n283), .CK(n440), .SN(1'b1), .Q(scl_o) );
  fd3qd1_hd clk_r_REG4_S4 ( .D(n285), .CK(n441), .SN(1'b1), .Q(bus_control) );
  fd3qd1_hd clk_r_REG33_S8 ( .D(n281), .CK(i_CLK), .SN(1'b1), .Q(
        data_out_valid) );
  fd3qd1_hd clk_r_REG34_S5 ( .D(n271), .CK(i_CLK), .SN(1'b1), .Q(cmd_ready) );
  fd3qd1_hd clk_r_REG30_S5 ( .D(n272), .CK(i_CLK), .SN(1'b1), .Q(data_in_ready) );
  fd3qd1_hd clk_r_REG9_S5 ( .D(delay_reg[7]), .CK(n441), .SN(1'b1), .Q(n244)
         );
  fd3qd1_hd clk_r_REG26_S5 ( .D(delay_reg[1]), .CK(n441), .SN(1'b1), .Q(n238)
         );
  fd3qd1_hd clk_r_REG11_S5 ( .D(delay_reg[16]), .CK(n441), .SN(1'b1), .Q(n122)
         );
  fd3qd1_hd clk_r_REG21_S4 ( .D(delay_reg[3]), .CK(n441), .SN(1'b1), .Q(n240)
         );
  fd3qd1_hd clk_r_REG20_S4 ( .D(delay_reg[4]), .CK(n441), .SN(1'b1), .Q(n241)
         );
  fd3qd1_hd clk_r_REG19_S4 ( .D(delay_reg[5]), .CK(n441), .SN(1'b1), .Q(n242)
         );
  fd3qd1_hd clk_r_REG8_S4 ( .D(delay_reg[6]), .CK(n441), .SN(1'b1), .Q(n243)
         );
  fds2eqd1_hd clk_r_REG71_S2 ( .CRN(1'b1), .D(n473), .E(n474), .CK(i_CLK), .Q(
        bus_active) );
  fds2eqd1_hd clk_r_REG3_S4 ( .CRN(1'b1), .D(n470), .E(n471), .CK(i_CLK), .Q(
        n237) );
  fd3qd1_hd clk_r_REG75_S1 ( .D(n43), .CK(i_CLK), .SN(1'b1), .Q(n270) );
  fd3qd1_hd clk_r_REG2_S3 ( .D(n142), .CK(i_CLK), .SN(1'b1), .Q(n138) );
  or3d1_hd U607 ( .A(n120), .B(1'b0), .C(N976), .Y(N975) );
  scg4d1_hd U86 ( .A(N1042), .B(1'b0), .C(N1054), .D(n436), .E(N1046), .F(n436), .G(N1044), .H(n436), .Y(n66) );
  nr2d1_hd U181 ( .A(1'b0), .B(n148), .Y(n95) );
  nr2d1_hd U195 ( .A(n91), .B(1'b0), .Y(n37) );
  clknd2d1_hd U518 ( .A(N553), .B(1'b1), .Y(n90) );
  clknd2d1_hd U540 ( .A(n85), .B(1'b1), .Y(n84) );
  clknd2d1_hd U547 ( .A(1'b1), .B(n69), .Y(n49) );
  clknd2d1_hd U638 ( .A(n39), .B(1'b1), .Y(n38) );
  nd3d1_hd U639 ( .A(1'b1), .B(alt5_n278), .C(n376), .Y(N977) );
  ad2d1_hd U332 ( .A(1'b1), .B(alt5_n133), .Y(alt5_n221) );
  ad2d1_hd U334 ( .A(1'b1), .B(alt5_n133), .Y(alt5_n254) );
  scg17d1_hd U84 ( .A(N1050), .B(n436), .C(n66), .D(1'b1), .Y(n65) );
  ivd2_hd U1 ( .A(n174), .Y(n218) );
  nr2d1_hd U2 ( .A(n153), .B(N132), .Y(phy_start_bit) );
  oa211d1_hd U8 ( .A(n443), .B(1'b1), .C(n445), .D(w_rstn), .Y(n476) );
  clknd2d1_hd U12 ( .A(n446), .B(1'b1), .Y(n445) );
  ao211d1_hd U15 ( .A(n22), .B(n458), .C(1'b0), .D(n120), .Y(n447) );
  oa21d2_hd U18 ( .A(alt5_n292), .B(n145), .C(n146), .Y(n98) );
  clknd2d1_hd U23 ( .A(N524), .B(N928), .Y(n460) );
  clknd2d1_hd U41 ( .A(n23), .B(n82), .Y(n461) );
  clknd2d1_hd U42 ( .A(alt5_n278), .B(n457), .Y(n462) );
  clknd2d1_hd U51 ( .A(n37), .B(N1029), .Y(n463) );
  nr2d2_hd U52 ( .A(N178), .B(N179), .Y(n312) );
  ivd1_hd U111 ( .A(n267), .Y(N1071) );
  or2d1_hd U115 ( .A(n212), .B(n208), .Y(n427) );
  nr2d1_hd U118 ( .A(alt5_n137), .B(alt5_n204), .Y(n428) );
  nr2d1_hd U119 ( .A(alt5_n126), .B(alt5_n125), .Y(n429) );
  nr2d1_hd U122 ( .A(alt5_n94), .B(alt5_n125), .Y(n430) );
  nr2d1_hd U123 ( .A(alt5_n166), .B(alt5_n165), .Y(n431) );
  nr2d1_hd U126 ( .A(alt5_n232), .B(alt5_n231), .Y(n432) );
  nr2d1_hd U127 ( .A(alt5_n151), .B(alt5_n204), .Y(n433) );
  nr2d1_hd U130 ( .A(alt5_n110), .B(alt5_n125), .Y(n434) );
  nr2d1_hd U131 ( .A(alt5_n225), .B(alt5_n231), .Y(n435) );
  or2d1_hd U154 ( .A(n472), .B(n270), .Y(n470) );
  scg13d1_hd U155 ( .A(n472), .B(n270), .C(n138), .Y(n471) );
  nr2d1_hd U158 ( .A(n120), .B(n144), .Y(n472) );
  ad2d1_hd U159 ( .A(w_rstn), .B(sda_negedge), .Y(n473) );
  nd2bd1_hd U162 ( .AN(n43), .B(n442), .Y(n474) );
  oa21d1_hd U163 ( .A(sda_posedge), .B(sda_negedge), .C(n269), .Y(n442) );
  oa211d1_hd U166 ( .A(alt5_n278), .B(n447), .C(n448), .D(alt5_n278), .Y(n446)
         );
  oa211d1_hd U167 ( .A(n22), .B(n449), .C(n450), .D(alt5_n278), .Y(n448) );
  oa21d1_hd U168 ( .A(n451), .B(n120), .C(n22), .Y(n450) );
  oa211d1_hd U169 ( .A(N524), .B(n452), .C(n453), .D(N928), .Y(n449) );
  oa21d1_hd U170 ( .A(n454), .B(n455), .C(N524), .Y(n453) );
  nr3d1_hd U171 ( .A(n23), .B(n82), .C(n44), .Y(n454) );
  ao211d1_hd U173 ( .A(n82), .B(N525), .C(n23), .D(n456), .Y(n452) );
  oa211d1_hd U175 ( .A(N525), .B(n44), .C(n457), .D(N526), .Y(n456) );
  oa211d1_hd U176 ( .A(n451), .B(n44), .C(n459), .D(n457), .Y(n458) );
  scg22d1_hd U179 ( .A(N525), .B(N526), .C(n460), .D(n461), .Y(n459) );
  nr2d1_hd U184 ( .A(n455), .B(n460), .Y(n451) );
  nd3d1_hd U186 ( .A(N525), .B(N526), .C(n457), .Y(n455) );
  ivd1_hd U187 ( .A(N498), .Y(n457) );
  ao22d1_hd U188 ( .A(alt5_n278), .B(n462), .C(alt5_n370), .D(n120), .Y(n443)
         );
  scg22d1_hd U189 ( .A(n37), .B(N629), .C(n145), .D(n463), .Y(n477) );
  scg9d1_hd U191 ( .A(N1034), .B(n464), .C(n37), .Y(n478) );
  ao211d1_hd U196 ( .A(N928), .B(n465), .C(n466), .D(n467), .Y(n464) );
  nr2bd1_hd U199 ( .AN(n82), .B(n151), .Y(n467) );
  ao21d1_hd U200 ( .A(n468), .B(N631), .C(N928), .Y(n466) );
  nr2d1_hd U204 ( .A(n23), .B(n44), .Y(n468) );
  nd3d1_hd U205 ( .A(phy_start_bit), .B(N524), .C(N526), .Y(n465) );
  or2d1_hd U207 ( .A(n18), .B(n43), .Y(n480) );
  ad2d1_hd U217 ( .A(n71), .B(n175), .Y(n481) );
  ad2d1_hd U219 ( .A(n71), .B(n155), .Y(n482) );
  ad2d1_hd U223 ( .A(n71), .B(n165), .Y(n483) );
  ad2d1_hd U228 ( .A(n71), .B(n159), .Y(n484) );
  nd2bd1_hd U229 ( .AN(n43), .B(N132), .Y(n486) );
  ad2d1_hd U230 ( .A(n266), .B(n312), .Y(n487) );
  ad2d1_hd U232 ( .A(n225), .B(n312), .Y(n488) );
  ad2d1_hd U233 ( .A(n226), .B(n312), .Y(n489) );
  ad2d1_hd U234 ( .A(n229), .B(n312), .Y(n490) );
  ad2d1_hd U235 ( .A(n230), .B(n312), .Y(n491) );
  ad2d1_hd U236 ( .A(n231), .B(n312), .Y(n492) );
  ad2d1_hd U237 ( .A(n232), .B(n312), .Y(n493) );
  ad2d1_hd U238 ( .A(n233), .B(n312), .Y(n494) );
  ivd1_hd U239 ( .A(n469), .Y(n496) );
  scg16d1_hd U240 ( .A(n184), .B(n182), .C(n432), .Y(n469) );
  oa21d1_hd U242 ( .A(n174), .B(n223), .C(n177), .Y(n497) );
  ad2d1_hd U244 ( .A(cmd_write_multiple), .B(n427), .Y(n498) );
  ad2d1_hd U245 ( .A(cmd_stop), .B(n427), .Y(n499) );
  ad2d1_hd U274 ( .A(cmd_read), .B(n427), .Y(n500) );
  nr2bd1_hd U282 ( .AN(n433), .B(n220), .Y(n502) );
endmodule


module mpr121_controller_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  had1_hd U2 ( .A(A[8]), .B(n2), .CO(n1), .S(SUM[8]) );
  had1_hd U3 ( .A(A[7]), .B(n3), .CO(n2), .S(SUM[7]) );
  had1_hd U4 ( .A(A[6]), .B(n4), .CO(n3), .S(SUM[6]) );
  had1_hd U5 ( .A(A[5]), .B(n5), .CO(n4), .S(SUM[5]) );
  had1_hd U6 ( .A(A[4]), .B(n6), .CO(n5), .S(SUM[4]) );
  had1_hd U7 ( .A(A[3]), .B(n7), .CO(n6), .S(SUM[3]) );
  had1_hd U8 ( .A(A[2]), .B(n8), .CO(n7), .S(SUM[2]) );
  had1_hd U9 ( .A(A[1]), .B(A[0]), .CO(n8), .S(SUM[1]) );
  xo2d1_hd U13 ( .A(n1), .B(A[9]), .Y(SUM[9]) );
  ivd1_hd U14 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mpr121_controller_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mpr121_controller_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mpr121_controller_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mpr121_controller_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mpr121_controller_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module mpr121_controller ( o_MPR121_DATA_OUT, o_MPR121_REG_ADDR, 
        i_MPR121_DATA_IN, i_MPR121_WRITE_ENABLE, i_MPR121_READ_ENABLE, 
        o_MPR121_INIT_SET, o_MPR121_BUSY, o_MPR121_FAIL, i_I2C_SCL_IN, 
        i_I2C_SDA_IN, o_I2C_SCL_OUT, o_I2C_SDA_OUT, o_I2C_SCL_EN, o_I2C_SDA_EN, 
        i_CLK, i_RSTN );
  output [7:0] o_MPR121_DATA_OUT;
  input [7:0] o_MPR121_REG_ADDR;
  input [7:0] i_MPR121_DATA_IN;
  input i_MPR121_WRITE_ENABLE, i_MPR121_READ_ENABLE, i_I2C_SCL_IN,
         i_I2C_SDA_IN, i_CLK, i_RSTN;
  output o_MPR121_INIT_SET, o_MPR121_BUSY, o_MPR121_FAIL, o_I2C_SCL_OUT,
         o_I2C_SDA_OUT, o_I2C_SCL_EN, o_I2C_SDA_EN;
  wire   w_rstn, r_i2c_start, r_i2c_read, r_i2c_write, r_i2c_write_multiple,
         r_i2c_stop, r_i2c_cmd_valid, r_i2c_data_in_valid, w_i2c_data_in_ready,
         r_i2c_data_in_last, w_i2c_data_out_valid, r_i2c_data_out_ready,
         r_lstate_0_, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N307, N308, N309, N310, N311,
         N312, N315, N324, n40, n46, n47, n78, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n92, n93, n96, n97, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n23,
         n26, n185, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n251,
         n253, n254, n255, n256, n257, n258, n259, n260, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n273;
  wire   [7:0] r_i2c_data_in;
  wire   [7:0] w_i2c_data_out;
  wire   [5:0] r_pstate;
  wire   [9:0] r_clk_counter;
  wire   [7:0] r_i2c_reg_addr;
  wire   [7:0] r_i2c_reg_data_in;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  i2c_master i2c_master ( .i_CLK(i_CLK), .i_RSTN(n26), .cmd_start(r_i2c_start), 
        .cmd_read(r_i2c_read), .cmd_write(r_i2c_write), .cmd_write_multiple(
        r_i2c_write_multiple), .cmd_stop(r_i2c_stop), .cmd_valid(
        r_i2c_cmd_valid), .data_in(r_i2c_data_in), .data_in_valid(
        r_i2c_data_in_valid), .data_in_ready(w_i2c_data_in_ready), 
        .data_in_last(r_i2c_data_in_last), .data_out(w_i2c_data_out), 
        .data_out_valid(w_i2c_data_out_valid), .data_out_ready(
        r_i2c_data_out_ready), .scl_i(i_I2C_SCL_IN), .scl_o(o_I2C_SCL_OUT), 
        .scl_t(o_I2C_SCL_EN), .sda_i(i_I2C_SDA_IN), .sda_o(o_I2C_SDA_OUT), 
        .sda_t(o_I2C_SDA_EN), .missed_ack(o_MPR121_FAIL) );
  clknd2d1_hd U141 ( .A(r_pstate[2]), .B(n114), .Y(n129) );
  clknd2d1_hd U142 ( .A(n161), .B(n84), .Y(n128) );
  clknd2d1_hd U143 ( .A(r_pstate[1]), .B(n161), .Y(n119) );
  clknd2d1_hd U144 ( .A(n83), .B(n146), .Y(n158) );
  clknd2d1_hd U145 ( .A(r_pstate[4]), .B(n160), .Y(n134) );
  clknd2d1_hd U146 ( .A(w_i2c_data_in_ready), .B(n136), .Y(n145) );
  clknd2d1_hd U147 ( .A(n160), .B(n148), .Y(n107) );
  clknd2d1_hd U148 ( .A(n116), .B(n147), .Y(n137) );
  clknd2d1_hd U149 ( .A(i_MPR121_WRITE_ENABLE), .B(n111), .Y(n138) );
  clknd2d1_hd U150 ( .A(n139), .B(n85), .Y(n82) );
  clknd2d1_hd U151 ( .A(n120), .B(n141), .Y(n108) );
  clknd2d1_hd U152 ( .A(n112), .B(n102), .Y(n121) );
  clknd2d1_hd U153 ( .A(n112), .B(n145), .Y(n96) );
  clknd2d1_hd U154 ( .A(r_lstate_0_), .B(n86), .Y(n111) );
  clknd2d1_hd U157 ( .A(n123), .B(n145), .Y(n144) );
  clknd2d1_hd U158 ( .A(n105), .B(i_MPR121_READ_ENABLE), .Y(n131) );
  scg2d1_hd U169 ( .A(n103), .B(n109), .C(o_MPR121_INIT_SET), .D(n89), .Y(n46)
         );
  clknd2d1_hd U184 ( .A(n127), .B(n93), .Y(n97) );
  ivd1_hd U193 ( .A(n96), .Y(n92) );
  oa22ad1_hd U195 ( .A(n103), .B(n104), .C(n105), .D(n106), .Y(n47) );
  oa211d1_hd U196 ( .A(r_pstate[0]), .B(n107), .C(n108), .D(o_MPR121_BUSY), 
        .Y(n104) );
  ivd1_hd U197 ( .A(n110), .Y(n89) );
  ivd1_hd U198 ( .A(n111), .Y(n109) );
  scg22d1_hd U206 ( .A(r_i2c_cmd_valid), .B(n122), .C(n121), .D(n123), .Y(n40)
         );
  nr2d1_hd U217 ( .A(n107), .B(n128), .Y(n110) );
  nr2d1_hd U218 ( .A(n129), .B(n128), .Y(n117) );
  ivd1_hd U219 ( .A(n130), .Y(n127) );
  nr2d1_hd U220 ( .A(n105), .B(n81), .Y(n88) );
  oa211d1_hd U221 ( .A(i_MPR121_WRITE_ENABLE), .B(n131), .C(n132), .D(n133), 
        .Y(N312) );
  scg18d1_hd U222 ( .A(n105), .B(i_MPR121_WRITE_ENABLE), .C(N310), .D(n134), 
        .E(n135), .Y(N311) );
  nr2d1_hd U223 ( .A(n136), .B(n78), .Y(n135) );
  oa211d1_hd U224 ( .A(n137), .B(n138), .C(n122), .D(n82), .Y(N310) );
  ivd1_hd U225 ( .A(n137), .Y(n85) );
  nd2bd1_hd U226 ( .AN(n140), .B(n141), .Y(n122) );
  oa211d1_hd U227 ( .A(w_i2c_data_in_ready), .B(n99), .C(n132), .D(n93), .Y(
        N309) );
  ivd1_hd U228 ( .A(n136), .Y(n93) );
  scg22d1_hd U229 ( .A(r_pstate[0]), .B(r_pstate[1]), .C(i_MPR121_READ_ENABLE), 
        .D(n120), .Y(n132) );
  oa211d1_hd U230 ( .A(n87), .B(n106), .C(n142), .D(n143), .Y(N308) );
  ao21d1_hd U231 ( .A(n103), .B(n138), .C(n144), .Y(n143) );
  oa21d1_hd U232 ( .A(n114), .B(n115), .C(n146), .Y(n123) );
  ivd1_hd U233 ( .A(N324), .Y(n86) );
  nr2d1_hd U234 ( .A(n139), .B(n137), .Y(n103) );
  nr4d1_hd U235 ( .A(r_pstate[5]), .B(r_pstate[2]), .C(n148), .D(n149), .Y(
        n147) );
  nr2d1_hd U236 ( .A(n150), .B(r_clk_counter[9]), .Y(n139) );
  ao211d1_hd U237 ( .A(n151), .B(n152), .C(n153), .D(n154), .Y(n150) );
  nd4d1_hd U238 ( .A(r_clk_counter[5]), .B(r_clk_counter[4]), .C(
        r_clk_counter[8]), .D(r_clk_counter[7]), .Y(n154) );
  ivd1_hd U239 ( .A(r_clk_counter[6]), .Y(n153) );
  ivd1_hd U240 ( .A(r_clk_counter[3]), .Y(n152) );
  oa21d1_hd U241 ( .A(r_clk_counter[1]), .B(r_clk_counter[0]), .C(
        r_clk_counter[2]), .Y(n151) );
  ao211d1_hd U242 ( .A(n120), .B(r_pstate[1]), .C(n155), .D(n130), .Y(n142) );
  or2d1_hd U243 ( .A(i_MPR121_WRITE_ENABLE), .B(i_MPR121_READ_ENABLE), .Y(n106) );
  oa211d1_hd U244 ( .A(n156), .B(n108), .C(n100), .D(n157), .Y(N307) );
  ao211d1_hd U245 ( .A(n80), .B(n81), .C(n155), .D(n101), .Y(n157) );
  ivd1_hd U246 ( .A(n102), .Y(n101) );
  nd3bd1_hd U247 ( .AN(n119), .B(w_i2c_data_out_valid), .C(n120), .Y(n102) );
  nr2bd1_hd U248 ( .AN(w_i2c_data_in_ready), .B(n99), .Y(n155) );
  oa21d1_hd U249 ( .A(n118), .B(n115), .C(n141), .Y(n99) );
  ivd1_hd U250 ( .A(n134), .Y(n115) );
  ivd1_hd U251 ( .A(n158), .Y(n81) );
  ao21d1_hd U252 ( .A(w_i2c_data_in_ready), .B(n130), .C(n96), .Y(n100) );
  nr2d1_hd U253 ( .A(n128), .B(n140), .Y(n136) );
  nd3d1_hd U254 ( .A(r_pstate[4]), .B(r_pstate[2]), .C(n159), .Y(n140) );
  nr2d1_hd U255 ( .A(r_pstate[5]), .B(r_pstate[3]), .Y(n159) );
  oa21d1_hd U256 ( .A(n160), .B(n114), .C(n116), .Y(n112) );
  ivd1_hd U257 ( .A(n128), .Y(n116) );
  ao21d1_hd U258 ( .A(n133), .B(n134), .C(n119), .Y(n130) );
  ivd1_hd U259 ( .A(n118), .Y(n133) );
  nr2d1_hd U260 ( .A(n162), .B(r_pstate[2]), .Y(n118) );
  nr2d1_hd U261 ( .A(n161), .B(n84), .Y(n141) );
  ivd1_hd U262 ( .A(r_pstate[1]), .Y(n84) );
  ivd1_hd U263 ( .A(n129), .Y(n120) );
  ivd1_hd U264 ( .A(n162), .Y(n114) );
  nd3d1_hd U265 ( .A(r_pstate[5]), .B(n148), .C(n149), .Y(n162) );
  ivd1_hd U266 ( .A(r_pstate[3]), .Y(n149) );
  ivd1_hd U267 ( .A(i_MPR121_READ_ENABLE), .Y(n156) );
  nr2bd1_hd U268 ( .AN(i_MPR121_DATA_IN[7]), .B(n87), .Y(N294) );
  scg6d1_hd U269 ( .A(n105), .B(i_MPR121_DATA_IN[6]), .C(n78), .Y(N293) );
  scg6d1_hd U270 ( .A(n105), .B(i_MPR121_DATA_IN[5]), .C(n78), .Y(N292) );
  nr2bd1_hd U271 ( .AN(i_MPR121_DATA_IN[4]), .B(n87), .Y(N291) );
  nr2bd1_hd U272 ( .AN(i_MPR121_DATA_IN[3]), .B(n87), .Y(N290) );
  nr2bd1_hd U273 ( .AN(i_MPR121_DATA_IN[2]), .B(n87), .Y(N289) );
  scg6d1_hd U274 ( .A(n105), .B(i_MPR121_DATA_IN[1]), .C(n78), .Y(N288) );
  scg6d1_hd U275 ( .A(n105), .B(i_MPR121_DATA_IN[0]), .C(n78), .Y(N287) );
  scg6d1_hd U276 ( .A(n105), .B(o_MPR121_REG_ADDR[7]), .C(n78), .Y(N286) );
  nr2d1_hd U277 ( .A(n80), .B(n158), .Y(n78) );
  nr2d1_hd U278 ( .A(r_pstate[1]), .B(n161), .Y(n146) );
  ivd1_hd U279 ( .A(n107), .Y(n83) );
  nr2bd1_hd U281 ( .AN(o_MPR121_REG_ADDR[6]), .B(n87), .Y(N285) );
  nr2bd1_hd U282 ( .AN(o_MPR121_REG_ADDR[5]), .B(n87), .Y(N284) );
  nr2bd1_hd U283 ( .AN(o_MPR121_REG_ADDR[4]), .B(n87), .Y(N283) );
  nr2bd1_hd U284 ( .AN(o_MPR121_REG_ADDR[3]), .B(n87), .Y(N282) );
  nr2bd1_hd U285 ( .AN(o_MPR121_REG_ADDR[2]), .B(n87), .Y(N281) );
  nr2bd1_hd U286 ( .AN(o_MPR121_REG_ADDR[1]), .B(n87), .Y(N280) );
  ivd1_hd U287 ( .A(n105), .Y(n87) );
  ad2d1_hd U288 ( .A(o_MPR121_REG_ADDR[0]), .B(n105), .Y(N279) );
  ivd1_hd U290 ( .A(r_pstate[4]), .Y(n148) );
  nr3d1_hd U291 ( .A(r_pstate[2]), .B(r_pstate[5]), .C(r_pstate[3]), .Y(n160)
         );
  ivd1_hd U292 ( .A(r_pstate[0]), .Y(n161) );
  ivd1_hd U23 ( .A(n185), .Y(n23) );
  ivd1_hd U26 ( .A(n185), .Y(n26) );
  ivd1_hd U57 ( .A(w_rstn), .Y(n185) );
  mpr121_controller_DW01_inc_0 add_x_2 ( .A(r_clk_counter), .SUM({N192, N191, 
        N190, N189, N188, N187, N186, N185, N184, N183}) );
  SNPS_CLOCK_GATE_HIGH_mpr121_controller_10 clk_gate_r_i2c_write_reg_0 ( .CLK(
        i_CLK), .EN(n251), .ENCLK(n203), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mpr121_controller_11 clk_gate_o_MPR121_DATA_OUT_reg_7__0 ( 
        .CLK(i_CLK), .EN(n101), .ENCLK(n202), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mpr121_controller_12 clk_gate_r_i2c_data_in_reg_0__0 ( 
        .CLK(i_CLK), .EN(n198), .ENCLK(n201), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mpr121_controller_13 clk_gate_r_clk_counter_reg_8__0 ( 
        .CLK(i_CLK), .EN(n273), .ENCLK(n200), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mpr121_controller_14 clk_gate_r_i2c_reg_addr_reg_0__0 ( 
        .CLK(i_CLK), .EN(N315), .ENCLK(n199), .TE(1'b0) );
  fd2qd1_hd r_lstate_reg_0_ ( .D(n204), .CK(i_CLK), .RN(n26), .Q(r_lstate_0_)
         );
  fd1qd1_hd r_i2c_reg_data_in_reg_5_ ( .D(N292), .CK(n199), .Q(
        r_i2c_reg_data_in[5]) );
  fd1qd1_hd r_i2c_reg_data_in_reg_7_ ( .D(N294), .CK(n199), .Q(
        r_i2c_reg_data_in[7]) );
  fd1qd1_hd r_i2c_reg_data_in_reg_3_ ( .D(N290), .CK(n199), .Q(
        r_i2c_reg_data_in[3]) );
  fd1qd1_hd r_i2c_reg_data_in_reg_2_ ( .D(N289), .CK(n199), .Q(
        r_i2c_reg_data_in[2]) );
  fd1qd1_hd r_i2c_reg_addr_reg_6_ ( .D(N285), .CK(n199), .Q(r_i2c_reg_addr[6])
         );
  fd1qd1_hd r_i2c_reg_addr_reg_4_ ( .D(N283), .CK(n199), .Q(r_i2c_reg_addr[4])
         );
  fd1qd1_hd r_i2c_reg_addr_reg_2_ ( .D(N281), .CK(n199), .Q(r_i2c_reg_addr[2])
         );
  fd1qd1_hd r_i2c_reg_data_in_reg_4_ ( .D(N291), .CK(n199), .Q(
        r_i2c_reg_data_in[4]) );
  fd1qd1_hd r_i2c_reg_addr_reg_5_ ( .D(N284), .CK(n199), .Q(r_i2c_reg_addr[5])
         );
  fd1qd1_hd r_i2c_reg_addr_reg_3_ ( .D(N282), .CK(n199), .Q(r_i2c_reg_addr[3])
         );
  fd1qd1_hd r_i2c_reg_addr_reg_1_ ( .D(N280), .CK(n199), .Q(r_i2c_reg_addr[1])
         );
  fd1qd1_hd r_i2c_reg_addr_reg_0_ ( .D(N279), .CK(n199), .Q(r_i2c_reg_addr[0])
         );
  fd1qd1_hd r_i2c_reg_data_in_reg_6_ ( .D(N293), .CK(n199), .Q(
        r_i2c_reg_data_in[6]) );
  fd1qd1_hd r_i2c_reg_data_in_reg_1_ ( .D(N288), .CK(n199), .Q(
        r_i2c_reg_data_in[1]) );
  fd1qd1_hd r_i2c_reg_data_in_reg_0_ ( .D(N287), .CK(n199), .Q(
        r_i2c_reg_data_in[0]) );
  fd1qd1_hd r_i2c_reg_addr_reg_7_ ( .D(N286), .CK(n199), .Q(r_i2c_reg_addr[7])
         );
  fd2qd1_hd r_i2c_write_multiple_reg ( .D(n115), .CK(n203), .RN(w_rstn), .Q(
        r_i2c_write_multiple) );
  fd2qd1_hd r_i2c_write_reg ( .D(n118), .CK(n203), .RN(n23), .Q(r_i2c_write)
         );
  fd2qd1_hd r_i2c_read_reg ( .D(r_pstate[2]), .CK(n203), .RN(n23), .Q(
        r_i2c_read) );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_6_ ( .D(w_i2c_data_out[6]), .CK(n202), .RN(
        n23), .Q(o_MPR121_DATA_OUT[6]) );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_4_ ( .D(w_i2c_data_out[4]), .CK(n202), .RN(
        n23), .Q(o_MPR121_DATA_OUT[4]) );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_2_ ( .D(w_i2c_data_out[2]), .CK(n202), .RN(
        n23), .Q(o_MPR121_DATA_OUT[2]) );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_0_ ( .D(w_i2c_data_out[0]), .CK(n202), .RN(
        n23), .Q(o_MPR121_DATA_OUT[0]) );
  fd2qd1_hd r_i2c_start_reg ( .D(n249), .CK(n203), .RN(n26), .Q(r_i2c_start)
         );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_7_ ( .D(w_i2c_data_out[7]), .CK(n202), .RN(
        n26), .Q(o_MPR121_DATA_OUT[7]) );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_5_ ( .D(w_i2c_data_out[5]), .CK(n202), .RN(
        n26), .Q(o_MPR121_DATA_OUT[5]) );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_3_ ( .D(w_i2c_data_out[3]), .CK(n202), .RN(
        n26), .Q(o_MPR121_DATA_OUT[3]) );
  fd2qd1_hd o_MPR121_DATA_OUT_reg_1_ ( .D(w_i2c_data_out[1]), .CK(n202), .RN(
        n26), .Q(o_MPR121_DATA_OUT[1]) );
  fd2qd1_hd r_i2c_data_in_last_reg ( .D(n210), .CK(i_CLK), .RN(n26), .Q(
        r_i2c_data_in_last) );
  fd2qd1_hd r_i2c_data_in_reg_0_ ( .D(n260), .CK(n201), .RN(n23), .Q(
        r_i2c_data_in[0]) );
  fd2qd1_hd r_i2c_cmd_valid_reg ( .D(n40), .CK(i_CLK), .RN(n26), .Q(
        r_i2c_cmd_valid) );
  fd2qd1_hd r_i2c_stop_reg ( .D(n206), .CK(i_CLK), .RN(w_rstn), .Q(r_i2c_stop)
         );
  fd2qd1_hd r_i2c_data_out_ready_reg ( .D(n207), .CK(i_CLK), .RN(n23), .Q(
        r_i2c_data_out_ready) );
  fd2qd1_hd r_i2c_data_in_valid_reg ( .D(n209), .CK(i_CLK), .RN(n23), .Q(
        r_i2c_data_in_valid) );
  fd2qd1_hd o_MPR121_INIT_SET_reg ( .D(n46), .CK(n200), .RN(n23), .Q(
        o_MPR121_INIT_SET) );
  fd2qd1_hd r_clk_counter_reg_7_ ( .D(n270), .CK(n200), .RN(n26), .Q(
        r_clk_counter[7]) );
  fd2qd1_hd r_clk_counter_reg_6_ ( .D(n269), .CK(n200), .RN(n23), .Q(
        r_clk_counter[6]) );
  fd2qd1_hd r_i2c_data_in_reg_7_ ( .D(n259), .CK(n201), .RN(w_rstn), .Q(
        r_i2c_data_in[7]) );
  fd2qd1_hd r_i2c_data_in_reg_6_ ( .D(n258), .CK(n201), .RN(w_rstn), .Q(
        r_i2c_data_in[6]) );
  fd2qd1_hd r_i2c_data_in_reg_5_ ( .D(n257), .CK(n201), .RN(n26), .Q(
        r_i2c_data_in[5]) );
  fd2qd1_hd r_i2c_data_in_reg_4_ ( .D(n256), .CK(n201), .RN(n26), .Q(
        r_i2c_data_in[4]) );
  fd2qd1_hd r_i2c_data_in_reg_3_ ( .D(n255), .CK(n201), .RN(w_rstn), .Q(
        r_i2c_data_in[3]) );
  fd2qd1_hd r_i2c_data_in_reg_2_ ( .D(n254), .CK(n201), .RN(w_rstn), .Q(
        r_i2c_data_in[2]) );
  fd2qd1_hd r_i2c_data_in_reg_1_ ( .D(n253), .CK(n201), .RN(w_rstn), .Q(
        r_i2c_data_in[1]) );
  fd2qd1_hd r_clk_counter_reg_5_ ( .D(n268), .CK(n200), .RN(n26), .Q(
        r_clk_counter[5]) );
  fd2qd1_hd r_clk_counter_reg_4_ ( .D(n267), .CK(n200), .RN(n23), .Q(
        r_clk_counter[4]) );
  fd2qd1_hd r_clk_counter_reg_3_ ( .D(n266), .CK(n200), .RN(n26), .Q(
        r_clk_counter[3]) );
  fd2qd1_hd r_clk_counter_reg_2_ ( .D(n265), .CK(n200), .RN(n23), .Q(
        r_clk_counter[2]) );
  fd2qd1_hd r_clk_counter_reg_1_ ( .D(n264), .CK(n200), .RN(n26), .Q(
        r_clk_counter[1]) );
  fd2qd1_hd r_clk_counter_reg_0_ ( .D(n263), .CK(n200), .RN(n23), .Q(
        r_clk_counter[0]) );
  fd2qd1_hd r_clk_counter_reg_9_ ( .D(n262), .CK(n200), .RN(n23), .Q(
        r_clk_counter[9]) );
  fd2qd1_hd r_clk_counter_reg_8_ ( .D(n271), .CK(n200), .RN(n23), .Q(
        r_clk_counter[8]) );
  fd2qd1_hd r_lstate_reg_1_ ( .D(n205), .CK(i_CLK), .RN(n26), .Q(N324) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(N307), .CK(i_CLK), .RN(w_rstn), .Q(
        r_pstate[0]) );
  fd2qd1_hd r_pstate_reg_2_ ( .D(N309), .CK(i_CLK), .RN(w_rstn), .Q(
        r_pstate[2]) );
  fd2qd1_hd r_pstate_reg_5_ ( .D(N312), .CK(i_CLK), .RN(w_rstn), .Q(
        r_pstate[5]) );
  fd2qd1_hd o_MPR121_BUSY_reg ( .D(n47), .CK(i_CLK), .RN(w_rstn), .Q(
        o_MPR121_BUSY) );
  fd2qd1_hd r_pstate_reg_1_ ( .D(N308), .CK(i_CLK), .RN(w_rstn), .Q(
        r_pstate[1]) );
  fd2qd1_hd r_pstate_reg_4_ ( .D(N311), .CK(i_CLK), .RN(w_rstn), .Q(
        r_pstate[4]) );
  fd2qd1_hd r_pstate_reg_3_ ( .D(n208), .CK(i_CLK), .RN(w_rstn), .Q(
        r_pstate[3]) );
  nr2bd1_hd U1 ( .AN(w_rstn), .B(n88), .Y(N315) );
  mx2d1_hd U2 ( .D0(r_pstate[3]), .D1(n245), .S(n246), .Y(n208) );
  scg2d1_hd U3 ( .A(n136), .B(r_i2c_reg_data_in[1]), .C(r_i2c_reg_addr[1]), 
        .D(n215), .Y(n253) );
  scg2d1_hd U4 ( .A(n136), .B(r_i2c_reg_data_in[2]), .C(r_i2c_reg_addr[2]), 
        .D(n215), .Y(n254) );
  scg2d1_hd U5 ( .A(n136), .B(r_i2c_reg_data_in[3]), .C(r_i2c_reg_addr[3]), 
        .D(n215), .Y(n255) );
  scg2d1_hd U6 ( .A(n136), .B(r_i2c_reg_data_in[4]), .C(r_i2c_reg_addr[4]), 
        .D(n215), .Y(n256) );
  scg2d1_hd U7 ( .A(n136), .B(r_i2c_reg_data_in[5]), .C(r_i2c_reg_addr[5]), 
        .D(n215), .Y(n257) );
  scg2d1_hd U8 ( .A(n136), .B(r_i2c_reg_data_in[6]), .C(r_i2c_reg_addr[6]), 
        .D(n215), .Y(n258) );
  scg2d1_hd U9 ( .A(r_i2c_reg_addr[7]), .B(n215), .C(r_i2c_reg_data_in[7]), 
        .D(n136), .Y(n259) );
  clknd2d1_hd U10 ( .A(r_pstate[1]), .B(n137), .Y(n233) );
  clknd2d1_hd U11 ( .A(r_pstate[1]), .B(n137), .Y(n236) );
  mx2d1_hd U12 ( .D0(r_i2c_data_in_valid), .D1(n97), .S(n244), .Y(n209) );
  mx2d1_hd U13 ( .D0(r_i2c_data_out_ready), .D1(n247), .S(n121), .Y(n207) );
  mx2d1_hd U14 ( .D0(r_i2c_stop), .D1(n247), .S(n121), .Y(n206) );
  mx2d1_hd U15 ( .D0(r_i2c_data_in_last), .D1(n242), .S(n243), .Y(n210) );
  mx2d1_hd U16 ( .D0(n136), .D1(n116), .S(n118), .Y(n242) );
  mx2d1_hd U17 ( .D0(r_lstate_0_), .D1(n78), .S(n248), .Y(n204) );
  mx2d1_hd U18 ( .D0(N324), .D1(n105), .S(n248), .Y(n205) );
  nr2ad1_hd U19 ( .A(n119), .B(n107), .Y(n105) );
  nr4d2_hd U20 ( .A(r_clk_counter[6]), .B(r_clk_counter[8]), .C(
        r_clk_counter[7]), .D(r_clk_counter[9]), .Y(n80) );
  ad2d1_hd U21 ( .A(n88), .B(n89), .Y(n197) );
  scg8d1_hd U22 ( .A(w_i2c_data_in_ready), .B(n97), .C(n117), .D(n110), .Y(
        n198) );
  scg14d1_hd U24 ( .A(n116), .B(n118), .C(n92), .Y(n243) );
  oa21d1_hd U25 ( .A(w_i2c_data_in_ready), .B(n99), .C(n211), .Y(n244) );
  ao21d1_hd U27 ( .A(n130), .B(w_i2c_data_in_ready), .C(n96), .Y(n211) );
  nr2d1_hd U28 ( .A(r_pstate[5]), .B(n212), .Y(n245) );
  nd4d1_hd U29 ( .A(r_pstate[2]), .B(n141), .C(r_pstate[4]), .D(n149), .Y(n212) );
  oa211d1_hd U30 ( .A(n139), .B(n213), .C(n116), .D(n214), .Y(n246) );
  nr3d1_hd U31 ( .A(r_pstate[2]), .B(r_pstate[5]), .C(n148), .Y(n214) );
  ivd1_hd U32 ( .A(n138), .Y(n213) );
  nr2bd1_hd U33 ( .AN(n120), .B(n119), .Y(n247) );
  nd2bd1_hd U34 ( .AN(n78), .B(n197), .Y(n248) );
  or2d1_hd U35 ( .A(n114), .B(n115), .Y(n249) );
  scg9d1_hd U36 ( .A(n160), .B(n114), .C(n116), .Y(n251) );
  ivd1_hd U37 ( .A(n127), .Y(n215) );
  oa22d1_hd U38 ( .A(n127), .B(n216), .C(n93), .D(n217), .Y(n260) );
  ivd1_hd U39 ( .A(r_i2c_reg_data_in[0]), .Y(n217) );
  ivd1_hd U40 ( .A(r_i2c_reg_addr[0]), .Y(n216) );
  ao21d1_hd U41 ( .A(n218), .B(n219), .C(n220), .Y(n262) );
  ivd1_hd U42 ( .A(N192), .Y(n220) );
  scg17d1_hd U43 ( .A(r_clk_counter[5]), .B(n221), .C(r_clk_counter[9]), .D(
        n85), .Y(n219) );
  ao21d1_hd U44 ( .A(n151), .B(n152), .C(n222), .Y(n221) );
  nd4d1_hd U45 ( .A(r_clk_counter[8]), .B(r_clk_counter[6]), .C(
        r_clk_counter[7]), .D(r_clk_counter[4]), .Y(n222) );
  scg18d1_hd U46 ( .A(n223), .B(r_clk_counter[9]), .C(r_clk_counter[8]), .D(
        n224), .E(n146), .Y(n218) );
  nr2d1_hd U47 ( .A(r_clk_counter[6]), .B(r_clk_counter[7]), .Y(n224) );
  nd2bd1_hd U48 ( .AN(n85), .B(r_pstate[1]), .Y(n223) );
  nr2bd1_hd U49 ( .AN(N183), .B(n225), .Y(n263) );
  ao22d1_hd U50 ( .A(n139), .B(n85), .C(n80), .D(n81), .Y(n225) );
  nr2bd1_hd U51 ( .AN(N184), .B(n226), .Y(n264) );
  ao22d1_hd U52 ( .A(n139), .B(n85), .C(n80), .D(n81), .Y(n226) );
  nr2bd1_hd U53 ( .AN(N185), .B(n227), .Y(n265) );
  ao22d1_hd U54 ( .A(n139), .B(n85), .C(n80), .D(n81), .Y(n227) );
  nr2bd1_hd U55 ( .AN(N186), .B(n228), .Y(n266) );
  ao22d1_hd U56 ( .A(n139), .B(n85), .C(n80), .D(n81), .Y(n228) );
  nr2bd1_hd U58 ( .AN(N187), .B(n229), .Y(n267) );
  ao22d1_hd U59 ( .A(n139), .B(n85), .C(n80), .D(n81), .Y(n229) );
  nr2bd1_hd U60 ( .AN(N188), .B(n230), .Y(n268) );
  ao22d1_hd U61 ( .A(n139), .B(n85), .C(n80), .D(n81), .Y(n230) );
  scg12d1_hd U62 ( .A(n231), .B(N189), .C(r_clk_counter[9]), .Y(n269) );
  oa22d1_hd U63 ( .A(r_clk_counter[7]), .B(n232), .C(n150), .D(n137), .Y(n231)
         );
  scg18d1_hd U64 ( .A(n233), .B(r_clk_counter[6]), .C(r_clk_counter[8]), .D(
        n146), .E(n83), .Y(n232) );
  scg12d1_hd U65 ( .A(n234), .B(N190), .C(r_clk_counter[9]), .Y(n270) );
  oa22d1_hd U66 ( .A(r_clk_counter[8]), .B(n235), .C(n150), .D(n137), .Y(n234)
         );
  scg18d1_hd U67 ( .A(n236), .B(r_clk_counter[7]), .C(r_clk_counter[6]), .D(
        n146), .E(n83), .Y(n235) );
  scg12d1_hd U68 ( .A(N191), .B(n237), .C(r_clk_counter[9]), .Y(n271) );
  scg16d1_hd U69 ( .A(n85), .B(n150), .C(n238), .Y(n237) );
  nd4d1_hd U70 ( .A(n83), .B(n146), .C(n239), .D(n240), .Y(n238) );
  oa21d1_hd U71 ( .A(n85), .B(n84), .C(r_clk_counter[8]), .Y(n240) );
  nr2d1_hd U72 ( .A(r_clk_counter[7]), .B(r_clk_counter[6]), .Y(n239) );
  scg17d1_hd U73 ( .A(n83), .B(n84), .C(n85), .D(n241), .Y(n273) );
  nd3d1_hd U74 ( .A(n81), .B(N188), .C(n80), .Y(n241) );
endmodule


module converter_i2f_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  had1_hd U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  had1_hd U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  had1_hd U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  had1_hd U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  had1_hd U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  had1_hd U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  xo2d1_hd U11 ( .A(n1), .B(A[7]), .Y(SUM[7]) );
  ivd1_hd U12 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module converter_i2f_DW01_inc_1 ( A, SUM );
  input [23:0] A;
  output [23:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;

  had1_hd U2 ( .A(A[22]), .B(n2), .CO(n1), .S(SUM[22]) );
  had1_hd U3 ( .A(A[21]), .B(n3), .CO(n2), .S(SUM[21]) );
  had1_hd U4 ( .A(A[20]), .B(n4), .CO(n3), .S(SUM[20]) );
  had1_hd U5 ( .A(A[19]), .B(n5), .CO(n4), .S(SUM[19]) );
  had1_hd U6 ( .A(A[18]), .B(n6), .CO(n5), .S(SUM[18]) );
  had1_hd U7 ( .A(A[17]), .B(n7), .CO(n6), .S(SUM[17]) );
  had1_hd U8 ( .A(A[16]), .B(n8), .CO(n7), .S(SUM[16]) );
  had1_hd U9 ( .A(A[15]), .B(n9), .CO(n8), .S(SUM[15]) );
  had1_hd U10 ( .A(A[14]), .B(n10), .CO(n9), .S(SUM[14]) );
  had1_hd U11 ( .A(A[13]), .B(n11), .CO(n10), .S(SUM[13]) );
  had1_hd U12 ( .A(A[12]), .B(n12), .CO(n11), .S(SUM[12]) );
  had1_hd U13 ( .A(A[11]), .B(n13), .CO(n12), .S(SUM[11]) );
  had1_hd U14 ( .A(A[10]), .B(n14), .CO(n13), .S(SUM[10]) );
  had1_hd U15 ( .A(A[9]), .B(n15), .CO(n14), .S(SUM[9]) );
  had1_hd U16 ( .A(A[8]), .B(n16), .CO(n15), .S(SUM[8]) );
  had1_hd U17 ( .A(A[7]), .B(n17), .CO(n16), .S(SUM[7]) );
  had1_hd U18 ( .A(A[6]), .B(n18), .CO(n17), .S(SUM[6]) );
  had1_hd U19 ( .A(A[5]), .B(n19), .CO(n18), .S(SUM[5]) );
  had1_hd U20 ( .A(A[4]), .B(n20), .CO(n19), .S(SUM[4]) );
  had1_hd U21 ( .A(A[3]), .B(n21), .CO(n20), .S(SUM[3]) );
  had1_hd U22 ( .A(A[2]), .B(n22), .CO(n21), .S(SUM[2]) );
  had1_hd U23 ( .A(A[1]), .B(A[0]), .CO(n22), .S(SUM[1]) );
  xo2d1_hd U27 ( .A(n1), .B(A[23]), .Y(SUM[23]) );
  ivd1_hd U28 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module converter_i2f_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62;

  had1_hd U2 ( .A(n33), .B(n2), .CO(n1), .S(DIFF[30]) );
  had1_hd U3 ( .A(n34), .B(n3), .CO(n2), .S(DIFF[29]) );
  had1_hd U4 ( .A(n35), .B(n4), .CO(n3), .S(DIFF[28]) );
  had1_hd U5 ( .A(n36), .B(n5), .CO(n4), .S(DIFF[27]) );
  had1_hd U6 ( .A(n37), .B(n6), .CO(n5), .S(DIFF[26]) );
  had1_hd U7 ( .A(n38), .B(n7), .CO(n6), .S(DIFF[25]) );
  had1_hd U8 ( .A(n39), .B(n8), .CO(n7), .S(DIFF[24]) );
  had1_hd U9 ( .A(n40), .B(n9), .CO(n8), .S(DIFF[23]) );
  had1_hd U10 ( .A(n41), .B(n10), .CO(n9), .S(DIFF[22]) );
  had1_hd U11 ( .A(n42), .B(n11), .CO(n10), .S(DIFF[21]) );
  had1_hd U12 ( .A(n43), .B(n12), .CO(n11), .S(DIFF[20]) );
  had1_hd U13 ( .A(n44), .B(n13), .CO(n12), .S(DIFF[19]) );
  had1_hd U14 ( .A(n45), .B(n14), .CO(n13), .S(DIFF[18]) );
  had1_hd U15 ( .A(n46), .B(n15), .CO(n14), .S(DIFF[17]) );
  had1_hd U16 ( .A(n47), .B(n16), .CO(n15), .S(DIFF[16]) );
  had1_hd U17 ( .A(n48), .B(n17), .CO(n16), .S(DIFF[15]) );
  had1_hd U18 ( .A(n49), .B(n18), .CO(n17), .S(DIFF[14]) );
  had1_hd U19 ( .A(n50), .B(n19), .CO(n18), .S(DIFF[13]) );
  had1_hd U20 ( .A(n51), .B(n20), .CO(n19), .S(DIFF[12]) );
  had1_hd U21 ( .A(n52), .B(n21), .CO(n20), .S(DIFF[11]) );
  had1_hd U22 ( .A(n53), .B(n22), .CO(n21), .S(DIFF[10]) );
  had1_hd U23 ( .A(n54), .B(n23), .CO(n22), .S(DIFF[9]) );
  had1_hd U24 ( .A(n55), .B(n24), .CO(n23), .S(DIFF[8]) );
  had1_hd U25 ( .A(n56), .B(n25), .CO(n24), .S(DIFF[7]) );
  had1_hd U26 ( .A(n57), .B(n26), .CO(n25), .S(DIFF[6]) );
  had1_hd U27 ( .A(n58), .B(n27), .CO(n26), .S(DIFF[5]) );
  had1_hd U28 ( .A(n59), .B(n28), .CO(n27), .S(DIFF[4]) );
  had1_hd U29 ( .A(n60), .B(n29), .CO(n28), .S(DIFF[3]) );
  had1_hd U30 ( .A(n61), .B(n30), .CO(n29), .S(DIFF[2]) );
  had1_hd U31 ( .A(n62), .B(n31), .CO(n30), .S(DIFF[1]) );
  nid1_hd U68 ( .A(B[0]), .Y(DIFF[0]) );
  ivd1_hd U69 ( .A(B[1]), .Y(n62) );
  ivd1_hd U70 ( .A(B[2]), .Y(n61) );
  ivd1_hd U71 ( .A(B[3]), .Y(n60) );
  ivd1_hd U72 ( .A(B[4]), .Y(n59) );
  ivd1_hd U73 ( .A(B[5]), .Y(n58) );
  ivd1_hd U74 ( .A(B[6]), .Y(n57) );
  ivd1_hd U75 ( .A(B[7]), .Y(n56) );
  ivd1_hd U76 ( .A(B[8]), .Y(n55) );
  ivd1_hd U77 ( .A(B[9]), .Y(n54) );
  ivd1_hd U78 ( .A(B[10]), .Y(n53) );
  ivd1_hd U79 ( .A(B[11]), .Y(n52) );
  ivd1_hd U80 ( .A(B[12]), .Y(n51) );
  ivd1_hd U81 ( .A(B[13]), .Y(n50) );
  ivd1_hd U82 ( .A(B[14]), .Y(n49) );
  ivd1_hd U83 ( .A(B[15]), .Y(n48) );
  ivd1_hd U84 ( .A(B[16]), .Y(n47) );
  ivd1_hd U85 ( .A(B[17]), .Y(n46) );
  ivd1_hd U86 ( .A(B[18]), .Y(n45) );
  ivd1_hd U87 ( .A(B[19]), .Y(n44) );
  ivd1_hd U88 ( .A(B[20]), .Y(n43) );
  ivd1_hd U89 ( .A(B[21]), .Y(n42) );
  ivd1_hd U90 ( .A(B[22]), .Y(n41) );
  ivd1_hd U91 ( .A(B[23]), .Y(n40) );
  ivd1_hd U92 ( .A(B[24]), .Y(n39) );
  ivd1_hd U93 ( .A(B[25]), .Y(n38) );
  ivd1_hd U94 ( .A(B[26]), .Y(n37) );
  ivd1_hd U95 ( .A(B[27]), .Y(n36) );
  ivd1_hd U96 ( .A(B[28]), .Y(n35) );
  ivd1_hd U97 ( .A(B[29]), .Y(n34) );
  ivd1_hd U98 ( .A(B[30]), .Y(n33) );
  ivd1_hd U99 ( .A(B[0]), .Y(n31) );
  xn2d1_hd U100 ( .A(n1), .B(B[31]), .Y(DIFF[31]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_i2f_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_i2f_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_i2f_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_i2f_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_i2f_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_i2f_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module converter_i2f ( i_A, i_A_STB, o_A_ACK, o_Z, o_Z_STB, i_Z_ACK, i_CLK, 
        i_RST );
  input [31:0] i_A;
  output [31:0] o_Z;
  input i_A_STB, i_Z_ACK, i_CLK, i_RST;
  output o_A_ACK, o_Z_STB;
  wire   n243, n244, n245, n246, n247, n248, n249, n250, n242, n251, N6, N23,
         N24, N25, N26, N27, N28, N31, N34, N37, N40, N43, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N118, N119, N120, N121, N122, N123, N124, N125, sticky, N127, N130,
         N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N180, N184,
         N185, N210, N211, N220, N229, N230, N231, N232, N233, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N293, N305, N308, N309, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n194, n195, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, state_1_, n12, n21, n22, n23, n24, n26,
         n27, n29, n30, n32, n33, n35, n36, n38, n39, n41, n42, n44, n45, n47,
         n48, n50, n51, n53, n54, n56, n57, n59, n60, n62, n63, n65, n66, n68,
         n69, n71, n72, n74, n75, n77, n78, n80, n81, n83, n84, n86, n87, n89,
         n90, n92, n93, n94, n96, n98, n100, n102, n104, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n196, n197, n232, n233, n234, n236, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285;
  wire   [31:0] value;
  wire   [7:0] z_e;
  wire   [23:0] z_m;
  wire   [7:0] z_r;

  ivd1_hd U3 ( .A(i_RST), .Y(n1) );
  ivd1_hd U4 ( .A(i_RST), .Y(n2) );
  ivd1_hd U5 ( .A(i_RST), .Y(n3) );
  ivd1_hd U6 ( .A(i_RST), .Y(n4) );
  ivd1_hd U7 ( .A(i_RST), .Y(n5) );
  ad2d1_hd U32 ( .A(n143), .B(n198), .Y(z_r[0]) );
  ao22d1_hd U34 ( .A(N6), .B(N125), .C(n199), .D(N161), .Y(n7) );
  ao22d1_hd U36 ( .A(N6), .B(N124), .C(n199), .D(N160), .Y(n9) );
  ao22d1_hd U38 ( .A(N6), .B(N123), .C(n199), .D(N159), .Y(n10) );
  ao22d1_hd U40 ( .A(N6), .B(N122), .C(n199), .D(N158), .Y(n11) );
  ao22d1_hd U42 ( .A(N6), .B(N121), .C(n199), .D(N157), .Y(n13) );
  ao22d1_hd U44 ( .A(N6), .B(N120), .C(n199), .D(N156), .Y(n14) );
  ao22d1_hd U46 ( .A(N6), .B(N119), .C(n199), .D(N155), .Y(n15) );
  ao22d1_hd U49 ( .A(N6), .B(N118), .C(n199), .D(N154), .Y(n16) );
  scg17d1_hd U50 ( .A(N257), .B(n17), .C(N220), .D(n18), .Y(N211) );
  ad2d1_hd U52 ( .A(n199), .B(N127), .Y(n17) );
  scg6d1_hd U53 ( .A(n19), .B(N6), .C(n198), .Y(N220) );
  scg5d1_hd U54 ( .A(n198), .B(n159), .C(n199), .D(N153), .E(N6), .F(n93), .Y(
        z_m[23]) );
  scg5d1_hd U55 ( .A(n198), .B(n145), .C(n199), .D(N152), .E(N6), .F(n90), .Y(
        z_m[22]) );
  scg5d1_hd U56 ( .A(n198), .B(n144), .C(n199), .D(N151), .E(N6), .F(n87), .Y(
        z_m[21]) );
  scg5d1_hd U57 ( .A(n198), .B(n115), .C(n199), .D(N150), .E(N6), .F(n84), .Y(
        z_m[20]) );
  scg5d1_hd U58 ( .A(n198), .B(n116), .C(n199), .D(N149), .E(N6), .F(n81), .Y(
        z_m[19]) );
  scg5d1_hd U59 ( .A(n198), .B(n117), .C(n199), .D(N148), .E(N6), .F(n78), .Y(
        z_m[18]) );
  scg5d1_hd U60 ( .A(n198), .B(n118), .C(n199), .D(N147), .E(N6), .F(n75), .Y(
        z_m[17]) );
  scg5d1_hd U61 ( .A(n198), .B(n119), .C(n199), .D(N146), .E(N6), .F(n72), .Y(
        z_m[16]) );
  scg5d1_hd U62 ( .A(n198), .B(n120), .C(n199), .D(N145), .E(N6), .F(n69), .Y(
        z_m[15]) );
  scg5d1_hd U63 ( .A(n198), .B(n121), .C(n199), .D(N144), .E(N6), .F(n66), .Y(
        z_m[14]) );
  scg5d1_hd U64 ( .A(n198), .B(n122), .C(n199), .D(N143), .E(N6), .F(n63), .Y(
        z_m[13]) );
  scg5d1_hd U65 ( .A(n198), .B(n123), .C(n199), .D(N142), .E(N6), .F(n60), .Y(
        z_m[12]) );
  scg5d1_hd U66 ( .A(n198), .B(n124), .C(n199), .D(N141), .E(N6), .F(n57), .Y(
        z_m[11]) );
  scg5d1_hd U67 ( .A(n198), .B(n125), .C(n199), .D(N140), .E(N6), .F(n54), .Y(
        z_m[10]) );
  scg5d1_hd U68 ( .A(n198), .B(n126), .C(n199), .D(N139), .E(N6), .F(n51), .Y(
        z_m[9]) );
  scg5d1_hd U69 ( .A(n198), .B(n127), .C(n199), .D(N138), .E(N6), .F(n48), .Y(
        z_m[8]) );
  scg5d1_hd U70 ( .A(n198), .B(n128), .C(n199), .D(N137), .E(N6), .F(n45), .Y(
        z_m[7]) );
  scg5d1_hd U71 ( .A(n198), .B(n129), .C(n199), .D(N136), .E(N6), .F(n42), .Y(
        z_m[6]) );
  scg5d1_hd U72 ( .A(n198), .B(n130), .C(n199), .D(N135), .E(N6), .F(n39), .Y(
        z_m[5]) );
  scg5d1_hd U73 ( .A(n198), .B(n131), .C(n199), .D(N134), .E(N6), .F(n36), .Y(
        z_m[4]) );
  scg5d1_hd U74 ( .A(n198), .B(n132), .C(n199), .D(N133), .E(N6), .F(n33), .Y(
        z_m[3]) );
  scg5d1_hd U75 ( .A(n198), .B(n133), .C(n199), .D(N132), .E(N6), .F(n30), .Y(
        z_m[2]) );
  scg5d1_hd U76 ( .A(n198), .B(n134), .C(n199), .D(N131), .E(N6), .F(n27), .Y(
        z_m[1]) );
  scg5d1_hd U77 ( .A(n198), .B(n135), .C(n199), .D(N130), .E(N6), .F(n108), 
        .Y(z_m[0]) );
  or2d1_hd U79 ( .A(N185), .B(N305), .Y(state_1_) );
  ivd1_hd U81 ( .A(n195), .Y(n8) );
  scg16d1_hd U84 ( .A(n202), .B(n251), .C(n20), .Y(N180) );
  nr3d1_hd U85 ( .A(N229), .B(N184), .C(N293), .Y(n20) );
  nr2bd1_hd U87 ( .AN(N6), .B(n19), .Y(N229) );
  ivd1_hd U88 ( .A(n94), .Y(n19) );
  nr2d1_hd U89 ( .A(n194), .B(n6), .Y(n243) );
  nr2bd1_hd U90 ( .AN(N82), .B(n6), .Y(value[31]) );
  or2d1_hd U107 ( .A(n168), .B(N286), .Y(N287) );
  or2d1_hd U108 ( .A(n169), .B(N285), .Y(N286) );
  or2d1_hd U109 ( .A(n170), .B(N284), .Y(N285) );
  clknd2d1_hd U110 ( .A(n195), .B(n194), .Y(n18) );
  ad2d1_hd U111 ( .A(n27), .B(N256), .Y(N257) );
  ad2d1_hd U112 ( .A(n30), .B(N255), .Y(N256) );
  ad2d1_hd U113 ( .A(n33), .B(N254), .Y(N255) );
  or2d1_hd U114 ( .A(n197), .B(N259), .Y(N260) );
  or2d1_hd U115 ( .A(n232), .B(N258), .Y(N259) );
  or2d1_hd U116 ( .A(n233), .B(n234), .Y(N258) );
  or2d1_hd U117 ( .A(n191), .B(N263), .Y(N264) );
  or2d1_hd U118 ( .A(n192), .B(N262), .Y(N263) );
  or2d1_hd U119 ( .A(n193), .B(N261), .Y(N262) );
  or2d1_hd U120 ( .A(n196), .B(N260), .Y(N261) );
  or2d1_hd U121 ( .A(n187), .B(N267), .Y(N268) );
  or2d1_hd U122 ( .A(n188), .B(N266), .Y(N267) );
  or2d1_hd U123 ( .A(n189), .B(N265), .Y(N266) );
  or2d1_hd U124 ( .A(n190), .B(N264), .Y(N265) );
  ad2d1_hd U125 ( .A(n84), .B(N237), .Y(N238) );
  ad2d1_hd U126 ( .A(n87), .B(N236), .Y(N237) );
  ad2d1_hd U127 ( .A(n90), .B(N235), .Y(N236) );
  ad2d1_hd U128 ( .A(n93), .B(n94), .Y(N235) );
  or2d1_hd U129 ( .A(n183), .B(N271), .Y(N272) );
  or2d1_hd U130 ( .A(n184), .B(N270), .Y(N271) );
  or2d1_hd U131 ( .A(n185), .B(N269), .Y(N270) );
  or2d1_hd U132 ( .A(n186), .B(N268), .Y(N269) );
  ad2d1_hd U133 ( .A(n72), .B(N241), .Y(N242) );
  ad2d1_hd U134 ( .A(n75), .B(N240), .Y(N241) );
  ad2d1_hd U135 ( .A(n78), .B(N239), .Y(N240) );
  ad2d1_hd U136 ( .A(n81), .B(N238), .Y(N239) );
  or2d1_hd U137 ( .A(n179), .B(N275), .Y(N276) );
  or2d1_hd U138 ( .A(n180), .B(N274), .Y(N275) );
  or2d1_hd U139 ( .A(n181), .B(N273), .Y(N274) );
  or2d1_hd U140 ( .A(n182), .B(N272), .Y(N273) );
  ad2d1_hd U141 ( .A(n60), .B(N245), .Y(N246) );
  ad2d1_hd U142 ( .A(n63), .B(N244), .Y(N245) );
  ad2d1_hd U143 ( .A(n66), .B(N243), .Y(N244) );
  ad2d1_hd U144 ( .A(n69), .B(N242), .Y(N243) );
  or2d1_hd U145 ( .A(n175), .B(N279), .Y(N280) );
  or2d1_hd U146 ( .A(n176), .B(N278), .Y(N279) );
  or2d1_hd U147 ( .A(n177), .B(N277), .Y(N278) );
  or2d1_hd U148 ( .A(n178), .B(N276), .Y(N277) );
  ad2d1_hd U149 ( .A(n48), .B(N249), .Y(N250) );
  ad2d1_hd U150 ( .A(n51), .B(N248), .Y(N249) );
  ad2d1_hd U151 ( .A(n54), .B(N247), .Y(N248) );
  ad2d1_hd U152 ( .A(n57), .B(N246), .Y(N247) );
  or2d1_hd U153 ( .A(n171), .B(N283), .Y(N284) );
  or2d1_hd U154 ( .A(n172), .B(N282), .Y(N283) );
  or2d1_hd U155 ( .A(n173), .B(N281), .Y(N282) );
  or2d1_hd U156 ( .A(n174), .B(N280), .Y(N281) );
  clknd2d1_hd U157 ( .A(n204), .B(N118), .Y(n206) );
  clknd2d1_hd U158 ( .A(n209), .B(n208), .Y(n211) );
  clknd2d1_hd U159 ( .A(n214), .B(n213), .Y(n217) );
  ad2d1_hd U160 ( .A(n36), .B(N253), .Y(N254) );
  ad2d1_hd U161 ( .A(n39), .B(N252), .Y(N253) );
  ad2d1_hd U162 ( .A(n42), .B(N251), .Y(N252) );
  ad2d1_hd U163 ( .A(n45), .B(N250), .Y(N251) );
  or2d1_hd U164 ( .A(n158), .B(n27), .Y(N309) );
  or2d1_hd U165 ( .A(n109), .B(sticky), .Y(N308) );
  clknd2d1_hd U166 ( .A(n226), .B(n225), .Y(n228) );
  nid2_hd U167 ( .A(n200), .Y(N6) );
  or2d1_hd U168 ( .A(n111), .B(n110), .Y(N230) );
  clknd2d1_hd U169 ( .A(n221), .B(n220), .Y(n223) );
  or2d1_hd U170 ( .A(n165), .B(N24), .Y(N31) );
  or2d1_hd U171 ( .A(N23), .B(n164), .Y(N37) );
  or2d1_hd U172 ( .A(n165), .B(N24), .Y(N34) );
  ivd1_hd U173 ( .A(n164), .Y(N24) );
  ivd1_hd U174 ( .A(n165), .Y(N23) );
  ivd1_hd U175 ( .A(n163), .Y(N25) );
  scg2d1_hd U176 ( .A(n234), .B(N81), .C(n233), .D(n6), .Y(value[30]) );
  scg2d1_hd U177 ( .A(n234), .B(N80), .C(n232), .D(n6), .Y(value[29]) );
  scg2d1_hd U178 ( .A(n234), .B(N51), .C(n167), .D(n6), .Y(value[0]) );
  scg2d1_hd U179 ( .A(n234), .B(N52), .C(n168), .D(n6), .Y(value[1]) );
  scg2d1_hd U180 ( .A(n234), .B(N53), .C(n169), .D(n6), .Y(value[2]) );
  scg2d1_hd U181 ( .A(n234), .B(N54), .C(n170), .D(n6), .Y(value[3]) );
  scg2d1_hd U182 ( .A(n234), .B(N55), .C(n171), .D(n6), .Y(value[4]) );
  scg2d1_hd U183 ( .A(n234), .B(N56), .C(n172), .D(n6), .Y(value[5]) );
  scg2d1_hd U184 ( .A(n234), .B(N57), .C(n173), .D(n6), .Y(value[6]) );
  scg2d1_hd U185 ( .A(n234), .B(N58), .C(n174), .D(n6), .Y(value[7]) );
  scg2d1_hd U186 ( .A(n234), .B(N59), .C(n175), .D(n6), .Y(value[8]) );
  scg2d1_hd U187 ( .A(n234), .B(N60), .C(n176), .D(n6), .Y(value[9]) );
  scg2d1_hd U188 ( .A(n234), .B(N61), .C(n177), .D(n6), .Y(value[10]) );
  scg2d1_hd U189 ( .A(n234), .B(N62), .C(n178), .D(n6), .Y(value[11]) );
  scg2d1_hd U190 ( .A(n234), .B(N63), .C(n179), .D(n6), .Y(value[12]) );
  scg2d1_hd U191 ( .A(n234), .B(N64), .C(n180), .D(n6), .Y(value[13]) );
  scg2d1_hd U192 ( .A(n234), .B(N65), .C(n181), .D(n6), .Y(value[14]) );
  scg2d1_hd U193 ( .A(n234), .B(N66), .C(n182), .D(n6), .Y(value[15]) );
  scg2d1_hd U194 ( .A(n234), .B(N67), .C(n183), .D(n6), .Y(value[16]) );
  scg2d1_hd U195 ( .A(n234), .B(N68), .C(n184), .D(n6), .Y(value[17]) );
  scg2d1_hd U196 ( .A(n234), .B(N69), .C(n185), .D(n6), .Y(value[18]) );
  scg2d1_hd U197 ( .A(n234), .B(N70), .C(n186), .D(n6), .Y(value[19]) );
  scg2d1_hd U198 ( .A(n234), .B(N71), .C(n187), .D(n6), .Y(value[20]) );
  scg2d1_hd U199 ( .A(n234), .B(N72), .C(n188), .D(n6), .Y(value[21]) );
  scg2d1_hd U200 ( .A(n234), .B(N73), .C(n189), .D(n6), .Y(value[22]) );
  scg2d1_hd U201 ( .A(n234), .B(N74), .C(n190), .D(n6), .Y(value[23]) );
  scg2d1_hd U202 ( .A(n234), .B(N75), .C(n191), .D(n6), .Y(value[24]) );
  scg2d1_hd U203 ( .A(n234), .B(N76), .C(n192), .D(n6), .Y(value[25]) );
  scg2d1_hd U204 ( .A(n234), .B(N77), .C(n193), .D(n6), .Y(value[26]) );
  scg2d1_hd U205 ( .A(n234), .B(N78), .C(n196), .D(n6), .Y(value[27]) );
  scg2d1_hd U206 ( .A(n234), .B(N79), .C(n197), .D(n6), .Y(value[28]) );
  clknd2d1_hd U207 ( .A(n16), .B(n203), .Y(z_e[0]) );
  clknd2d1_hd U208 ( .A(n15), .B(n203), .Y(z_e[1]) );
  clknd2d1_hd U209 ( .A(n14), .B(n203), .Y(z_e[2]) );
  clknd2d1_hd U210 ( .A(n13), .B(n203), .Y(z_e[3]) );
  clknd2d1_hd U211 ( .A(n11), .B(n203), .Y(z_e[4]) );
  clknd2d1_hd U212 ( .A(n10), .B(n8), .Y(z_e[5]) );
  clknd2d1_hd U213 ( .A(n9), .B(n8), .Y(z_e[6]) );
  clknd2d1_hd U214 ( .A(n7), .B(n8), .Y(z_e[7]) );
  xo2d1_hd U215 ( .A(n150), .B(n218), .Y(N125) );
  or2d1_hd U216 ( .A(n165), .B(n164), .Y(N28) );
  xo2d1_hd U217 ( .A(n150), .B(n231), .Y(n244) );
  clknd2d1_hd U218 ( .A(n215), .B(n230), .Y(n231) );
  scg2d1_hd U219 ( .A(n198), .B(n142), .C(N6), .D(n166), .Y(z_r[1]) );
  scg2d1_hd U220 ( .A(n198), .B(n141), .C(N6), .D(n114), .Y(z_r[2]) );
  scg2d1_hd U221 ( .A(n198), .B(n140), .C(N6), .D(n113), .Y(z_r[3]) );
  scg2d1_hd U222 ( .A(n198), .B(n139), .C(N6), .D(n112), .Y(z_r[4]) );
  scg2d1_hd U223 ( .A(n198), .B(n138), .C(N6), .D(n111), .Y(z_r[5]) );
  scg2d1_hd U224 ( .A(n198), .B(n137), .C(N6), .D(n110), .Y(z_r[6]) );
  scg2d1_hd U225 ( .A(n198), .B(n136), .C(N6), .D(n109), .Y(z_r[7]) );
  or2d1_hd U226 ( .A(n166), .B(N233), .Y(sticky) );
  or2d1_hd U227 ( .A(n114), .B(N232), .Y(N233) );
  or2d1_hd U228 ( .A(n113), .B(N231), .Y(N232) );
  or2d1_hd U229 ( .A(n112), .B(N230), .Y(N231) );
  or2d1_hd U230 ( .A(N23), .B(n164), .Y(N40) );
  or2d1_hd U231 ( .A(n198), .B(n201), .Y(N305) );
  or2d1_hd U233 ( .A(N23), .B(N24), .Y(N43) );
  ad2d1_hd U234 ( .A(N23), .B(N24), .Y(N26) );
  ad2d1_hd U235 ( .A(N26), .B(N25), .Y(N27) );
  ivd2_hd U237 ( .A(n234), .Y(n6) );
  nr2d1_hd U412 ( .A(n167), .B(N287), .Y(n194) );
  nr2d1_hd U413 ( .A(N28), .B(N25), .Y(n195) );
  clknd2d1_hd U414 ( .A(o_A_ACK), .B(i_A_STB), .Y(n242) );
  clknd2d1_hd U415 ( .A(o_Z_STB), .B(i_Z_ACK), .Y(n251) );
  nr2d4_hd U416 ( .A(N31), .B(n163), .Y(n198) );
  nr2d4_hd U417 ( .A(N37), .B(n163), .Y(n199) );
  nr2d1_hd U418 ( .A(N34), .B(N25), .Y(n200) );
  or4d1_hd U421 ( .A(n195), .B(n198), .C(n199), .D(n201), .Y(N293) );
  ad2d1_hd U422 ( .A(n107), .B(N309), .Y(N127) );
  nr2d1_hd U423 ( .A(n195), .B(n198), .Y(n203) );
  ivd1_hd U425 ( .A(n157), .Y(N118) );
  ivd1_hd U426 ( .A(n156), .Y(n204) );
  ao22d1_hd U427 ( .A(n156), .B(N118), .C(n157), .D(n204), .Y(N119) );
  ivd1_hd U428 ( .A(n206), .Y(n205) );
  ao22d1_hd U429 ( .A(n155), .B(n205), .C(n206), .D(n220), .Y(N120) );
  nr2d1_hd U430 ( .A(n155), .B(n206), .Y(n209) );
  ivd1_hd U431 ( .A(n209), .Y(n207) );
  ivd1_hd U432 ( .A(n154), .Y(n208) );
  ao22d1_hd U433 ( .A(n154), .B(n209), .C(n207), .D(n208), .Y(N121) );
  ivd1_hd U434 ( .A(n211), .Y(n210) );
  ao22d1_hd U435 ( .A(n153), .B(n210), .C(n211), .D(n225), .Y(N122) );
  nr2d1_hd U436 ( .A(n153), .B(n211), .Y(n214) );
  ivd1_hd U437 ( .A(n214), .Y(n212) );
  ivd1_hd U438 ( .A(n152), .Y(n213) );
  ao22d1_hd U439 ( .A(n152), .B(n214), .C(n212), .D(n213), .Y(N123) );
  ivd1_hd U440 ( .A(n217), .Y(n216) );
  ivd1_hd U441 ( .A(n151), .Y(n215) );
  ao22d1_hd U442 ( .A(n151), .B(n216), .C(n217), .D(n215), .Y(N124) );
  nr2d1_hd U443 ( .A(n151), .B(n217), .Y(n218) );
  ao22d1_hd U444 ( .A(n156), .B(N118), .C(n157), .D(n204), .Y(n250) );
  nr2d1_hd U445 ( .A(n156), .B(n157), .Y(n221) );
  ivd1_hd U446 ( .A(n221), .Y(n219) );
  ivd1_hd U447 ( .A(n155), .Y(n220) );
  ao22d1_hd U448 ( .A(n155), .B(n221), .C(n219), .D(n220), .Y(n249) );
  ivd1_hd U449 ( .A(n223), .Y(n222) );
  ao22d1_hd U450 ( .A(n154), .B(n222), .C(n223), .D(n208), .Y(n248) );
  nr2d1_hd U451 ( .A(n154), .B(n223), .Y(n226) );
  ivd1_hd U452 ( .A(n226), .Y(n224) );
  ivd1_hd U453 ( .A(n153), .Y(n225) );
  ao22d1_hd U454 ( .A(n153), .B(n226), .C(n224), .D(n225), .Y(n247) );
  ivd1_hd U455 ( .A(n228), .Y(n227) );
  ao22d1_hd U456 ( .A(n152), .B(n227), .C(n228), .D(n213), .Y(n246) );
  nr2d1_hd U457 ( .A(n152), .B(n228), .Y(n230) );
  ivd1_hd U458 ( .A(n230), .Y(n229) );
  ao22d1_hd U459 ( .A(n151), .B(n230), .C(n229), .D(n215), .Y(n245) );
  ivd1_hd U1 ( .A(i_RST), .Y(n12) );
  ivd1_hd U2 ( .A(i_RST), .Y(n21) );
  ivd1_hd U8 ( .A(i_RST), .Y(n22) );
  ivd1_hd U9 ( .A(i_RST), .Y(n23) );
  ivd1_hd U10 ( .A(i_RST), .Y(n24) );
  ivd6_hd U11 ( .A(n1) );
  ivd6_hd U12 ( .A(n2) );
  ivd6_hd U13 ( .A(n5) );
  ivd6_hd U14 ( .A(n4) );
  ivd6_hd U15 ( .A(n3) );
  fds2eqd1_hd clk_r_REG85_S3 ( .CRN(n23), .D(state_1_), .E(N180), .CK(i_CLK), 
        .Q(n164) );
  fd1eqd1_hd clk_r_REG107_S4 ( .D(z_e[0]), .E(N211), .CK(n256), .Q(n157) );
  fd1eqd1_hd clk_r_REG104_S4 ( .D(z_e[1]), .E(N211), .CK(n256), .Q(n156) );
  fd1eqd1_hd clk_r_REG101_S4 ( .D(z_e[2]), .E(N211), .CK(n256), .Q(n155) );
  fd1eqd1_hd clk_r_REG98_S4 ( .D(z_e[3]), .E(N211), .CK(n256), .Q(n154) );
  fd1eqd1_hd clk_r_REG95_S4 ( .D(z_e[4]), .E(N211), .CK(n256), .Q(n153) );
  fd1eqd1_hd clk_r_REG92_S4 ( .D(z_e[5]), .E(N211), .CK(n256), .Q(n152) );
  fd1eqd1_hd clk_r_REG89_S4 ( .D(z_e[6]), .E(N211), .CK(n256), .Q(n151) );
  fd1eqd1_hd clk_r_REG86_S4 ( .D(z_e[7]), .E(N211), .CK(n256), .Q(n150) );
  fd1eqd1_hd clk_r_REG61_S3 ( .D(z_m[23]), .E(N210), .CK(i_CLK), .Q(n94) );
  fd1eqd1_hd clk_r_REG15_S3 ( .D(z_m[0]), .E(N210), .CK(i_CLK), .Q(n27) );
  fd1qd1_hd clk_r_REG87_S5 ( .D(n244), .CK(n252), .Q(n149) );
  fd1qd1_hd clk_r_REG90_S5 ( .D(n245), .CK(n252), .Q(n96) );
  fd1qd1_hd clk_r_REG93_S5 ( .D(n246), .CK(n252), .Q(n98) );
  fd1qd1_hd clk_r_REG96_S5 ( .D(n247), .CK(n252), .Q(n100) );
  fd1qd1_hd clk_r_REG2_S3 ( .D(n162), .CK(n252), .Q(n161) );
  fd1qd1_hd clk_r_REG16_S4 ( .D(n27), .CK(n252), .Q(n26) );
  fd1qd1_hd clk_r_REG18_S4 ( .D(n30), .CK(n252), .Q(n29) );
  fd1qd1_hd clk_r_REG20_S4 ( .D(n33), .CK(n252), .Q(n32) );
  fd1qd1_hd clk_r_REG22_S4 ( .D(n36), .CK(n252), .Q(n35) );
  fd1qd1_hd clk_r_REG24_S4 ( .D(n39), .CK(n252), .Q(n38) );
  fd1qd1_hd clk_r_REG26_S4 ( .D(n42), .CK(n252), .Q(n41) );
  fd1qd1_hd clk_r_REG28_S4 ( .D(n45), .CK(n252), .Q(n44) );
  fd1qd1_hd clk_r_REG30_S4 ( .D(n48), .CK(n252), .Q(n47) );
  fd1qd1_hd clk_r_REG32_S4 ( .D(n51), .CK(n252), .Q(n50) );
  fd1qd1_hd clk_r_REG34_S4 ( .D(n54), .CK(n252), .Q(n53) );
  fd1qd1_hd clk_r_REG36_S4 ( .D(n57), .CK(n252), .Q(n56) );
  fd1qd1_hd clk_r_REG38_S4 ( .D(n60), .CK(n252), .Q(n59) );
  fd1qd1_hd clk_r_REG40_S4 ( .D(n63), .CK(n252), .Q(n62) );
  fd1qd1_hd clk_r_REG42_S4 ( .D(n66), .CK(n252), .Q(n65) );
  fd1qd1_hd clk_r_REG44_S4 ( .D(n69), .CK(n252), .Q(n68) );
  fd1qd1_hd clk_r_REG46_S4 ( .D(n72), .CK(n252), .Q(n71) );
  fd1qd1_hd clk_r_REG48_S4 ( .D(n75), .CK(n252), .Q(n74) );
  fd1qd1_hd clk_r_REG50_S4 ( .D(n78), .CK(n252), .Q(n77) );
  fd1qd1_hd clk_r_REG52_S4 ( .D(n81), .CK(n252), .Q(n80) );
  fd1qd1_hd clk_r_REG54_S4 ( .D(n84), .CK(n252), .Q(n83) );
  fd1qd1_hd clk_r_REG56_S4 ( .D(n87), .CK(n252), .Q(n86) );
  fd1qd1_hd clk_r_REG58_S4 ( .D(n90), .CK(n252), .Q(n89) );
  fd1qd1_hd clk_r_REG60_S4 ( .D(n93), .CK(n252), .Q(n92) );
  fd1qd1_hd clk_r_REG99_S5 ( .D(n248), .CK(n252), .Q(n102) );
  fd1qd1_hd clk_r_REG102_S5 ( .D(n249), .CK(n252), .Q(n104) );
  fd1qd1_hd clk_r_REG105_S5 ( .D(n250), .CK(n252), .Q(n106) );
  fd1qd1_hd clk_r_REG108_S5 ( .D(N118), .CK(n252), .Q(n236) );
  fd1qd1_hd clk_r_REG3_S4 ( .D(n161), .CK(n253), .Q(o_Z[31]) );
  fd1qd1_hd clk_r_REG62_S5 ( .D(n92), .CK(n253), .Q(o_Z[22]) );
  fd1qd1_hd clk_r_REG63_S5 ( .D(n89), .CK(n253), .Q(o_Z[21]) );
  fd1qd1_hd clk_r_REG64_S5 ( .D(n86), .CK(n253), .Q(o_Z[20]) );
  fd1qd1_hd clk_r_REG65_S5 ( .D(n83), .CK(n253), .Q(o_Z[19]) );
  fd1qd1_hd clk_r_REG66_S5 ( .D(n80), .CK(n253), .Q(o_Z[18]) );
  fd1qd1_hd clk_r_REG67_S5 ( .D(n77), .CK(n253), .Q(o_Z[17]) );
  fd1qd1_hd clk_r_REG68_S5 ( .D(n74), .CK(n253), .Q(o_Z[16]) );
  fd1qd1_hd clk_r_REG69_S5 ( .D(n71), .CK(n253), .Q(o_Z[15]) );
  fd1qd1_hd clk_r_REG70_S5 ( .D(n68), .CK(n253), .Q(o_Z[14]) );
  fd1qd1_hd clk_r_REG71_S5 ( .D(n65), .CK(n253), .Q(o_Z[13]) );
  fd1qd1_hd clk_r_REG72_S5 ( .D(n62), .CK(n253), .Q(o_Z[12]) );
  fd1qd1_hd clk_r_REG73_S5 ( .D(n59), .CK(n253), .Q(o_Z[11]) );
  fd1qd1_hd clk_r_REG74_S5 ( .D(n56), .CK(n253), .Q(o_Z[10]) );
  fd1qd1_hd clk_r_REG75_S5 ( .D(n53), .CK(n253), .Q(o_Z[9]) );
  fd1qd1_hd clk_r_REG76_S5 ( .D(n50), .CK(n253), .Q(o_Z[8]) );
  fd1qd1_hd clk_r_REG77_S5 ( .D(n47), .CK(n253), .Q(o_Z[7]) );
  fd1qd1_hd clk_r_REG78_S5 ( .D(n44), .CK(n253), .Q(o_Z[6]) );
  fd1qd1_hd clk_r_REG79_S5 ( .D(n41), .CK(n253), .Q(o_Z[5]) );
  fd1qd1_hd clk_r_REG80_S5 ( .D(n38), .CK(n253), .Q(o_Z[4]) );
  fd1qd1_hd clk_r_REG81_S5 ( .D(n35), .CK(n253), .Q(o_Z[3]) );
  fd1qd1_hd clk_r_REG82_S5 ( .D(n32), .CK(n253), .Q(o_Z[2]) );
  fd1qd1_hd clk_r_REG83_S5 ( .D(n29), .CK(n253), .Q(o_Z[1]) );
  fd1qd1_hd clk_r_REG84_S5 ( .D(n26), .CK(n253), .Q(o_Z[0]) );
  fd1qd1_hd clk_r_REG88_S6 ( .D(n149), .CK(n253), .Q(o_Z[30]) );
  fd1qd1_hd clk_r_REG91_S6 ( .D(n96), .CK(n253), .Q(o_Z[29]) );
  fd1qd1_hd clk_r_REG94_S6 ( .D(n98), .CK(n253), .Q(o_Z[28]) );
  fd1qd1_hd clk_r_REG97_S6 ( .D(n100), .CK(n253), .Q(o_Z[27]) );
  fd1qd1_hd clk_r_REG100_S6 ( .D(n102), .CK(n253), .Q(o_Z[26]) );
  fd1qd1_hd clk_r_REG103_S6 ( .D(n104), .CK(n253), .Q(o_Z[25]) );
  fd1qd1_hd clk_r_REG106_S6 ( .D(n106), .CK(n253), .Q(o_Z[24]) );
  fd1qd1_hd clk_r_REG109_S6 ( .D(n236), .CK(n253), .Q(o_Z[23]) );
  fd1qd1_hd clk_r_REG173_S1 ( .D(i_A[0]), .CK(n254), .Q(n167) );
  fd1qd1_hd clk_r_REG172_S1 ( .D(i_A[1]), .CK(n254), .Q(n168) );
  fd1qd1_hd clk_r_REG171_S1 ( .D(i_A[2]), .CK(n254), .Q(n169) );
  fd1qd1_hd clk_r_REG170_S1 ( .D(i_A[3]), .CK(n254), .Q(n170) );
  fd1qd1_hd clk_r_REG169_S1 ( .D(i_A[4]), .CK(n254), .Q(n171) );
  fd1qd1_hd clk_r_REG168_S1 ( .D(i_A[5]), .CK(n254), .Q(n172) );
  fd1qd1_hd clk_r_REG167_S1 ( .D(i_A[6]), .CK(n254), .Q(n173) );
  fd1qd1_hd clk_r_REG166_S1 ( .D(i_A[7]), .CK(n254), .Q(n174) );
  fd1qd1_hd clk_r_REG165_S1 ( .D(i_A[8]), .CK(n254), .Q(n175) );
  fd1qd1_hd clk_r_REG164_S1 ( .D(i_A[9]), .CK(n254), .Q(n176) );
  fd1qd1_hd clk_r_REG163_S1 ( .D(i_A[10]), .CK(n254), .Q(n177) );
  fd1qd1_hd clk_r_REG162_S1 ( .D(i_A[11]), .CK(n254), .Q(n178) );
  fd1qd1_hd clk_r_REG161_S1 ( .D(i_A[12]), .CK(n254), .Q(n179) );
  fd1qd1_hd clk_r_REG160_S1 ( .D(i_A[13]), .CK(n254), .Q(n180) );
  fd1qd1_hd clk_r_REG159_S1 ( .D(i_A[14]), .CK(n254), .Q(n181) );
  fd1qd1_hd clk_r_REG158_S1 ( .D(i_A[15]), .CK(n254), .Q(n182) );
  fd1qd1_hd clk_r_REG157_S1 ( .D(i_A[16]), .CK(n254), .Q(n183) );
  fd1qd1_hd clk_r_REG156_S1 ( .D(i_A[17]), .CK(n254), .Q(n184) );
  fd1qd1_hd clk_r_REG155_S1 ( .D(i_A[18]), .CK(n254), .Q(n185) );
  fd1qd1_hd clk_r_REG154_S1 ( .D(i_A[19]), .CK(n254), .Q(n186) );
  fd1qd1_hd clk_r_REG153_S1 ( .D(i_A[20]), .CK(n254), .Q(n187) );
  fd1qd1_hd clk_r_REG152_S1 ( .D(i_A[21]), .CK(n254), .Q(n188) );
  fd1qd1_hd clk_r_REG151_S1 ( .D(i_A[22]), .CK(n254), .Q(n189) );
  fd1qd1_hd clk_r_REG150_S1 ( .D(i_A[23]), .CK(n254), .Q(n190) );
  fd1qd1_hd clk_r_REG149_S1 ( .D(i_A[24]), .CK(n254), .Q(n191) );
  fd1qd1_hd clk_r_REG148_S1 ( .D(i_A[25]), .CK(n254), .Q(n192) );
  fd1qd1_hd clk_r_REG147_S1 ( .D(i_A[26]), .CK(n254), .Q(n193) );
  fd1qd1_hd clk_r_REG146_S1 ( .D(i_A[27]), .CK(n254), .Q(n196) );
  fd1qd1_hd clk_r_REG145_S1 ( .D(i_A[28]), .CK(n254), .Q(n197) );
  fd1qd1_hd clk_r_REG144_S1 ( .D(i_A[29]), .CK(n254), .Q(n232) );
  fd1qd1_hd clk_r_REG143_S1 ( .D(i_A[30]), .CK(n254), .Q(n233) );
  fd1qd2_hd clk_r_REG0_S1 ( .D(i_A[31]), .CK(n254), .Q(n234) );
  fd1qd1_hd clk_r_REG141_S2 ( .D(value[28]), .CK(n255), .Q(n115) );
  fd1qd1_hd clk_r_REG140_S2 ( .D(value[27]), .CK(n255), .Q(n116) );
  fd1qd1_hd clk_r_REG139_S2 ( .D(value[26]), .CK(n255), .Q(n117) );
  fd1qd1_hd clk_r_REG138_S2 ( .D(value[25]), .CK(n255), .Q(n118) );
  fd1qd1_hd clk_r_REG137_S2 ( .D(value[24]), .CK(n255), .Q(n119) );
  fd1qd1_hd clk_r_REG136_S2 ( .D(value[23]), .CK(n255), .Q(n120) );
  fd1qd1_hd clk_r_REG135_S2 ( .D(value[22]), .CK(n255), .Q(n121) );
  fd1qd1_hd clk_r_REG134_S2 ( .D(value[21]), .CK(n255), .Q(n122) );
  fd1qd1_hd clk_r_REG133_S2 ( .D(value[20]), .CK(n255), .Q(n123) );
  fd1qd1_hd clk_r_REG132_S2 ( .D(value[19]), .CK(n255), .Q(n124) );
  fd1qd1_hd clk_r_REG131_S2 ( .D(value[18]), .CK(n255), .Q(n125) );
  fd1qd1_hd clk_r_REG130_S2 ( .D(value[17]), .CK(n255), .Q(n126) );
  fd1qd1_hd clk_r_REG129_S2 ( .D(value[16]), .CK(n255), .Q(n127) );
  fd1qd1_hd clk_r_REG128_S2 ( .D(value[15]), .CK(n255), .Q(n128) );
  fd1qd1_hd clk_r_REG127_S2 ( .D(value[14]), .CK(n255), .Q(n129) );
  fd1qd1_hd clk_r_REG126_S2 ( .D(value[13]), .CK(n255), .Q(n130) );
  fd1qd1_hd clk_r_REG125_S2 ( .D(value[12]), .CK(n255), .Q(n131) );
  fd1qd1_hd clk_r_REG124_S2 ( .D(value[11]), .CK(n255), .Q(n132) );
  fd1qd1_hd clk_r_REG123_S2 ( .D(value[10]), .CK(n255), .Q(n133) );
  fd1qd1_hd clk_r_REG122_S2 ( .D(value[9]), .CK(n255), .Q(n134) );
  fd1qd1_hd clk_r_REG121_S2 ( .D(value[8]), .CK(n255), .Q(n135) );
  fd1qd1_hd clk_r_REG120_S2 ( .D(value[7]), .CK(n255), .Q(n136) );
  fd1qd1_hd clk_r_REG119_S2 ( .D(value[6]), .CK(n255), .Q(n137) );
  fd1qd1_hd clk_r_REG118_S2 ( .D(value[5]), .CK(n255), .Q(n138) );
  fd1qd1_hd clk_r_REG117_S2 ( .D(value[4]), .CK(n255), .Q(n139) );
  fd1qd1_hd clk_r_REG116_S2 ( .D(value[3]), .CK(n255), .Q(n140) );
  fd1qd1_hd clk_r_REG115_S2 ( .D(value[2]), .CK(n255), .Q(n141) );
  fd1qd1_hd clk_r_REG114_S2 ( .D(value[1]), .CK(n255), .Q(n142) );
  fd1qd1_hd clk_r_REG113_S2 ( .D(value[0]), .CK(n255), .Q(n143) );
  fd1qd1_hd clk_r_REG112_S2 ( .D(value[29]), .CK(n255), .Q(n144) );
  fd1qd1_hd clk_r_REG111_S2 ( .D(value[30]), .CK(n255), .Q(n145) );
  fd1qd1_hd clk_r_REG142_S2 ( .D(value[31]), .CK(n255), .Q(n159) );
  fd1qd1_hd clk_r_REG17_S3 ( .D(z_m[1]), .CK(n256), .Q(n30) );
  fd1qd1_hd clk_r_REG19_S3 ( .D(z_m[2]), .CK(n256), .Q(n33) );
  fd1qd1_hd clk_r_REG21_S3 ( .D(z_m[3]), .CK(n256), .Q(n36) );
  fd1qd1_hd clk_r_REG23_S3 ( .D(z_m[4]), .CK(n256), .Q(n39) );
  fd1qd1_hd clk_r_REG25_S3 ( .D(z_m[5]), .CK(n256), .Q(n42) );
  fd1qd1_hd clk_r_REG27_S3 ( .D(z_m[6]), .CK(n256), .Q(n45) );
  fd1qd1_hd clk_r_REG29_S3 ( .D(z_m[7]), .CK(n256), .Q(n48) );
  fd1qd1_hd clk_r_REG31_S3 ( .D(z_m[8]), .CK(n256), .Q(n51) );
  fd1qd1_hd clk_r_REG33_S3 ( .D(z_m[9]), .CK(n256), .Q(n54) );
  fd1qd1_hd clk_r_REG35_S3 ( .D(z_m[10]), .CK(n256), .Q(n57) );
  fd1qd1_hd clk_r_REG37_S3 ( .D(z_m[11]), .CK(n256), .Q(n60) );
  fd1qd1_hd clk_r_REG39_S3 ( .D(z_m[12]), .CK(n256), .Q(n63) );
  fd1qd1_hd clk_r_REG41_S3 ( .D(z_m[13]), .CK(n256), .Q(n66) );
  fd1qd1_hd clk_r_REG43_S3 ( .D(z_m[14]), .CK(n256), .Q(n69) );
  fd1qd1_hd clk_r_REG45_S3 ( .D(z_m[15]), .CK(n256), .Q(n72) );
  fd1qd1_hd clk_r_REG47_S3 ( .D(z_m[16]), .CK(n256), .Q(n75) );
  fd1qd1_hd clk_r_REG49_S3 ( .D(z_m[17]), .CK(n256), .Q(n78) );
  fd1qd1_hd clk_r_REG51_S3 ( .D(z_m[18]), .CK(n256), .Q(n81) );
  fd1qd1_hd clk_r_REG53_S3 ( .D(z_m[19]), .CK(n256), .Q(n84) );
  fd1qd1_hd clk_r_REG55_S3 ( .D(z_m[20]), .CK(n256), .Q(n87) );
  fd1qd1_hd clk_r_REG57_S3 ( .D(z_m[21]), .CK(n256), .Q(n90) );
  fd1qd1_hd clk_r_REG59_S3 ( .D(z_m[22]), .CK(n256), .Q(n93) );
  fd1qd1_hd clk_r_REG13_S3 ( .D(z_r[7]), .CK(n257), .Q(n108) );
  fd1qd1_hd clk_r_REG12_S3 ( .D(z_r[6]), .CK(n257), .Q(n109) );
  fd1qd1_hd clk_r_REG11_S3 ( .D(z_r[5]), .CK(n257), .Q(n110) );
  fd1qd1_hd clk_r_REG9_S3 ( .D(z_r[4]), .CK(n257), .Q(n111) );
  fd1qd1_hd clk_r_REG8_S3 ( .D(z_r[3]), .CK(n257), .Q(n112) );
  fd1qd1_hd clk_r_REG7_S3 ( .D(z_r[2]), .CK(n257), .Q(n113) );
  fd1qd1_hd clk_r_REG6_S3 ( .D(z_r[1]), .CK(n257), .Q(n114) );
  fd1qd1_hd clk_r_REG5_S3 ( .D(z_r[0]), .CK(n257), .Q(n166) );
  fd1eqd1_hd clk_r_REG110_S2 ( .D(n264), .E(n279), .CK(i_CLK), .Q(n163) );
  fd1eqd1_hd clk_r_REG174_S1 ( .D(n262), .E(n281), .CK(i_CLK), .Q(o_A_ACK) );
  fd1eqd1_hd clk_r_REG175_S1 ( .D(n260), .E(n283), .CK(i_CLK), .Q(o_Z_STB) );
  fd1eqd1_hd clk_r_REG1_S2 ( .D(n243), .E(n195), .CK(i_CLK), .Q(n162) );
  fd1eqd1_hd clk_r_REG4_S2 ( .D(n258), .E(n285), .CK(i_CLK), .Q(n165) );
  fd1eqd1_hd clk_r_REG14_S4 ( .D(n108), .E(N229), .CK(i_CLK), .Q(n107) );
  fd1eqd1_hd clk_r_REG10_S4 ( .D(N308), .E(N229), .CK(i_CLK), .Q(n158) );
  converter_i2f_DW01_inc_0 add_x_4 ( .A({n150, n151, n152, n153, n154, n155, 
        n156, n157}), .SUM({N161, N160, N159, N158, N157, N156, N155, N154})
         );
  converter_i2f_DW01_inc_1 add_x_3 ( .A({n94, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, n36, 
        n33, n30, n27}), .SUM({N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, 
        N133, N132, N131, N130}) );
  converter_i2f_DW01_sub_0 sub_x_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({n234, n233, n232, n197, n196, n193, n192, n191, n190, 
        n189, n188, n187, n186, n185, n184, n183, n182, n181, n180, n179, n178, 
        n177, n176, n175, n174, n173, n172, n171, n170, n169, n168, n167}), 
        .CI(1'b0), .DIFF({N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55, N54, N53, N52, N51}) );
  SNPS_CLOCK_GATE_HIGH_converter_i2f_12 clk_gate_clk_r_REG13_S3_0 ( .CLK(i_CLK), .EN(N220), .ENCLK(n257), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_i2f_13 clk_gate_clk_r_REG17_S3_0 ( .CLK(i_CLK), .EN(N210), .ENCLK(n256), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_i2f_14 clk_gate_clk_r_REG141_S2_0 ( .CLK(
        i_CLK), .EN(N185), .ENCLK(n255), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_i2f_15 clk_gate_clk_r_REG173_S1_0 ( .CLK(
        i_CLK), .EN(N184), .ENCLK(n254), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_i2f_16 clk_gate_clk_r_REG3_S4_0 ( .CLK(i_CLK), 
        .EN(n202), .ENCLK(n253), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_i2f_17 clk_gate_clk_r_REG87_S5_0 ( .CLK(i_CLK), .EN(n201), .ENCLK(n252), .TE(1'b0) );
  clknd2d1_hd U16 ( .A(n19), .B(n163), .Y(n268) );
  clknd2d1_hd U17 ( .A(n164), .B(N23), .Y(n274) );
  clknd2d1_hd U18 ( .A(N24), .B(n242), .Y(n272) );
  nr2d1_hd U19 ( .A(N40), .B(N25), .Y(n201) );
  nr2d1_hd U20 ( .A(N43), .B(n163), .Y(n202) );
  nr2bd1_hd U21 ( .AN(N27), .B(n242), .Y(N184) );
  nr2d1_hd U22 ( .A(n194), .B(n8), .Y(N185) );
  clknd2d1_hd U23 ( .A(n164), .B(n277), .Y(n276) );
  clknd2d1_hd U24 ( .A(n163), .B(n194), .Y(n275) );
  ivd1_hd U25 ( .A(n259), .Y(n258) );
  clknd2d1_hd U26 ( .A(n24), .B(n284), .Y(n259) );
  ivd1_hd U27 ( .A(n261), .Y(n260) );
  clknd2d1_hd U28 ( .A(n12), .B(n282), .Y(n261) );
  ivd1_hd U29 ( .A(n263), .Y(n262) );
  clknd2d1_hd U30 ( .A(n21), .B(n280), .Y(n263) );
  ivd1_hd U31 ( .A(n265), .Y(n264) );
  clknd2d1_hd U33 ( .A(n22), .B(n278), .Y(n265) );
  scg13d1_hd U35 ( .A(N220), .B(n17), .C(n18), .Y(N210) );
  scg9d1_hd U37 ( .A(n266), .B(n267), .C(n22), .Y(n278) );
  ao211d1_hd U39 ( .A(n164), .B(n268), .C(n165), .D(n269), .Y(n267) );
  ao21d1_hd U41 ( .A(n194), .B(n270), .C(n164), .Y(n269) );
  ivd1_hd U43 ( .A(n242), .Y(n270) );
  nr2d1_hd U45 ( .A(n271), .B(n163), .Y(n266) );
  oa22d1_hd U47 ( .A(n165), .B(n272), .C(N23), .D(N24), .Y(n271) );
  oa211d1_hd U48 ( .A(n164), .B(n273), .C(n22), .D(n274), .Y(n279) );
  scg12d1_hd U51 ( .A(n242), .B(n194), .C(n165), .Y(n273) );
  ad2d1_hd U78 ( .A(n242), .B(n21), .Y(n280) );
  nd2bd1_hd U80 ( .AN(N27), .B(n21), .Y(n281) );
  ad2d1_hd U82 ( .A(n251), .B(n12), .Y(n282) );
  nd2bd1_hd U83 ( .AN(n202), .B(n12), .Y(n283) );
  ad2d1_hd U86 ( .A(n163), .B(n24), .Y(n284) );
  oa211d1_hd U91 ( .A(n164), .B(n275), .C(n24), .D(n276), .Y(n285) );
  ao22d1_hd U92 ( .A(n163), .B(n19), .C(n251), .D(N25), .Y(n277) );
endmodule


module float_adder_DW01_inc_0 ( A, SUM );
  input [23:0] A;
  output [23:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;

  had1_hd U2 ( .A(A[22]), .B(n2), .CO(n1), .S(SUM[22]) );
  had1_hd U3 ( .A(A[21]), .B(n3), .CO(n2), .S(SUM[21]) );
  had1_hd U4 ( .A(A[20]), .B(n4), .CO(n3), .S(SUM[20]) );
  had1_hd U5 ( .A(A[19]), .B(n5), .CO(n4), .S(SUM[19]) );
  had1_hd U6 ( .A(A[18]), .B(n6), .CO(n5), .S(SUM[18]) );
  had1_hd U7 ( .A(A[17]), .B(n7), .CO(n6), .S(SUM[17]) );
  had1_hd U8 ( .A(A[16]), .B(n8), .CO(n7), .S(SUM[16]) );
  had1_hd U9 ( .A(A[15]), .B(n9), .CO(n8), .S(SUM[15]) );
  had1_hd U10 ( .A(A[14]), .B(n10), .CO(n9), .S(SUM[14]) );
  had1_hd U11 ( .A(A[13]), .B(n11), .CO(n10), .S(SUM[13]) );
  had1_hd U12 ( .A(A[12]), .B(n12), .CO(n11), .S(SUM[12]) );
  had1_hd U13 ( .A(A[11]), .B(n13), .CO(n12), .S(SUM[11]) );
  had1_hd U14 ( .A(A[10]), .B(n14), .CO(n13), .S(SUM[10]) );
  had1_hd U15 ( .A(A[9]), .B(n15), .CO(n14), .S(SUM[9]) );
  had1_hd U16 ( .A(A[8]), .B(n16), .CO(n15), .S(SUM[8]) );
  had1_hd U17 ( .A(A[7]), .B(n17), .CO(n16), .S(SUM[7]) );
  had1_hd U18 ( .A(A[6]), .B(n18), .CO(n17), .S(SUM[6]) );
  had1_hd U19 ( .A(A[5]), .B(n19), .CO(n18), .S(SUM[5]) );
  had1_hd U20 ( .A(A[4]), .B(n20), .CO(n19), .S(SUM[4]) );
  had1_hd U21 ( .A(A[3]), .B(n21), .CO(n20), .S(SUM[3]) );
  had1_hd U22 ( .A(A[2]), .B(n22), .CO(n21), .S(SUM[2]) );
  had1_hd U23 ( .A(A[1]), .B(A[0]), .CO(n22), .S(SUM[1]) );
  xo2d1_hd U27 ( .A(n1), .B(A[23]), .Y(SUM[23]) );
  ivd1_hd U28 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module float_adder_DP_OP_131_125_8359_0 ( I1, O1, U488_Y, i_CLK, IN0 );
  input [7:0] I1;
  output [8:0] O1;
  input U488_Y, i_CLK, IN0;
  wire   n2, n3, n4, n5, n6, n7, n29, n30, n1, n8, n9, n10, n11, n12, n13, n14
;

  had1_hd U4 ( .A(n13), .B(n3), .CO(n2), .S(O1[6]) );
  had1_hd U5 ( .A(n12), .B(n4), .CO(n3), .S(O1[5]) );
  had1_hd U6 ( .A(n11), .B(n5), .CO(n4), .S(O1[4]) );
  had1_hd U7 ( .A(n10), .B(n6), .CO(n5), .S(O1[3]) );
  had1_hd U8 ( .A(n9), .B(n7), .CO(n6), .S(O1[2]) );
  had1_hd U9 ( .A(n8), .B(n1), .CO(n7), .S(O1[1]) );
  nr2d1_hd U13 ( .A(n14), .B(n2), .Y(O1[8]) );
  ao22d1_hd U14 ( .A(n14), .B(n29), .C(n2), .D(n30), .Y(O1[7]) );
  ivd1_hd U15 ( .A(n14), .Y(n30) );
  ivd1_hd U16 ( .A(n2), .Y(n29) );
  ivd1_hd U17 ( .A(n1), .Y(O1[0]) );
  fd1qd1_hd clk_r_REG247_S1 ( .D(I1[7]), .CK(IN0), .Q(n14) );
  fd1qd1_hd clk_r_REG248_S1 ( .D(I1[6]), .CK(IN0), .Q(n13) );
  fd1qd1_hd clk_r_REG249_S1 ( .D(I1[5]), .CK(IN0), .Q(n12) );
  fd1qd1_hd clk_r_REG250_S1 ( .D(I1[4]), .CK(IN0), .Q(n11) );
  fd1qd1_hd clk_r_REG251_S1 ( .D(I1[3]), .CK(IN0), .Q(n10) );
  fd1qd1_hd clk_r_REG252_S1 ( .D(I1[2]), .CK(IN0), .Q(n9) );
  fd1qd1_hd clk_r_REG253_S1 ( .D(I1[1]), .CK(IN0), .Q(n8) );
  fd1qd1_hd clk_r_REG254_S1 ( .D(I1[0]), .CK(IN0), .Q(n1) );
endmodule


module float_adder_DP_OP_132_126_1283_0 ( I1, O1 );
  input [9:0] I1;
  output [9:0] O1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  had1_hd U2 ( .A(I1[8]), .B(n2), .CO(n1), .S(O1[8]) );
  had1_hd U3 ( .A(I1[7]), .B(n3), .CO(n2), .S(O1[7]) );
  had1_hd U4 ( .A(I1[6]), .B(n4), .CO(n3), .S(O1[6]) );
  had1_hd U5 ( .A(I1[5]), .B(n5), .CO(n4), .S(O1[5]) );
  had1_hd U6 ( .A(I1[4]), .B(n6), .CO(n5), .S(O1[4]) );
  had1_hd U7 ( .A(I1[3]), .B(n7), .CO(n6), .S(O1[3]) );
  had1_hd U8 ( .A(I1[2]), .B(n8), .CO(n7), .S(O1[2]) );
  had1_hd U9 ( .A(I1[1]), .B(I1[0]), .CO(n8), .S(O1[1]) );
  xo2d1_hd U13 ( .A(I1[9]), .B(n1), .Y(O1[9]) );
  ivd1_hd U14 ( .A(I1[0]), .Y(O1[0]) );
endmodule


module float_adder_DP_OP_128_128_163_0 ( I1, O1, U488_Y, i_CLK, IN0 );
  input [7:0] I1;
  output [8:0] O1;
  input U488_Y, i_CLK, IN0;
  wire   n2, n3, n4, n5, n6, n7, n29, n30, n1, n8, n9, n10, n11, n12, n13, n14
;

  had1_hd U4 ( .A(n13), .B(n3), .CO(n2), .S(O1[6]) );
  had1_hd U5 ( .A(n12), .B(n4), .CO(n3), .S(O1[5]) );
  had1_hd U6 ( .A(n11), .B(n5), .CO(n4), .S(O1[4]) );
  had1_hd U7 ( .A(n10), .B(n6), .CO(n5), .S(O1[3]) );
  had1_hd U8 ( .A(n9), .B(n7), .CO(n6), .S(O1[2]) );
  had1_hd U9 ( .A(n8), .B(n1), .CO(n7), .S(O1[1]) );
  nr2d1_hd U13 ( .A(n14), .B(n2), .Y(O1[8]) );
  ao22d1_hd U14 ( .A(n14), .B(n29), .C(n2), .D(n30), .Y(O1[7]) );
  ivd1_hd U15 ( .A(n14), .Y(n30) );
  ivd1_hd U16 ( .A(n2), .Y(n29) );
  ivd1_hd U17 ( .A(n1), .Y(O1[0]) );
  fd1qd1_hd clk_r_REG122_S1 ( .D(I1[7]), .CK(IN0), .Q(n14) );
  fd1qd1_hd clk_r_REG215_S1 ( .D(I1[6]), .CK(IN0), .Q(n13) );
  fd1qd1_hd clk_r_REG216_S1 ( .D(I1[5]), .CK(IN0), .Q(n12) );
  fd1qd1_hd clk_r_REG217_S1 ( .D(I1[4]), .CK(IN0), .Q(n11) );
  fd1qd1_hd clk_r_REG218_S1 ( .D(I1[3]), .CK(IN0), .Q(n10) );
  fd1qd1_hd clk_r_REG219_S1 ( .D(I1[2]), .CK(IN0), .Q(n9) );
  fd1qd1_hd clk_r_REG220_S1 ( .D(I1[1]), .CK(IN0), .Q(n8) );
  fd1qd1_hd clk_r_REG221_S1 ( .D(I1[0]), .CK(IN0), .Q(n1) );
endmodule


module float_adder_DP_OP_129_129_1948_0 ( I1, O1 );
  input [9:0] I1;
  output [9:0] O1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  had1_hd U2 ( .A(I1[8]), .B(n2), .CO(n1), .S(O1[8]) );
  had1_hd U3 ( .A(I1[7]), .B(n3), .CO(n2), .S(O1[7]) );
  had1_hd U4 ( .A(I1[6]), .B(n4), .CO(n3), .S(O1[6]) );
  had1_hd U5 ( .A(I1[5]), .B(n5), .CO(n4), .S(O1[5]) );
  had1_hd U6 ( .A(I1[4]), .B(n6), .CO(n5), .S(O1[4]) );
  had1_hd U7 ( .A(I1[3]), .B(n7), .CO(n6), .S(O1[3]) );
  had1_hd U8 ( .A(I1[2]), .B(n8), .CO(n7), .S(O1[2]) );
  had1_hd U9 ( .A(I1[1]), .B(I1[0]), .CO(n8), .S(O1[1]) );
  xo2d1_hd U13 ( .A(I1[9]), .B(n1), .Y(O1[9]) );
  ivd1_hd U14 ( .A(I1[0]), .Y(O1[0]) );
endmodule


module float_adder_DP_OP_143_130_3257_0 ( I1, I2, O1 );
  input [9:0] I1;
  output [9:0] O1;
  input I2;
  wire   n2, n3, n4, n5, n6, n7, n8, n9;

  fad1_hd U3 ( .A(I2), .B(I1[8]), .CI(n3), .CO(n2), .S(O1[8]) );
  fad1_hd U4 ( .A(I2), .B(I1[7]), .CI(n4), .CO(n3), .S(O1[7]) );
  fad1_hd U5 ( .A(I2), .B(I1[6]), .CI(n5), .CO(n4), .S(O1[6]) );
  fad1_hd U6 ( .A(I2), .B(I1[5]), .CI(n6), .CO(n5), .S(O1[5]) );
  fad1_hd U7 ( .A(I2), .B(I1[4]), .CI(n7), .CO(n6), .S(O1[4]) );
  fad1_hd U8 ( .A(I2), .B(I1[3]), .CI(n8), .CO(n7), .S(O1[3]) );
  fad1_hd U9 ( .A(I2), .B(I1[2]), .CI(n9), .CO(n8), .S(O1[2]) );
  fad1_hd U10 ( .A(I2), .B(I1[1]), .CI(I1[0]), .CO(n9), .S(O1[1]) );
  xo3d1_hd U14 ( .A(n2), .B(I1[9]), .C(I2), .Y(O1[9]) );
  ivd1_hd U15 ( .A(I1[0]), .Y(O1[0]) );
endmodule


module float_adder_DP_OP_43_133_2142_0 ( I1, I2, I3, O1 );
  input [26:0] I1;
  input [26:0] I2;
  output [27:0] O1;
  input I3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n142;

  xo2d1_hd U59 ( .A(I3), .B(I2[3]), .Y(n55) );
  xo2d1_hd U60 ( .A(I3), .B(I2[10]), .Y(n48) );
  xo2d1_hd U61 ( .A(I3), .B(I2[5]), .Y(n53) );
  ivd1_hd U62 ( .A(I3), .Y(n142) );
  fad4_hd U65 ( .A(n41), .B(I1[17]), .CI(n11), .CO(n10), .S(O1[17]) );
  fad4_hd U70 ( .A(n44), .B(I1[14]), .CI(n14), .CO(n13), .S(O1[14]) );
  fad4_hd U72 ( .A(n39), .B(I1[19]), .CI(n9), .CO(n8), .S(O1[19]) );
  fad4_hd U77 ( .A(n33), .B(I1[25]), .CI(n3), .CO(n2), .S(O1[25]) );
  xo2d1_hd U80 ( .A(I3), .B(I2[12]), .Y(n46) );
  xo2d1_hd U81 ( .A(I3), .B(I2[19]), .Y(n39) );
  xo2d1_hd U82 ( .A(I3), .B(I2[9]), .Y(n49) );
  xo2d1_hd U84 ( .A(I3), .B(I2[26]), .Y(n32) );
  xo2d1_hd U85 ( .A(I3), .B(I2[25]), .Y(n33) );
  xo2d1_hd U86 ( .A(I3), .B(I2[24]), .Y(n34) );
  xo2d1_hd U87 ( .A(I3), .B(I2[23]), .Y(n35) );
  xo2d1_hd U89 ( .A(I3), .B(I2[22]), .Y(n36) );
  xo2d1_hd U91 ( .A(I3), .B(I2[21]), .Y(n37) );
  xo2d1_hd U93 ( .A(I3), .B(I2[20]), .Y(n38) );
  xo2d1_hd U94 ( .A(I3), .B(I2[18]), .Y(n40) );
  xo2d1_hd U95 ( .A(I3), .B(I2[17]), .Y(n41) );
  xo2d1_hd U96 ( .A(I3), .B(I2[16]), .Y(n42) );
  xo2d1_hd U98 ( .A(I3), .B(I2[15]), .Y(n43) );
  xo2d1_hd U99 ( .A(I3), .B(I2[14]), .Y(n44) );
  xo2d1_hd U100 ( .A(I3), .B(I2[13]), .Y(n45) );
  xo2d1_hd U101 ( .A(I3), .B(I2[11]), .Y(n47) );
  xo2d1_hd U102 ( .A(I3), .B(I2[8]), .Y(n50) );
  xo2d1_hd U103 ( .A(I3), .B(I2[7]), .Y(n51) );
  xo2d1_hd U104 ( .A(I3), .B(I2[6]), .Y(n52) );
  xo2d1_hd U105 ( .A(I3), .B(I2[4]), .Y(n54) );
  xo2d1_hd U106 ( .A(I3), .B(I2[2]), .Y(n56) );
  xo2d1_hd U107 ( .A(I3), .B(I2[1]), .Y(n57) );
  fad2_hd U108 ( .A(n54), .B(I1[4]), .CI(n24), .CO(n23), .S(O1[4]) );
  fad4_hd U110 ( .A(n48), .B(I1[10]), .CI(n18), .CO(n17), .S(O1[10]) );
  fad4_hd U3 ( .A(n35), .B(I1[23]), .CI(n5), .CO(n4), .S(O1[23]) );
  xo2d4_hd U5 ( .A(I3), .B(I2[0]), .Y(n58) );
  fad4_hd U6 ( .A(n36), .B(I1[22]), .CI(n6), .CO(n5), .S(O1[22]) );
  fad2_hd U8 ( .A(n32), .B(I1[26]), .CI(n2), .CO(n1), .S(O1[26]) );
  fad2_hd U9 ( .A(n42), .B(I1[16]), .CI(n12), .CO(n11), .S(O1[16]) );
  fad2_hd U10 ( .A(n45), .B(I1[13]), .CI(n15), .CO(n14), .S(O1[13]) );
  fad2_hd U11 ( .A(n47), .B(I1[11]), .CI(n17), .CO(n16), .S(O1[11]) );
  fad2_hd U13 ( .A(n51), .B(I1[7]), .CI(n21), .CO(n20), .S(O1[7]) );
  fad4_hd U16 ( .A(n57), .B(I1[1]), .CI(n27), .CO(n26), .S(O1[1]) );
  fad2_hd U17 ( .A(I1[0]), .B(I3), .CI(n58), .CO(n27), .S(O1[0]) );
  fad2_hd U1 ( .A(n55), .B(I1[3]), .CI(n25), .CO(n24), .S(O1[3]) );
  fad2_hd U2 ( .A(n40), .B(I1[18]), .CI(n10), .CO(n9), .S(O1[18]) );
  fad4_hd U4 ( .A(n52), .B(I1[6]), .CI(n22), .CO(n21), .S(O1[6]) );
  fad4_hd U7 ( .A(n53), .B(I1[5]), .CI(n23), .CO(n22), .S(O1[5]) );
  fad4_hd U12 ( .A(n56), .B(I1[2]), .CI(n26), .CO(n25), .S(O1[2]) );
  fad4_hd U14 ( .A(n34), .B(I1[24]), .CI(n4), .CO(n3), .S(O1[24]) );
  fad4_hd U15 ( .A(n37), .B(I1[21]), .CI(n7), .CO(n6), .S(O1[21]) );
  fad4_hd U18 ( .A(n38), .B(I1[20]), .CI(n8), .CO(n7), .S(O1[20]) );
  fad4_hd U19 ( .A(n49), .B(I1[9]), .CI(n19), .CO(n18), .S(O1[9]) );
  fad4_hd U20 ( .A(n50), .B(I1[8]), .CI(n20), .CO(n19), .S(O1[8]) );
  fad1_hd U21 ( .A(n46), .B(I1[12]), .CI(n16), .CO(n15), .S(O1[12]) );
  fad1_hd U22 ( .A(n43), .B(I1[15]), .CI(n13), .CO(n12), .S(O1[15]) );
  xn2d1_hd U23 ( .A(n142), .B(n1), .Y(O1[27]) );
endmodule


module float_adder_DW_cmp_6 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE, 
        U780_Y, i_CLK, U786_Y, IN0, IN1, IN2 );
  input [26:0] A;
  input [26:0] B;
  input TC, GE_LT, GE_GT_EQ, U780_Y, i_CLK, U786_Y, IN0, IN1, IN2;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n199, n200,
         n201, n202, n11;

  nr2bd1_hd U140 ( .AN(B[1]), .B(A[1]), .Y(n101) );
  nd2bd1_hd U141 ( .AN(B[1]), .B(A[1]), .Y(n102) );
  nr2bd1_hd U142 ( .AN(B[2]), .B(A[2]), .Y(n98) );
  nr2bd1_hd U143 ( .AN(B[3]), .B(A[3]), .Y(n96) );
  nd2bd1_hd U144 ( .AN(B[2]), .B(A[2]), .Y(n99) );
  nd2bd1_hd U145 ( .AN(B[3]), .B(A[3]), .Y(n97) );
  clknd2d1_hd U146 ( .A(n201), .B(n199), .Y(n8) );
  oa21d1_hd U147 ( .A(n103), .B(n101), .C(n102), .Y(n100) );
  nr2bd1_hd U148 ( .AN(B[0]), .B(A[0]), .Y(n103) );
  nr2d1_hd U149 ( .A(n98), .B(n96), .Y(n94) );
  oa21d1_hd U150 ( .A(n96), .B(n99), .C(n97), .Y(n95) );
  nr2d1_hd U151 ( .A(n91), .B(n89), .Y(n87) );
  nr2d1_hd U152 ( .A(n112), .B(A[4]), .Y(n91) );
  nr2d1_hd U153 ( .A(n113), .B(A[5]), .Y(n89) );
  oa21d1_hd U154 ( .A(n89), .B(n92), .C(n90), .Y(n88) );
  ao21d1_hd U157 ( .A(n100), .B(n94), .C(n95), .Y(n93) );
  clknd2d1_hd U158 ( .A(n72), .B(n66), .Y(n64) );
  ao21d1_hd U160 ( .A(n66), .B(n73), .C(n67), .Y(n65) );
  nr2d1_hd U161 ( .A(n116), .B(A[8]), .Y(n76) );
  clknd2d1_hd U162 ( .A(n112), .B(A[4]), .Y(n92) );
  or2d1_hd U163 ( .A(n132), .B(A[24]), .Y(n201) );
  nr2d1_hd U164 ( .A(n76), .B(n74), .Y(n72) );
  nr2d1_hd U165 ( .A(n11), .B(IN2), .Y(n6) );
  nr2d1_hd U167 ( .A(n125), .B(A[17]), .Y(n44) );
  nr2d1_hd U168 ( .A(n117), .B(A[9]), .Y(n74) );
  clknd2d1_hd U169 ( .A(n113), .B(A[5]), .Y(n90) );
  ad2d1_hd U170 ( .A(n133), .B(A[25]), .Y(n202) );
  nr2d1_hd U171 ( .A(n56), .B(n54), .Y(n52) );
  clknd2d1_hd U172 ( .A(n11), .B(IN2), .Y(n7) );
  ao21d1_hd U173 ( .A(n199), .B(n200), .C(n202), .Y(n9) );
  oa21d1_hd U174 ( .A(n9), .B(n6), .C(n7), .Y(n5) );
  ivd1_hd U177 ( .A(B[23]), .Y(n131) );
  ivd1_hd U178 ( .A(B[19]), .Y(n127) );
  ivd1_hd U179 ( .A(B[21]), .Y(n129) );
  ivd1_hd U180 ( .A(B[22]), .Y(n130) );
  ivd1_hd U181 ( .A(B[5]), .Y(n113) );
  ivd1_hd U182 ( .A(B[7]), .Y(n115) );
  ivd1_hd U183 ( .A(B[4]), .Y(n112) );
  ivd1_hd U184 ( .A(B[6]), .Y(n114) );
  nr2d1_hd U185 ( .A(n115), .B(A[7]), .Y(n83) );
  ivd1_hd U186 ( .A(B[15]), .Y(n123) );
  ivd1_hd U187 ( .A(B[11]), .Y(n119) );
  ivd1_hd U188 ( .A(B[13]), .Y(n121) );
  ivd1_hd U189 ( .A(B[14]), .Y(n122) );
  ivd1_hd U190 ( .A(B[9]), .Y(n117) );
  ivd1_hd U191 ( .A(B[10]), .Y(n118) );
  nr2d1_hd U192 ( .A(n119), .B(A[11]), .Y(n68) );
  ivd1_hd U193 ( .A(B[12]), .Y(n120) );
  nr2d1_hd U194 ( .A(n121), .B(A[13]), .Y(n60) );
  ivd1_hd U195 ( .A(B[17]), .Y(n125) );
  ivd1_hd U196 ( .A(B[18]), .Y(n126) );
  nr2d1_hd U197 ( .A(n127), .B(A[19]), .Y(n38) );
  ivd1_hd U198 ( .A(B[20]), .Y(n128) );
  nr2d1_hd U199 ( .A(n129), .B(A[21]), .Y(n30) );
  ivd1_hd U200 ( .A(B[25]), .Y(n133) );
  ad2d1_hd U201 ( .A(n132), .B(A[24]), .Y(n200) );
  ivd1_hd U202 ( .A(B[26]), .Y(n134) );
  clknd2d1_hd U203 ( .A(n130), .B(A[22]), .Y(n27) );
  clknd2d1_hd U204 ( .A(n131), .B(A[23]), .Y(n25) );
  nr2d1_hd U205 ( .A(n131), .B(A[23]), .Y(n24) );
  oa21d1_hd U206 ( .A(n44), .B(n47), .C(n45), .Y(n43) );
  clknd2d1_hd U207 ( .A(n125), .B(A[17]), .Y(n45) );
  clknd2d1_hd U208 ( .A(n124), .B(A[16]), .Y(n47) );
  oa21d1_hd U209 ( .A(n38), .B(n41), .C(n39), .Y(n37) );
  clknd2d1_hd U210 ( .A(n127), .B(A[19]), .Y(n39) );
  clknd2d1_hd U211 ( .A(n126), .B(A[18]), .Y(n41) );
  oa21d1_hd U212 ( .A(n30), .B(n33), .C(n31), .Y(n29) );
  clknd2d1_hd U213 ( .A(n129), .B(A[21]), .Y(n31) );
  clknd2d1_hd U214 ( .A(n128), .B(A[20]), .Y(n33) );
  nr2d1_hd U215 ( .A(n26), .B(n24), .Y(n22) );
  nr2d1_hd U216 ( .A(n130), .B(A[22]), .Y(n26) );
  oa21d1_hd U217 ( .A(n83), .B(n86), .C(n84), .Y(n82) );
  clknd2d1_hd U218 ( .A(n115), .B(A[7]), .Y(n84) );
  clknd2d1_hd U219 ( .A(n114), .B(A[6]), .Y(n86) );
  nr2d1_hd U221 ( .A(n114), .B(A[6]), .Y(n85) );
  clknd2d1_hd U222 ( .A(n122), .B(A[14]), .Y(n57) );
  clknd2d1_hd U223 ( .A(n123), .B(A[15]), .Y(n55) );
  nr2d1_hd U224 ( .A(n123), .B(A[15]), .Y(n54) );
  oa21d1_hd U225 ( .A(n74), .B(n77), .C(n75), .Y(n73) );
  clknd2d1_hd U226 ( .A(n117), .B(A[9]), .Y(n75) );
  clknd2d1_hd U227 ( .A(n116), .B(A[8]), .Y(n77) );
  oa21d1_hd U228 ( .A(n68), .B(n71), .C(n69), .Y(n67) );
  clknd2d1_hd U229 ( .A(n119), .B(A[11]), .Y(n69) );
  clknd2d1_hd U230 ( .A(n118), .B(A[10]), .Y(n71) );
  oa21d1_hd U231 ( .A(n60), .B(n63), .C(n61), .Y(n59) );
  clknd2d1_hd U232 ( .A(n121), .B(A[13]), .Y(n61) );
  clknd2d1_hd U233 ( .A(n120), .B(A[12]), .Y(n63) );
  nr2d1_hd U234 ( .A(n122), .B(A[14]), .Y(n56) );
  ivd1_hd U235 ( .A(B[8]), .Y(n116) );
  nr2d1_hd U236 ( .A(n70), .B(n68), .Y(n66) );
  nr2d1_hd U237 ( .A(n118), .B(A[10]), .Y(n70) );
  nr2d1_hd U238 ( .A(n62), .B(n60), .Y(n58) );
  nr2d1_hd U239 ( .A(n120), .B(A[12]), .Y(n62) );
  ivd1_hd U240 ( .A(B[24]), .Y(n132) );
  ivd1_hd U241 ( .A(B[16]), .Y(n124) );
  nr2d1_hd U242 ( .A(n40), .B(n38), .Y(n36) );
  nr2d1_hd U243 ( .A(n126), .B(A[18]), .Y(n40) );
  nr2d1_hd U244 ( .A(n32), .B(n30), .Y(n28) );
  nr2d1_hd U245 ( .A(n128), .B(A[20]), .Y(n32) );
  oa21d1_hd U246 ( .A(n35), .B(n20), .C(n21), .Y(n19) );
  ao21d1_hd U247 ( .A(n22), .B(n29), .C(n23), .Y(n21) );
  ao21d1_hd U248 ( .A(n36), .B(n43), .C(n37), .Y(n35) );
  oa21d1_hd U249 ( .A(n24), .B(n27), .C(n25), .Y(n23) );
  ao21d1_hd U250 ( .A(n52), .B(n59), .C(n53), .Y(n51) );
  oa21d1_hd U251 ( .A(n54), .B(n57), .C(n55), .Y(n53) );
  nr2d1_hd U252 ( .A(n34), .B(n20), .Y(n18) );
  clknd2d1_hd U253 ( .A(n42), .B(n36), .Y(n34) );
  nr2d1_hd U254 ( .A(n46), .B(n44), .Y(n42) );
  nr2d1_hd U255 ( .A(n124), .B(A[16]), .Y(n46) );
  or2d1_hd U256 ( .A(n133), .B(A[25]), .Y(n199) );
  nr2d1_hd U1 ( .A(n85), .B(n83), .Y(n81) );
  clknd2d1_hd U2 ( .A(n58), .B(n52), .Y(n50) );
  clknd2d1_hd U3 ( .A(n28), .B(n22), .Y(n20) );
  oa21d1_hd U4 ( .A(n65), .B(n50), .C(n51), .Y(n49) );
  oa21d1_hd U5 ( .A(n93), .B(n79), .C(n80), .Y(n78) );
  clknd2d1_hd U6 ( .A(n87), .B(n81), .Y(n79) );
  ao21d1_hd U7 ( .A(n81), .B(n88), .C(n82), .Y(n80) );
  nr2d1_hd U8 ( .A(n64), .B(n50), .Y(n48) );
  nr2d1_hd U9 ( .A(n8), .B(n6), .Y(n4) );
  ao21d1_hd U12 ( .A(n19), .B(n4), .C(n5), .Y(n3) );
  fd1qd1_hd clk_r_REG212_S5 ( .D(n134), .CK(IN1), .Q(n11) );
  ao21d1_hd U10 ( .A(n78), .B(n48), .C(n49), .Y(n1) );
  oa21d2_hd U11 ( .A(n1), .B(n2), .C(n3), .Y(GE_LT_GT_LE) );
  nd2d1_hd U13 ( .A(n18), .B(n4), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_12_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_10_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_9_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_7_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_4_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_3_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_2_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_1_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_adder_0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module float_adder ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n695,
         n728, guard, round_bit, sticky, z_s, N47, N87, N220, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N443,
         N444, N445, N446, N447, N448, N449, N450, N511, N516, N543, N545,
         N573, N574, N585, N596, N629, N664, N667, N668, C85_DATA2_0,
         C85_DATA2_1, C85_DATA2_2, C85_DATA2_3, C85_DATA2_4, C85_DATA2_5,
         C85_DATA2_6, C85_DATA2_7, C85_DATA2_8, C85_DATA2_9, C82_DATA2_0,
         C82_DATA2_1, C82_DATA2_2, C82_DATA2_3, C82_DATA2_4, C82_DATA2_5,
         C82_DATA2_6, C82_DATA2_7, n6, n7, n8, n9, n10, n11, C1_DATA1_8,
         C1_DATA1_7, C1_DATA1_6, C1_DATA1_5, C1_DATA1_4, C1_DATA1_3,
         C1_DATA1_2, C1_DATA1_1, C1_DATA1_0, C1_DATA2_9, C1_DATA2_8,
         C1_DATA2_7, C1_DATA2_6, C1_DATA2_5, C1_DATA2_4, C1_DATA2_3,
         C1_DATA2_2, C1_DATA2_1, C1_DATA2_0, C2_Z_26, C2_Z_25, C2_Z_24,
         C2_Z_23, C2_Z_22, C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17,
         C2_Z_16, C2_Z_15, C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9,
         C2_Z_8, C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1,
         C2_Z_0, C3_Z_26, C3_Z_25, C3_Z_24, C3_Z_23, C3_Z_22, C3_Z_21, C3_Z_20,
         C3_Z_19, C3_Z_18, C3_Z_17, C3_Z_16, C3_Z_15, C3_Z_14, C3_Z_13,
         C3_Z_12, C3_Z_11, C3_Z_10, C3_Z_9, C3_Z_8, C3_Z_7, C3_Z_6, C3_Z_5,
         C3_Z_4, C3_Z_3, C3_Z_2, C3_Z_1, C3_Z_0, C1_Z_7, C1_Z_6, C1_Z_5,
         C1_Z_4, C1_Z_3, C1_Z_2, C1_Z_1, C1_Z_0, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n176, n177, n179, n182, n183, n185, n186,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n401, n402, n403,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n1, n2, n3, n4, n5,
         n12, n13, n14, n15, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n134, n136, n138, n140, n142, n144, n146, n148,
         n150, n152, n154, n156, n158, n160, n162, n164, n166, n168, n170,
         n172, n187, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n589, n591, n593, n595, n597, n599,
         n601, n603, n605, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n743, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n789, n795;
  wire   [3:0] state;
  wire   [8:0] a_e;
  wire   [25:0] a_m;
  wire   [9:0] b_e;
  wire   [25:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;

  ivd1_hd U26 ( .A(i_RST), .Y(n6) );
  ivd1_hd U27 ( .A(i_RST), .Y(n7) );
  ivd1_hd U28 ( .A(i_RST), .Y(n8) );
  ivd1_hd U29 ( .A(i_RST), .Y(n9) );
  ivd1_hd U30 ( .A(i_RST), .Y(n10) );
  ivd1_hd U31 ( .A(i_RST), .Y(n11) );
  mx2id1_hd U261 ( .D0(n384), .D1(n491), .S(n486), .YN(C3_Z_5) );
  mx2id1_hd U262 ( .D0(n388), .D1(n419), .S(n486), .YN(C3_Z_3) );
  or2d1_hd U263 ( .A(n130), .B(n426), .Y(n84) );
  mx2id1_hd U264 ( .D0(n374), .D1(n510), .S(n486), .YN(C3_Z_10) );
  mx2id1_hd U265 ( .D0(n510), .D1(n374), .S(n486), .YN(C2_Z_10) );
  mx2id1_hd U266 ( .D0(n491), .D1(n384), .S(n486), .YN(C2_Z_5) );
  nr2d1_hd U267 ( .A(n130), .B(n428), .Y(N543) );
  mx2id1_hd U269 ( .D0(n508), .D1(n370), .S(n486), .YN(C2_Z_12) );
  mx2id1_hd U270 ( .D0(n370), .D1(n508), .S(n486), .YN(C3_Z_12) );
  clknd2d1_hd U271 ( .A(n191), .B(n190), .Y(n194) );
  clknd2d1_hd U272 ( .A(n197), .B(n196), .Y(n200) );
  clknd2d1_hd U273 ( .A(n203), .B(n202), .Y(n204) );
  mx2id1_hd U276 ( .D0(n501), .D1(n356), .S(n486), .YN(C2_Z_19) );
  mx2id1_hd U277 ( .D0(n356), .D1(n501), .S(n486), .YN(C3_Z_19) );
  mx2id1_hd U278 ( .D0(n487), .D1(n376), .S(n486), .YN(C2_Z_9) );
  mx2id1_hd U279 ( .D0(n376), .D1(n487), .S(n486), .YN(C3_Z_9) );
  clknd2d1_hd U280 ( .A(n430), .B(n315), .Y(n519) );
  clknd2d1_hd U281 ( .A(n458), .B(n459), .Y(n457) );
  clknd2d1_hd U282 ( .A(n113), .B(n112), .Y(n436) );
  clknd2d1_hd U283 ( .A(n585), .B(n473), .Y(n461) );
  clknd2d1_hd U284 ( .A(n582), .B(n475), .Y(n450) );
  clknd2d1_hd U285 ( .A(n127), .B(n474), .Y(n468) );
  clknd2d1_hd U286 ( .A(n583), .B(n480), .Y(n456) );
  clknd2d1_hd U287 ( .A(n132), .B(n448), .Y(n445) );
  clknd2d1_hd U288 ( .A(n587), .B(n481), .Y(n478) );
  clknd2d1_hd U289 ( .A(n18), .B(n479), .Y(n441) );
  clknd2d1_hd U290 ( .A(n423), .B(n424), .Y(n315) );
  clknd2d1_hd U291 ( .A(n410), .B(n343), .Y(n518) );
  clknd2d1_hd U292 ( .A(n523), .B(n524), .Y(n344) );
  clknd2d1_hd U293 ( .A(n438), .B(n425), .Y(n413) );
  clknd2d1_hd U294 ( .A(n434), .B(n484), .Y(n485) );
  clknd2d2_hd U295 ( .A(N543), .B(n392), .Y(n334) );
  clknd2d1_hd U296 ( .A(n208), .B(n207), .Y(n211) );
  clknd2d1_hd U297 ( .A(n214), .B(n213), .Y(n217) );
  clknd2d1_hd U298 ( .A(n220), .B(n219), .Y(n221) );
  clknd2d1_hd U299 ( .A(n333), .B(n334), .Y(n321) );
  clknd2d1_hd U300 ( .A(n223), .B(n636), .Y(n230) );
  clknd2d1_hd U301 ( .A(n280), .B(n281), .Y(n279) );
  ivd1_hd U302 ( .A(N220), .Y(n186) );
  scg13d1_hd U303 ( .A(n511), .B(n185), .C(n186), .Y(n183) );
  ivd1_hd U304 ( .A(n541), .Y(n185) );
  or2d1_hd U305 ( .A(n512), .B(n541), .Y(n176) );
  ad2d1_hd U308 ( .A(n661), .B(n565), .Y(n177) );
  nr2d1_hd U309 ( .A(n661), .B(n565), .Y(n182) );
  ivd1_hd U310 ( .A(n565), .Y(n313) );
  ivd1_hd U311 ( .A(n661), .Y(n311) );
  ivd2_hd U312 ( .A(N543), .Y(n293) );
  scg2d1_hd U313 ( .A(n393), .B(C1_DATA2_7), .C(n660), .D(C1_DATA1_7), .Y(
        a_e[7]) );
  scg2d1_hd U314 ( .A(n393), .B(n549), .C(n660), .D(n559), .Y(b_e[7]) );
  scg2d1_hd U315 ( .A(n66), .B(n741), .C(C85_DATA2_0), .D(n279), .Y(z_e[0]) );
  scg2d1_hd U316 ( .A(n581), .B(n741), .C(C85_DATA2_1), .D(n279), .Y(z_e[1])
         );
  scg2d1_hd U317 ( .A(n580), .B(n741), .C(C85_DATA2_2), .D(n279), .Y(z_e[2])
         );
  scg2d1_hd U318 ( .A(n579), .B(n741), .C(C85_DATA2_3), .D(n279), .Y(z_e[3])
         );
  scg2d1_hd U319 ( .A(n578), .B(n741), .C(C85_DATA2_4), .D(n279), .Y(z_e[4])
         );
  scg2d1_hd U320 ( .A(n577), .B(n741), .C(C85_DATA2_5), .D(n279), .Y(z_e[5])
         );
  scg2d1_hd U321 ( .A(n119), .B(n393), .C(n660), .D(n637), .Y(b_m[3]) );
  scg2d1_hd U322 ( .A(n118), .B(n393), .C(n660), .D(n638), .Y(b_m[4]) );
  scg2d1_hd U323 ( .A(n64), .B(n393), .C(n660), .D(n639), .Y(b_m[5]) );
  scg2d1_hd U324 ( .A(n116), .B(n393), .C(n660), .D(n663), .Y(a_m[3]) );
  scg2d1_hd U325 ( .A(n115), .B(n393), .C(n660), .D(n664), .Y(a_m[4]) );
  scg2d1_hd U326 ( .A(n110), .B(n393), .C(n660), .D(n665), .Y(a_m[5]) );
  clknd2d1_hd U327 ( .A(n226), .B(n227), .Y(N668) );
  clknd2d1_hd U328 ( .A(n429), .B(n85), .Y(state[0]) );
  clknd2d1_hd U329 ( .A(i_Z_ACK), .B(o_Z_STB), .Y(n728) );
  mx2id1_hd U331 ( .D0(n688), .D1(n687), .S(n486), .YN(C2_Z_26) );
  mx2id1_hd U332 ( .D0(n687), .D1(n688), .S(n486), .YN(C3_Z_26) );
  mx2id1_hd U333 ( .D0(n495), .D1(n345), .S(n486), .YN(C2_Z_25) );
  mx2id1_hd U334 ( .D0(n345), .D1(n495), .S(n486), .YN(C3_Z_25) );
  mx2id1_hd U335 ( .D0(n496), .D1(n346), .S(n486), .YN(C2_Z_24) );
  mx2id1_hd U336 ( .D0(n346), .D1(n496), .S(n486), .YN(C3_Z_24) );
  clknd2d1_hd U337 ( .A(n296), .B(n565), .Y(n295) );
  clknd2d1_hd U338 ( .A(n328), .B(n319), .Y(n704) );
  clknd2d1_hd U339 ( .A(n327), .B(n319), .Y(n703) );
  clknd2d1_hd U340 ( .A(n326), .B(n319), .Y(n702) );
  clknd2d1_hd U341 ( .A(n325), .B(n319), .Y(n701) );
  clknd2d1_hd U342 ( .A(n324), .B(n319), .Y(n700) );
  clknd2d1_hd U343 ( .A(n323), .B(n319), .Y(n699) );
  clknd2d1_hd U344 ( .A(n322), .B(n319), .Y(n698) );
  clknd2d1_hd U345 ( .A(n318), .B(n319), .Y(n697) );
  xo2d1_hd U346 ( .A(n113), .B(n221), .Y(N450) );
  xo2d1_hd U347 ( .A(C1_Z_7), .B(n204), .Y(C82_DATA2_7) );
  scg2d1_hd U348 ( .A(n576), .B(n741), .C(C85_DATA2_6), .D(n279), .Y(z_e[6])
         );
  scg2d1_hd U349 ( .A(n128), .B(n741), .C(C85_DATA2_7), .D(n279), .Y(z_e[7])
         );
  scg2d1_hd U350 ( .A(n131), .B(n741), .C(C85_DATA2_8), .D(n279), .Y(z_e[8])
         );
  scg2d1_hd U351 ( .A(n18), .B(n741), .C(C85_DATA2_9), .D(n279), .Y(z_e[9]) );
  mx2id1_hd U352 ( .D0(n497), .D1(n348), .S(n486), .YN(C2_Z_23) );
  mx2id1_hd U353 ( .D0(n348), .D1(n497), .S(n486), .YN(C3_Z_23) );
  mx2id1_hd U354 ( .D0(n498), .D1(n350), .S(n486), .YN(C2_Z_22) );
  mx2id1_hd U355 ( .D0(n350), .D1(n498), .S(n486), .YN(C3_Z_22) );
  mx2id1_hd U356 ( .D0(n499), .D1(n352), .S(n486), .YN(C2_Z_21) );
  mx2id1_hd U357 ( .D0(n352), .D1(n499), .S(n486), .YN(C3_Z_21) );
  mx2id1_hd U358 ( .D0(n500), .D1(n354), .S(n486), .YN(C2_Z_20) );
  mx2id1_hd U359 ( .D0(n354), .D1(n500), .S(n486), .YN(C3_Z_20) );
  mx2id1_hd U360 ( .D0(n502), .D1(n358), .S(n486), .YN(C2_Z_18) );
  mx2id1_hd U361 ( .D0(n358), .D1(n502), .S(n486), .YN(C3_Z_18) );
  mx2id1_hd U362 ( .D0(n503), .D1(n360), .S(n486), .YN(C2_Z_17) );
  mx2id1_hd U363 ( .D0(n360), .D1(n503), .S(n486), .YN(C3_Z_17) );
  mx2id1_hd U364 ( .D0(n504), .D1(n362), .S(n486), .YN(C2_Z_16) );
  mx2id1_hd U365 ( .D0(n362), .D1(n504), .S(n486), .YN(C3_Z_16) );
  mx2id1_hd U366 ( .D0(n505), .D1(n364), .S(n486), .YN(C2_Z_15) );
  mx2id1_hd U367 ( .D0(n364), .D1(n505), .S(n486), .YN(C3_Z_15) );
  mx2id1_hd U368 ( .D0(n506), .D1(n366), .S(n486), .YN(C2_Z_14) );
  mx2id1_hd U369 ( .D0(n366), .D1(n506), .S(n486), .YN(C3_Z_14) );
  mx2id1_hd U370 ( .D0(n507), .D1(n368), .S(n486), .YN(C2_Z_13) );
  mx2id1_hd U371 ( .D0(n368), .D1(n507), .S(n486), .YN(C3_Z_13) );
  mx2id1_hd U372 ( .D0(n509), .D1(n372), .S(n486), .YN(C2_Z_11) );
  mx2id1_hd U373 ( .D0(n372), .D1(n509), .S(n486), .YN(C3_Z_11) );
  mx2id1_hd U374 ( .D0(n488), .D1(n378), .S(n486), .YN(C2_Z_8) );
  mx2id1_hd U375 ( .D0(n378), .D1(n488), .S(n486), .YN(C3_Z_8) );
  mx2id1_hd U376 ( .D0(n489), .D1(n380), .S(n486), .YN(C2_Z_7) );
  mx2id1_hd U377 ( .D0(n380), .D1(n489), .S(n486), .YN(C3_Z_7) );
  mx2id1_hd U378 ( .D0(n490), .D1(n382), .S(n486), .YN(C2_Z_6) );
  mx2id1_hd U379 ( .D0(n382), .D1(n490), .S(n486), .YN(C3_Z_6) );
  mx2id1_hd U380 ( .D0(n492), .D1(n386), .S(n486), .YN(C2_Z_4) );
  mx2id1_hd U381 ( .D0(n386), .D1(n492), .S(n486), .YN(C3_Z_4) );
  mx2id1_hd U382 ( .D0(n420), .D1(n414), .S(n486), .YN(C2_Z_2) );
  mx2id1_hd U383 ( .D0(n414), .D1(n420), .S(n486), .YN(C3_Z_2) );
  mx2id1_hd U384 ( .D0(n511), .D1(n512), .S(n486), .YN(C2_Z_1) );
  oa211d1_hd U385 ( .A(n186), .B(n512), .C(n183), .D(n176), .Y(C3_Z_1) );
  mx2id1_hd U386 ( .D0(n313), .D1(n311), .S(n486), .YN(z_s) );
  scg2d1_hd U387 ( .A(n109), .B(n393), .C(n660), .D(n666), .Y(a_m[6]) );
  scg2d1_hd U388 ( .A(n108), .B(n393), .C(n660), .D(n667), .Y(a_m[7]) );
  scg2d1_hd U389 ( .A(n83), .B(n393), .C(n660), .D(n668), .Y(a_m[8]) );
  scg2d1_hd U390 ( .A(n82), .B(n393), .C(n660), .D(n669), .Y(a_m[9]) );
  scg2d1_hd U391 ( .A(n81), .B(n393), .C(n660), .D(n670), .Y(a_m[10]) );
  scg2d1_hd U392 ( .A(n80), .B(n393), .C(n660), .D(n671), .Y(a_m[11]) );
  scg2d1_hd U393 ( .A(n79), .B(n393), .C(n660), .D(n672), .Y(a_m[12]) );
  scg2d1_hd U394 ( .A(n78), .B(n393), .C(n660), .D(n673), .Y(a_m[13]) );
  scg2d1_hd U395 ( .A(n77), .B(n393), .C(n660), .D(n674), .Y(a_m[14]) );
  scg2d1_hd U396 ( .A(n76), .B(n393), .C(n660), .D(n675), .Y(a_m[15]) );
  scg2d1_hd U397 ( .A(n75), .B(n393), .C(n660), .D(n676), .Y(a_m[16]) );
  scg2d1_hd U398 ( .A(n74), .B(n393), .C(n660), .D(n677), .Y(a_m[17]) );
  scg2d1_hd U399 ( .A(n73), .B(n393), .C(n660), .D(n678), .Y(a_m[18]) );
  scg2d1_hd U400 ( .A(n72), .B(n393), .C(n660), .D(n679), .Y(a_m[19]) );
  scg2d1_hd U401 ( .A(n71), .B(n393), .C(n660), .D(n680), .Y(a_m[20]) );
  scg2d1_hd U402 ( .A(n70), .B(n393), .C(n660), .D(n681), .Y(a_m[21]) );
  scg2d1_hd U403 ( .A(n69), .B(n393), .C(n660), .D(n682), .Y(a_m[22]) );
  scg2d1_hd U404 ( .A(n68), .B(n393), .C(n660), .D(n683), .Y(a_m[23]) );
  scg2d1_hd U405 ( .A(n67), .B(n393), .C(n660), .D(n684), .Y(a_m[24]) );
  scg2d1_hd U407 ( .A(n743), .B(n393), .C(n660), .D(n685), .Y(a_m[25]) );
  scg2d1_hd U408 ( .A(n393), .B(C1_DATA2_0), .C(n660), .D(C1_DATA1_0), .Y(
        a_e[0]) );
  scg2d1_hd U409 ( .A(n393), .B(n542), .C(n660), .D(n552), .Y(b_e[0]) );
  scg2d1_hd U410 ( .A(n63), .B(n393), .C(n660), .D(n640), .Y(b_m[6]) );
  scg2d1_hd U411 ( .A(n62), .B(n393), .C(n660), .D(n641), .Y(b_m[7]) );
  scg2d1_hd U412 ( .A(n61), .B(n393), .C(n660), .D(n642), .Y(b_m[8]) );
  scg2d1_hd U413 ( .A(n60), .B(n393), .C(n660), .D(n643), .Y(b_m[9]) );
  scg2d1_hd U414 ( .A(n59), .B(n393), .C(n660), .D(n644), .Y(b_m[10]) );
  scg2d1_hd U415 ( .A(n58), .B(n393), .C(n660), .D(n645), .Y(b_m[11]) );
  scg2d1_hd U416 ( .A(n57), .B(n393), .C(n660), .D(n646), .Y(b_m[12]) );
  scg2d1_hd U417 ( .A(n56), .B(n393), .C(n660), .D(n647), .Y(b_m[13]) );
  scg2d1_hd U418 ( .A(n55), .B(n393), .C(n660), .D(n648), .Y(b_m[14]) );
  scg2d1_hd U419 ( .A(n54), .B(n393), .C(n660), .D(n649), .Y(b_m[15]) );
  scg2d1_hd U420 ( .A(n53), .B(n393), .C(n660), .D(n650), .Y(b_m[16]) );
  scg2d1_hd U421 ( .A(n52), .B(n393), .C(n660), .D(n651), .Y(b_m[17]) );
  scg2d1_hd U422 ( .A(n51), .B(n393), .C(n660), .D(n652), .Y(b_m[18]) );
  scg2d1_hd U423 ( .A(n50), .B(n393), .C(n660), .D(n653), .Y(b_m[19]) );
  scg2d1_hd U424 ( .A(n49), .B(n393), .C(n660), .D(n654), .Y(b_m[20]) );
  scg2d1_hd U425 ( .A(n48), .B(n393), .C(n660), .D(n655), .Y(b_m[21]) );
  scg2d1_hd U426 ( .A(n47), .B(n393), .C(n660), .D(n656), .Y(b_m[22]) );
  scg2d1_hd U427 ( .A(n46), .B(n393), .C(n660), .D(n657), .Y(b_m[23]) );
  scg2d1_hd U428 ( .A(n45), .B(n393), .C(n660), .D(n658), .Y(b_m[24]) );
  scg2d1_hd U430 ( .A(n607), .B(n393), .C(n660), .D(n659), .Y(b_m[25]) );
  or2d1_hd U431 ( .A(n425), .B(n428), .Y(n85) );
  or2d1_hd U432 ( .A(n636), .B(n226), .Y(n86) );
  ao22d1_hd U433 ( .A(n393), .B(C1_DATA2_4), .C(n660), .D(C1_DATA1_4), .Y(n87)
         );
  ao22d1_hd U434 ( .A(n393), .B(C1_DATA2_5), .C(n660), .D(C1_DATA1_5), .Y(n88)
         );
  ao22d1_hd U435 ( .A(n393), .B(C1_DATA2_6), .C(n660), .D(C1_DATA1_6), .Y(n89)
         );
  oa21d2_hd U436 ( .A(n408), .B(n402), .C(n409), .Y(N574) );
  oa211d2_hd U438 ( .A(n229), .B(n85), .C(n282), .D(n227), .Y(N629) );
  ad2d2_hd U439 ( .A(n299), .B(n331), .Y(n339) );
  ivd1_hd U440 ( .A(n86), .Y(n90) );
  ivd1_hd U441 ( .A(n86), .Y(n91) );
  ad2d2_hd U443 ( .A(n130), .B(n438), .Y(n224) );
  ivd1_hd U444 ( .A(n85), .Y(n92) );
  ivd1_hd U445 ( .A(n85), .Y(n93) );
  ivd1_hd U446 ( .A(n85), .Y(n94) );
  ivd4_hd U447 ( .A(n413), .Y(n393) );
  clknd2d1_hd U450 ( .A(n740), .B(n293), .Y(b_e[1]) );
  clknd2d1_hd U453 ( .A(n739), .B(n293), .Y(b_e[2]) );
  clknd2d1_hd U456 ( .A(n738), .B(n293), .Y(b_e[3]) );
  clknd2d1_hd U459 ( .A(n737), .B(n293), .Y(b_e[4]) );
  clknd2d1_hd U462 ( .A(n736), .B(n293), .Y(b_e[5]) );
  clknd2d1_hd U465 ( .A(n735), .B(n293), .Y(b_e[6]) );
  clknd2d1_hd U468 ( .A(n734), .B(n293), .Y(a_e[1]) );
  clknd2d1_hd U471 ( .A(n733), .B(n293), .Y(a_e[2]) );
  clknd2d1_hd U474 ( .A(n732), .B(n293), .Y(a_e[3]) );
  clknd2d1_hd U475 ( .A(n87), .B(n293), .Y(a_e[4]) );
  clknd2d1_hd U476 ( .A(n88), .B(n293), .Y(a_e[5]) );
  clknd2d1_hd U477 ( .A(n89), .B(n293), .Y(a_e[6]) );
  ivd2_hd U482 ( .A(n230), .Y(n222) );
  ivd2_hd U483 ( .A(n333), .Y(n296) );
  clknd2d1_hd U484 ( .A(N543), .B(n391), .Y(n333) );
  clknd2d1_hd U485 ( .A(n315), .B(n316), .Y(n392) );
  nr2d4_hd U486 ( .A(n435), .B(n439), .Y(n232) );
  clknd2d1_hd U487 ( .A(n425), .B(n440), .Y(n435) );
  clknd2d1_hd U489 ( .A(i_AB_STB), .B(o_AB_ACK), .Y(n695) );
  clknd2d1_hd U492 ( .A(n566), .B(n434), .Y(n439) );
  mx2id1_hd U565 ( .D0(n513), .D1(n514), .S(n486), .YN(C2_Z_0) );
  ivd1_hd U568 ( .A(C1_Z_0), .Y(C82_DATA2_0) );
  ivd1_hd U569 ( .A(C1_Z_1), .Y(n188) );
  ao22d1_hd U570 ( .A(C1_Z_1), .B(C82_DATA2_0), .C(C1_Z_0), .D(n188), .Y(
        C82_DATA2_1) );
  nr2d1_hd U571 ( .A(C1_Z_1), .B(C1_Z_0), .Y(n191) );
  ivd1_hd U572 ( .A(n191), .Y(n189) );
  ivd1_hd U573 ( .A(C1_Z_2), .Y(n190) );
  ao22d1_hd U574 ( .A(C1_Z_2), .B(n191), .C(n189), .D(n190), .Y(C82_DATA2_2)
         );
  ivd1_hd U575 ( .A(n194), .Y(n193) );
  ivd1_hd U576 ( .A(C1_Z_3), .Y(n192) );
  ao22d1_hd U577 ( .A(C1_Z_3), .B(n193), .C(n194), .D(n192), .Y(C82_DATA2_3)
         );
  nr2d1_hd U578 ( .A(C1_Z_3), .B(n194), .Y(n197) );
  ivd1_hd U579 ( .A(n197), .Y(n195) );
  ivd1_hd U580 ( .A(C1_Z_4), .Y(n196) );
  ao22d1_hd U581 ( .A(C1_Z_4), .B(n197), .C(n195), .D(n196), .Y(C82_DATA2_4)
         );
  ivd1_hd U582 ( .A(n200), .Y(n199) );
  ivd1_hd U583 ( .A(C1_Z_5), .Y(n198) );
  ao22d1_hd U584 ( .A(C1_Z_5), .B(n199), .C(n200), .D(n198), .Y(C82_DATA2_5)
         );
  nr2d1_hd U585 ( .A(C1_Z_5), .B(n200), .Y(n202) );
  ivd1_hd U586 ( .A(n202), .Y(n201) );
  ivd1_hd U587 ( .A(C1_Z_6), .Y(n203) );
  ao22d1_hd U588 ( .A(C1_Z_6), .B(n202), .C(n201), .D(n203), .Y(C82_DATA2_6)
         );
  ivd1_hd U589 ( .A(n126), .Y(N443) );
  ivd1_hd U590 ( .A(n125), .Y(n205) );
  ao22d1_hd U591 ( .A(n125), .B(N443), .C(n126), .D(n205), .Y(N444) );
  nr2d1_hd U592 ( .A(n125), .B(n126), .Y(n208) );
  ivd1_hd U593 ( .A(n208), .Y(n206) );
  ivd1_hd U594 ( .A(n124), .Y(n207) );
  ao22d1_hd U595 ( .A(n124), .B(n208), .C(n206), .D(n207), .Y(N445) );
  ivd1_hd U596 ( .A(n211), .Y(n210) );
  ivd1_hd U597 ( .A(n123), .Y(n209) );
  ao22d1_hd U598 ( .A(n123), .B(n210), .C(n211), .D(n209), .Y(N446) );
  nr2d1_hd U599 ( .A(n123), .B(n211), .Y(n214) );
  ivd1_hd U600 ( .A(n214), .Y(n212) );
  ivd1_hd U601 ( .A(n122), .Y(n213) );
  ao22d1_hd U602 ( .A(n122), .B(n214), .C(n212), .D(n213), .Y(N447) );
  ivd1_hd U603 ( .A(n217), .Y(n216) );
  ivd1_hd U604 ( .A(n121), .Y(n215) );
  ao22d1_hd U605 ( .A(n121), .B(n216), .C(n217), .D(n215), .Y(N448) );
  nr2d1_hd U606 ( .A(n121), .B(n217), .Y(n219) );
  ivd1_hd U607 ( .A(n219), .Y(n218) );
  ivd1_hd U608 ( .A(n114), .Y(n220) );
  ao22d1_hd U609 ( .A(n114), .B(n219), .C(n218), .D(n220), .Y(N449) );
  scg5d1_hd U610 ( .A(n222), .B(n609), .C(n223), .D(n608), .E(n224), .F(n225), 
        .Y(sticky) );
  scg5d1_hd U611 ( .A(n90), .B(n609), .C(n222), .D(n610), .E(n13), .F(n224), 
        .Y(round_bit) );
  scg4d1_hd U612 ( .A(n93), .B(n14), .C(n222), .D(n611), .E(n22), .F(n224), 
        .G(n91), .H(n610), .Y(guard) );
  oa211d1_hd U613 ( .A(n229), .B(n85), .C(n226), .D(n227), .Y(N667) );
  scg15d1_hd U614 ( .A(n43), .B(n93), .C(n230), .D(n231), .Y(z_m[23]) );
  ao22d1_hd U615 ( .A(n223), .B(n634), .C(n232), .D(N431), .Y(n231) );
  scg15d1_hd U616 ( .A(n222), .B(n634), .C(n233), .D(n234), .Y(z_m[22]) );
  ao22d1_hd U617 ( .A(n232), .B(N430), .C(n91), .D(n633), .Y(n234) );
  ao22d1_hd U618 ( .A(n44), .B(n224), .C(n93), .D(n42), .Y(n233) );
  scg15d1_hd U619 ( .A(n222), .B(n633), .C(n235), .D(n236), .Y(z_m[21]) );
  ao22d1_hd U620 ( .A(n232), .B(N429), .C(n90), .D(n632), .Y(n236) );
  ao22d1_hd U621 ( .A(n94), .B(n41), .C(n224), .D(n43), .Y(n235) );
  scg15d1_hd U622 ( .A(n222), .B(n632), .C(n237), .D(n238), .Y(z_m[20]) );
  ao22d1_hd U623 ( .A(n232), .B(N428), .C(n91), .D(n631), .Y(n238) );
  ao22d1_hd U624 ( .A(n93), .B(n40), .C(n224), .D(n42), .Y(n237) );
  scg15d1_hd U625 ( .A(n222), .B(n631), .C(n239), .D(n240), .Y(z_m[19]) );
  ao22d1_hd U626 ( .A(n232), .B(N427), .C(n90), .D(n630), .Y(n240) );
  ao22d1_hd U627 ( .A(n94), .B(n39), .C(n224), .D(n41), .Y(n239) );
  scg15d1_hd U628 ( .A(n222), .B(n630), .C(n241), .D(n242), .Y(z_m[18]) );
  ao22d1_hd U629 ( .A(n232), .B(N426), .C(n91), .D(n629), .Y(n242) );
  ao22d1_hd U630 ( .A(n93), .B(n38), .C(n224), .D(n40), .Y(n241) );
  scg15d1_hd U631 ( .A(n222), .B(n629), .C(n243), .D(n244), .Y(z_m[17]) );
  ao22d1_hd U632 ( .A(n232), .B(N425), .C(n90), .D(n628), .Y(n244) );
  ao22d1_hd U633 ( .A(n94), .B(n37), .C(n224), .D(n39), .Y(n243) );
  scg15d1_hd U634 ( .A(n222), .B(n628), .C(n245), .D(n246), .Y(z_m[16]) );
  ao22d1_hd U635 ( .A(n232), .B(N424), .C(n91), .D(n627), .Y(n246) );
  ao22d1_hd U636 ( .A(n93), .B(n36), .C(n224), .D(n38), .Y(n245) );
  scg15d1_hd U637 ( .A(n222), .B(n627), .C(n247), .D(n248), .Y(z_m[15]) );
  ao22d1_hd U638 ( .A(n232), .B(N423), .C(n90), .D(n626), .Y(n248) );
  ao22d1_hd U639 ( .A(n94), .B(n35), .C(n224), .D(n37), .Y(n247) );
  scg15d1_hd U640 ( .A(n222), .B(n626), .C(n249), .D(n250), .Y(z_m[14]) );
  ao22d1_hd U641 ( .A(n232), .B(N422), .C(n91), .D(n625), .Y(n250) );
  ao22d1_hd U642 ( .A(n93), .B(n34), .C(n224), .D(n36), .Y(n249) );
  scg15d1_hd U643 ( .A(n222), .B(n625), .C(n251), .D(n252), .Y(z_m[13]) );
  ao22d1_hd U644 ( .A(n232), .B(N421), .C(n90), .D(n624), .Y(n252) );
  ao22d1_hd U645 ( .A(n94), .B(n33), .C(n224), .D(n35), .Y(n251) );
  scg15d1_hd U646 ( .A(n222), .B(n624), .C(n253), .D(n254), .Y(z_m[12]) );
  ao22d1_hd U647 ( .A(n232), .B(N420), .C(n91), .D(n623), .Y(n254) );
  ao22d1_hd U648 ( .A(n93), .B(n32), .C(n224), .D(n34), .Y(n253) );
  scg15d1_hd U649 ( .A(n222), .B(n623), .C(n255), .D(n256), .Y(z_m[11]) );
  ao22d1_hd U650 ( .A(n232), .B(N419), .C(n90), .D(n622), .Y(n256) );
  ao22d1_hd U651 ( .A(n94), .B(n31), .C(n224), .D(n33), .Y(n255) );
  scg15d1_hd U652 ( .A(n222), .B(n622), .C(n257), .D(n258), .Y(z_m[10]) );
  ao22d1_hd U653 ( .A(n232), .B(N418), .C(n91), .D(n621), .Y(n258) );
  ao22d1_hd U654 ( .A(n93), .B(n30), .C(n224), .D(n32), .Y(n257) );
  scg15d1_hd U655 ( .A(n222), .B(n621), .C(n259), .D(n260), .Y(z_m[9]) );
  ao22d1_hd U656 ( .A(n232), .B(N417), .C(n90), .D(n620), .Y(n260) );
  ao22d1_hd U657 ( .A(n94), .B(n29), .C(n224), .D(n31), .Y(n259) );
  scg15d1_hd U658 ( .A(n222), .B(n620), .C(n261), .D(n262), .Y(z_m[8]) );
  ao22d1_hd U659 ( .A(n232), .B(N416), .C(n91), .D(n619), .Y(n262) );
  ao22d1_hd U660 ( .A(n93), .B(n28), .C(n224), .D(n30), .Y(n261) );
  scg15d1_hd U661 ( .A(n222), .B(n619), .C(n263), .D(n264), .Y(z_m[7]) );
  ao22d1_hd U662 ( .A(n232), .B(N415), .C(n90), .D(n618), .Y(n264) );
  ao22d1_hd U663 ( .A(n94), .B(n27), .C(n224), .D(n29), .Y(n263) );
  scg15d1_hd U664 ( .A(n222), .B(n618), .C(n265), .D(n266), .Y(z_m[6]) );
  ao22d1_hd U665 ( .A(n232), .B(N414), .C(n91), .D(n617), .Y(n266) );
  ao22d1_hd U666 ( .A(n93), .B(n26), .C(n224), .D(n28), .Y(n265) );
  scg15d1_hd U667 ( .A(n222), .B(n617), .C(n267), .D(n268), .Y(z_m[5]) );
  ao22d1_hd U668 ( .A(n232), .B(N413), .C(n91), .D(n616), .Y(n268) );
  ao22d1_hd U669 ( .A(n94), .B(n25), .C(n224), .D(n27), .Y(n267) );
  scg15d1_hd U670 ( .A(n222), .B(n616), .C(n269), .D(n270), .Y(z_m[4]) );
  ao22d1_hd U671 ( .A(n232), .B(N412), .C(n90), .D(n615), .Y(n270) );
  ao22d1_hd U672 ( .A(n93), .B(n24), .C(n224), .D(n26), .Y(n269) );
  scg15d1_hd U673 ( .A(n222), .B(n615), .C(n271), .D(n272), .Y(z_m[3]) );
  ao22d1_hd U674 ( .A(n232), .B(N411), .C(n91), .D(n614), .Y(n272) );
  ao22d1_hd U675 ( .A(n94), .B(n563), .C(n224), .D(n25), .Y(n271) );
  scg6d1_hd U676 ( .A(n222), .B(n614), .C(n273), .Y(z_m[2]) );
  scg4d1_hd U677 ( .A(n94), .B(n23), .C(n232), .D(N410), .E(n24), .F(n224), 
        .G(n613), .H(n90), .Y(n273) );
  oa211d1_hd U678 ( .A(n85), .B(n274), .C(n275), .D(n276), .Y(z_m[1]) );
  ao22d1_hd U679 ( .A(n222), .B(n613), .C(n90), .D(n612), .Y(n276) );
  ao22d1_hd U680 ( .A(n224), .B(n563), .C(n232), .D(N409), .Y(n275) );
  scg15d1_hd U681 ( .A(n13), .B(n94), .C(n277), .D(n278), .Y(z_m[0]) );
  ao22d1_hd U682 ( .A(n224), .B(n23), .C(n232), .D(N408), .Y(n278) );
  ao22d1_hd U683 ( .A(n222), .B(n612), .C(n90), .D(n611), .Y(n277) );
  ivd1_hd U684 ( .A(n223), .Y(n226) );
  nd2bd1_hd U685 ( .AN(n283), .B(n224), .Y(n227) );
  ao211d1_hd U686 ( .A(n284), .B(n285), .C(n741), .D(n222), .Y(n282) );
  nr3d1_hd U687 ( .A(n228), .B(n286), .C(n287), .Y(n285) );
  nd4d1_hd U688 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n287) );
  nd4d1_hd U689 ( .A(n40), .B(n39), .C(n38), .D(n37), .Y(n286) );
  oa211d1_hd U690 ( .A(n22), .B(n225), .C(n232), .D(n13), .Y(n228) );
  or2d1_hd U691 ( .A(n14), .B(n15), .Y(n225) );
  nr4d1_hd U692 ( .A(n288), .B(n289), .C(n290), .D(n291), .Y(n284) );
  nd4d1_hd U693 ( .A(n28), .B(n27), .C(n26), .D(n25), .Y(n291) );
  nd4d1_hd U694 ( .A(n22), .B(n24), .C(n563), .D(n23), .Y(n290) );
  nd4d1_hd U695 ( .A(n36), .B(n35), .C(n34), .D(n33), .Y(n289) );
  nd4d1_hd U696 ( .A(n32), .B(n31), .C(n30), .D(n29), .Y(n288) );
  oa211d1_hd U697 ( .A(n292), .B(n293), .C(n294), .D(n295), .Y(n696) );
  oa211d1_hd U698 ( .A(n297), .B(n298), .C(n299), .D(n564), .Y(n294) );
  nd4d1_hd U699 ( .A(n300), .B(n301), .C(n302), .D(n303), .Y(n298) );
  nr4d1_hd U700 ( .A(n29), .B(n28), .C(n27), .D(n26), .Y(n303) );
  nr4d1_hd U701 ( .A(n25), .B(n24), .C(n563), .D(n23), .Y(n302) );
  nr4d1_hd U702 ( .A(n37), .B(n36), .C(n35), .D(n34), .Y(n301) );
  nr4d1_hd U703 ( .A(n33), .B(n32), .C(n31), .D(n30), .Y(n300) );
  nd4d1_hd U704 ( .A(n304), .B(n305), .C(n306), .D(n274), .Y(n297) );
  ivd1_hd U705 ( .A(n22), .Y(n274) );
  nr4d1_hd U706 ( .A(n41), .B(n40), .C(n39), .D(n38), .Y(n306) );
  nr2d1_hd U707 ( .A(n43), .B(n42), .Y(n305) );
  ao211d1_hd U708 ( .A(n661), .B(n307), .C(n308), .D(n309), .Y(n292) );
  ao211d1_hd U709 ( .A(n310), .B(n311), .C(n312), .D(n313), .Y(n308) );
  ivd1_hd U710 ( .A(n314), .Y(n312) );
  oa211d1_hd U711 ( .A(n315), .B(n313), .C(n316), .D(n317), .Y(n307) );
  ao22d1_hd U712 ( .A(N450), .B(n320), .C(C82_DATA2_7), .D(n321), .Y(n318) );
  ao22d1_hd U713 ( .A(N449), .B(n320), .C(C82_DATA2_6), .D(n321), .Y(n322) );
  ao22d1_hd U714 ( .A(N448), .B(n320), .C(C82_DATA2_5), .D(n321), .Y(n323) );
  ao22d1_hd U715 ( .A(N447), .B(n320), .C(C82_DATA2_4), .D(n321), .Y(n324) );
  ao22d1_hd U716 ( .A(N446), .B(n320), .C(C82_DATA2_3), .D(n321), .Y(n325) );
  ao22d1_hd U717 ( .A(N445), .B(n320), .C(C82_DATA2_2), .D(n321), .Y(n326) );
  ao22d1_hd U718 ( .A(N444), .B(n320), .C(C82_DATA2_1), .D(n321), .Y(n327) );
  ao21d1_hd U719 ( .A(N543), .B(n329), .C(n330), .Y(n319) );
  nr2d1_hd U720 ( .A(n331), .B(n332), .Y(n330) );
  ao22d1_hd U721 ( .A(N443), .B(n320), .C(C82_DATA2_0), .D(n321), .Y(n328) );
  nr2d1_hd U722 ( .A(n304), .B(n332), .Y(n320) );
  scg12d1_hd U723 ( .A(n125), .B(n335), .C(n126), .Y(n304) );
  ad4d1_hd U724 ( .A(n111), .B(n336), .C(n337), .D(n338), .Y(n335) );
  scg18d1_hd U725 ( .A(n43), .B(n339), .C(n340), .D(n341), .E(n342), .Y(n705)
         );
  nd4d1_hd U726 ( .A(n310), .B(n541), .C(n314), .D(N543), .Y(n342) );
  ao22d1_hd U727 ( .A(N543), .B(n309), .C(n67), .D(n296), .Y(n341) );
  oa22ad1_hd U728 ( .A(n343), .B(n317), .C(n344), .D(n314), .Y(n309) );
  nr2d1_hd U729 ( .A(n345), .B(n334), .Y(n340) );
  oa21d1_hd U730 ( .A(n346), .B(n334), .C(n347), .Y(n706) );
  ao22d1_hd U731 ( .A(n68), .B(n296), .C(n42), .D(n339), .Y(n347) );
  oa21d1_hd U732 ( .A(n348), .B(n334), .C(n349), .Y(n707) );
  ao22d1_hd U733 ( .A(n69), .B(n296), .C(n41), .D(n339), .Y(n349) );
  oa21d1_hd U734 ( .A(n350), .B(n334), .C(n351), .Y(n708) );
  ao22d1_hd U735 ( .A(n70), .B(n296), .C(n40), .D(n339), .Y(n351) );
  oa21d1_hd U736 ( .A(n352), .B(n334), .C(n353), .Y(n709) );
  ao22d1_hd U737 ( .A(n71), .B(n296), .C(n39), .D(n339), .Y(n353) );
  oa21d1_hd U738 ( .A(n354), .B(n334), .C(n355), .Y(n710) );
  ao22d1_hd U739 ( .A(n72), .B(n296), .C(n38), .D(n339), .Y(n355) );
  oa21d1_hd U740 ( .A(n356), .B(n334), .C(n357), .Y(n711) );
  ao22d1_hd U741 ( .A(n73), .B(n296), .C(n37), .D(n339), .Y(n357) );
  oa21d1_hd U742 ( .A(n358), .B(n334), .C(n359), .Y(n712) );
  ao22d1_hd U743 ( .A(n74), .B(n296), .C(n36), .D(n339), .Y(n359) );
  oa21d1_hd U744 ( .A(n360), .B(n334), .C(n361), .Y(n713) );
  ao22d1_hd U745 ( .A(n75), .B(n296), .C(n35), .D(n339), .Y(n361) );
  oa21d1_hd U746 ( .A(n362), .B(n334), .C(n363), .Y(n714) );
  ao22d1_hd U747 ( .A(n76), .B(n296), .C(n34), .D(n339), .Y(n363) );
  oa21d1_hd U748 ( .A(n364), .B(n334), .C(n365), .Y(n715) );
  ao22d1_hd U749 ( .A(n77), .B(n296), .C(n33), .D(n339), .Y(n365) );
  oa21d1_hd U750 ( .A(n366), .B(n334), .C(n367), .Y(n716) );
  ao22d1_hd U751 ( .A(n78), .B(n296), .C(n32), .D(n339), .Y(n367) );
  oa21d1_hd U752 ( .A(n368), .B(n334), .C(n369), .Y(n717) );
  ao22d1_hd U753 ( .A(n79), .B(n296), .C(n31), .D(n339), .Y(n369) );
  oa21d1_hd U754 ( .A(n370), .B(n334), .C(n371), .Y(n718) );
  ao22d1_hd U755 ( .A(n80), .B(n296), .C(n30), .D(n339), .Y(n371) );
  oa21d1_hd U756 ( .A(n372), .B(n334), .C(n373), .Y(n719) );
  ao22d1_hd U757 ( .A(n81), .B(n296), .C(n29), .D(n339), .Y(n373) );
  oa21d1_hd U758 ( .A(n374), .B(n334), .C(n375), .Y(n720) );
  ao22d1_hd U759 ( .A(n82), .B(n296), .C(n28), .D(n339), .Y(n375) );
  oa21d1_hd U760 ( .A(n376), .B(n334), .C(n377), .Y(n721) );
  ao22d1_hd U761 ( .A(n83), .B(n296), .C(n27), .D(n339), .Y(n377) );
  oa21d1_hd U762 ( .A(n378), .B(n334), .C(n379), .Y(n722) );
  ao22d1_hd U763 ( .A(n108), .B(n296), .C(n26), .D(n339), .Y(n379) );
  oa21d1_hd U764 ( .A(n380), .B(n334), .C(n381), .Y(n723) );
  ao22d1_hd U765 ( .A(n109), .B(n296), .C(n25), .D(n339), .Y(n381) );
  oa21d1_hd U766 ( .A(n382), .B(n334), .C(n383), .Y(n724) );
  ao22d1_hd U767 ( .A(n110), .B(n296), .C(n24), .D(n339), .Y(n383) );
  oa21d1_hd U768 ( .A(n384), .B(n334), .C(n385), .Y(n725) );
  ao22d1_hd U769 ( .A(n115), .B(n296), .C(n563), .D(n339), .Y(n385) );
  oa21d1_hd U770 ( .A(n386), .B(n334), .C(n387), .Y(n726) );
  ao22d1_hd U771 ( .A(n116), .B(n296), .C(n23), .D(n339), .Y(n387) );
  oa21d1_hd U772 ( .A(n388), .B(n334), .C(n389), .Y(n727) );
  ao22d1_hd U773 ( .A(n117), .B(n296), .C(n22), .D(n339), .Y(n389) );
  oa21d1_hd U774 ( .A(n113), .B(n112), .C(n390), .Y(n331) );
  ivd1_hd U775 ( .A(n332), .Y(n299) );
  scg15d1_hd U776 ( .A(n393), .B(n551), .C(n293), .D(n731), .Y(b_e[9]) );
  scg14d1_hd U777 ( .A(n393), .B(n550), .C(n731), .Y(b_e[8]) );
  scg14d1_hd U779 ( .A(n393), .B(C1_DATA2_8), .C(n730), .Y(a_e[8]) );
  oa21d1_hd U780 ( .A(n410), .B(n402), .C(n403), .Y(N573) );
  ivd1_hd U781 ( .A(n411), .Y(n402) );
  ao21d1_hd U782 ( .A(n412), .B(n393), .C(n660), .Y(n403) );
  nr2d1_hd U783 ( .A(n388), .B(n413), .Y(b_m[2]) );
  nr2d1_hd U784 ( .A(n414), .B(n413), .Y(b_m[1]) );
  nr2d1_hd U785 ( .A(n415), .B(n413), .Y(b_m[0]) );
  scg14d1_hd U786 ( .A(n411), .B(n408), .C(n409), .Y(N545) );
  ao21d1_hd U787 ( .A(n416), .B(n417), .C(n660), .Y(n409) );
  ivd1_hd U788 ( .A(n418), .Y(n416) );
  nr2d1_hd U789 ( .A(n419), .B(n413), .Y(a_m[2]) );
  nr2d1_hd U790 ( .A(n420), .B(n413), .Y(a_m[1]) );
  nr2d1_hd U791 ( .A(n421), .B(n413), .Y(a_m[0]) );
  nd2bd1_hd U792 ( .AN(N596), .B(n281), .Y(state[3]) );
  nr2d1_hd U793 ( .A(n224), .B(n232), .Y(n281) );
  nr3d1_hd U794 ( .A(n423), .B(n424), .C(n329), .Y(n422) );
  nd3bd1_hd U795 ( .AN(n741), .B(n280), .C(n413), .Y(state[2]) );
  nr2d1_hd U796 ( .A(n223), .B(n94), .Y(n280) );
  nr2d1_hd U797 ( .A(n425), .B(n426), .Y(n223) );
  nr4d1_hd U799 ( .A(n232), .B(n741), .C(N47), .D(n411), .Y(n429) );
  nr4d1_hd U800 ( .A(n424), .B(n423), .C(n293), .D(n329), .Y(n411) );
  ivd1_hd U801 ( .A(n430), .Y(n329) );
  scg1d1_hd U802 ( .A(n229), .B(n93), .C(N87), .D(n431), .F(n418), .G(n417), 
        .E(N516), .H(n432), .Y(N511) );
  scg13d1_hd U803 ( .A(n232), .B(n433), .C(n426), .Y(n432) );
  scg18d1_hd U804 ( .A(n224), .B(n283), .C(n741), .D(n332), .E(n293), .Y(n433)
         );
  nr2d1_hd U806 ( .A(n434), .B(n435), .Y(n427) );
  oa21d1_hd U807 ( .A(n436), .B(n437), .C(n111), .Y(n283) );
  scg12d1_hd U808 ( .A(n336), .B(n338), .C(n125), .Y(n437) );
  nr2d1_hd U809 ( .A(n412), .B(n413), .Y(n417) );
  nr3d1_hd U810 ( .A(n434), .B(n440), .C(n566), .Y(n438) );
  nr2bd1_hd U811 ( .AN(n441), .B(n442), .Y(n412) );
  ao22d1_hd U812 ( .A(n19), .B(n443), .C(n444), .D(n445), .Y(n442) );
  oa22d1_hd U813 ( .A(n446), .B(n447), .C(n132), .D(n448), .Y(n444) );
  ao22d1_hd U814 ( .A(n128), .B(n449), .C(n450), .D(n451), .Y(n447) );
  scg3d1_hd U815 ( .A(n576), .B(n452), .C(n577), .D(n453), .E(n454), .Y(n451)
         );
  oa211d1_hd U816 ( .A(n578), .B(n455), .C(n456), .D(n457), .Y(n454) );
  oa211d1_hd U817 ( .A(n460), .B(n580), .C(n461), .D(n462), .Y(n459) );
  scg17d1_hd U818 ( .A(n460), .B(n580), .C(n463), .D(n464), .Y(n462) );
  oa211d1_hd U819 ( .A(n581), .B(n465), .C(n466), .D(n66), .Y(n464) );
  ao22d1_hd U820 ( .A(n467), .B(n579), .C(n455), .D(n578), .Y(n458) );
  ivd1_hd U821 ( .A(n468), .Y(n446) );
  ao211d1_hd U822 ( .A(n65), .B(n469), .C(n470), .D(n471), .Y(n418) );
  nd4d1_hd U823 ( .A(n472), .B(n450), .C(n468), .D(n461), .Y(n471) );
  ao22d1_hd U824 ( .A(n584), .B(n476), .C(n586), .D(n477), .Y(n472) );
  nd4d1_hd U825 ( .A(n478), .B(n456), .C(n441), .D(n445), .Y(n470) );
  nr2d1_hd U826 ( .A(n66), .B(n463), .Y(n469) );
  nr2d1_hd U827 ( .A(n587), .B(n481), .Y(n463) );
  ivd1_hd U828 ( .A(n728), .Y(n431) );
  ao22d1_hd U829 ( .A(n337), .B(n482), .C(n390), .D(n483), .Y(n229) );
  ivd1_hd U830 ( .A(n44), .Y(n483) );
  ivd1_hd U831 ( .A(n111), .Y(n390) );
  scg15d1_hd U832 ( .A(n126), .B(n125), .C(n336), .D(n338), .Y(n482) );
  nr2d1_hd U833 ( .A(n123), .B(n124), .Y(n338) );
  nr3d1_hd U834 ( .A(n122), .B(n114), .C(n121), .Y(n336) );
  nr2d1_hd U835 ( .A(n44), .B(n436), .Y(n337) );
  nd3d1_hd U836 ( .A(n440), .B(n484), .C(n605), .Y(n426) );
  nr2d1_hd U837 ( .A(n485), .B(n435), .Y(N47) );
  ivd1_hd U838 ( .A(n129), .Y(n440) );
  nd2bd1_hd U839 ( .AN(n485), .B(n129), .Y(n428) );
  ivd1_hd U840 ( .A(n566), .Y(n484) );
  ivd1_hd U841 ( .A(n605), .Y(n434) );
  ivd1_hd U842 ( .A(n130), .Y(n425) );
  ivd1_hd U843 ( .A(n83), .Y(n487) );
  ivd1_hd U844 ( .A(n61), .Y(n376) );
  ivd1_hd U845 ( .A(n108), .Y(n488) );
  ivd1_hd U846 ( .A(n62), .Y(n378) );
  ivd1_hd U847 ( .A(n109), .Y(n489) );
  ivd1_hd U848 ( .A(n63), .Y(n380) );
  ivd1_hd U849 ( .A(n64), .Y(n382) );
  ivd1_hd U850 ( .A(n115), .Y(n491) );
  ivd1_hd U851 ( .A(n118), .Y(n384) );
  ivd1_hd U852 ( .A(n119), .Y(n386) );
  ivd1_hd U853 ( .A(n120), .Y(n388) );
  ivd1_hd U856 ( .A(n67), .Y(n495) );
  ivd1_hd U857 ( .A(n45), .Y(n345) );
  ivd1_hd U858 ( .A(n68), .Y(n496) );
  ivd1_hd U859 ( .A(n46), .Y(n346) );
  ivd1_hd U860 ( .A(n69), .Y(n497) );
  ivd1_hd U861 ( .A(n47), .Y(n348) );
  ivd1_hd U862 ( .A(n70), .Y(n498) );
  ivd1_hd U863 ( .A(n48), .Y(n350) );
  ivd1_hd U864 ( .A(n71), .Y(n499) );
  ivd1_hd U865 ( .A(n49), .Y(n352) );
  ivd1_hd U866 ( .A(n72), .Y(n500) );
  ivd1_hd U867 ( .A(n50), .Y(n354) );
  ivd1_hd U868 ( .A(n570), .Y(n420) );
  ivd1_hd U869 ( .A(n574), .Y(n414) );
  ivd1_hd U870 ( .A(n73), .Y(n501) );
  ivd1_hd U871 ( .A(n51), .Y(n356) );
  ivd1_hd U872 ( .A(n74), .Y(n502) );
  ivd1_hd U873 ( .A(n52), .Y(n358) );
  ivd1_hd U874 ( .A(n75), .Y(n503) );
  ivd1_hd U875 ( .A(n53), .Y(n360) );
  ivd1_hd U876 ( .A(n76), .Y(n504) );
  ivd1_hd U877 ( .A(n54), .Y(n362) );
  ivd1_hd U878 ( .A(n77), .Y(n505) );
  ivd1_hd U879 ( .A(n55), .Y(n364) );
  ivd1_hd U880 ( .A(n78), .Y(n506) );
  ivd1_hd U881 ( .A(n56), .Y(n366) );
  ivd1_hd U882 ( .A(n79), .Y(n507) );
  ivd1_hd U883 ( .A(n57), .Y(n368) );
  ivd1_hd U884 ( .A(n80), .Y(n508) );
  ivd1_hd U885 ( .A(n58), .Y(n370) );
  ivd1_hd U886 ( .A(n81), .Y(n509) );
  ivd1_hd U887 ( .A(n82), .Y(n510) );
  ivd1_hd U888 ( .A(n60), .Y(n374) );
  ivd1_hd U889 ( .A(n568), .Y(n511) );
  ivd1_hd U890 ( .A(n572), .Y(n512) );
  ivd1_hd U891 ( .A(n567), .Y(n513) );
  ivd1_hd U892 ( .A(n571), .Y(n514) );
  oa22d1_hd U893 ( .A(n515), .B(n449), .C(n474), .D(n516), .Y(C1_Z_7) );
  ivd1_hd U894 ( .A(n128), .Y(n474) );
  oa22d1_hd U895 ( .A(n515), .B(n452), .C(n475), .D(n516), .Y(C1_Z_6) );
  ivd1_hd U896 ( .A(n576), .Y(n475) );
  ivd1_hd U897 ( .A(n582), .Y(n452) );
  oa22d1_hd U898 ( .A(n515), .B(n453), .C(n480), .D(n516), .Y(C1_Z_5) );
  ivd1_hd U899 ( .A(n577), .Y(n480) );
  ivd1_hd U900 ( .A(n583), .Y(n453) );
  oa22d1_hd U901 ( .A(n515), .B(n455), .C(n476), .D(n516), .Y(C1_Z_4) );
  oa22d1_hd U902 ( .A(n515), .B(n467), .C(n473), .D(n516), .Y(C1_Z_3) );
  ivd1_hd U903 ( .A(n579), .Y(n473) );
  oa22d1_hd U904 ( .A(n515), .B(n460), .C(n477), .D(n516), .Y(C1_Z_2) );
  oa22d1_hd U905 ( .A(n515), .B(n465), .C(n481), .D(n516), .Y(C1_Z_1) );
  ivd1_hd U906 ( .A(n581), .Y(n481) );
  oa22d1_hd U907 ( .A(n515), .B(n466), .C(n517), .D(n516), .Y(C1_Z_0) );
  ivd1_hd U908 ( .A(n391), .Y(n516) );
  nr2d1_hd U909 ( .A(n518), .B(n519), .Y(n391) );
  ivd1_hd U910 ( .A(n392), .Y(n515) );
  nd2bd1_hd U911 ( .AN(n519), .B(n424), .Y(n316) );
  nr2d1_hd U912 ( .A(n314), .B(n310), .Y(n430) );
  ivd1_hd U913 ( .A(n317), .Y(n310) );
  nd4d1_hd U914 ( .A(n520), .B(n479), .C(n466), .D(n521), .Y(n317) );
  ivd1_hd U915 ( .A(n65), .Y(n466) );
  ivd1_hd U916 ( .A(n19), .Y(n479) );
  ivd1_hd U917 ( .A(n132), .Y(n520) );
  nr4d1_hd U918 ( .A(n18), .B(n131), .C(n66), .D(n522), .Y(n314) );
  nr2d1_hd U919 ( .A(n408), .B(n344), .Y(n424) );
  nr4d1_hd U920 ( .A(n570), .B(n743), .C(n525), .D(n526), .Y(n524) );
  nd4d1_hd U921 ( .A(n527), .B(n528), .C(n529), .D(n530), .Y(n526) );
  nr4d1_hd U922 ( .A(n70), .B(n80), .C(n69), .D(n81), .Y(n530) );
  nr4d1_hd U923 ( .A(n109), .B(n67), .C(n115), .D(n68), .Y(n529) );
  nr4d1_hd U924 ( .A(n72), .B(n78), .C(n73), .D(n76), .Y(n528) );
  nr4d1_hd U925 ( .A(n83), .B(n79), .C(n108), .D(n74), .Y(n527) );
  nd4d1_hd U926 ( .A(n421), .B(n419), .C(n490), .D(n492), .Y(n525) );
  ivd1_hd U927 ( .A(n116), .Y(n492) );
  ivd1_hd U928 ( .A(n110), .Y(n490) );
  ivd1_hd U929 ( .A(n117), .Y(n419) );
  nr2d1_hd U930 ( .A(n567), .B(n568), .Y(n421) );
  nr4d1_hd U931 ( .A(n71), .B(n77), .C(n75), .D(n82), .Y(n523) );
  or4d1_hd U932 ( .A(n443), .B(n448), .C(n517), .D(n522), .Y(n408) );
  nd4d1_hd U933 ( .A(n128), .B(n531), .C(n477), .D(n476), .Y(n522) );
  ivd1_hd U934 ( .A(n578), .Y(n476) );
  ivd1_hd U935 ( .A(n580), .Y(n477) );
  nr4d1_hd U936 ( .A(n576), .B(n577), .C(n579), .D(n581), .Y(n531) );
  ivd1_hd U937 ( .A(n66), .Y(n517) );
  ivd1_hd U938 ( .A(n131), .Y(n448) );
  ivd1_hd U939 ( .A(n18), .Y(n443) );
  ivd1_hd U940 ( .A(n518), .Y(n423) );
  nr2d1_hd U941 ( .A(n532), .B(n533), .Y(n343) );
  nd4d1_hd U942 ( .A(n415), .B(n534), .C(n535), .D(n372), .Y(n533) );
  ivd1_hd U943 ( .A(n59), .Y(n372) );
  nr4d1_hd U944 ( .A(n574), .B(n607), .C(n63), .D(n45), .Y(n535) );
  nr4d1_hd U945 ( .A(n119), .B(n47), .C(n51), .D(n57), .Y(n534) );
  nr2d1_hd U946 ( .A(n571), .B(n572), .Y(n415) );
  nd4d1_hd U947 ( .A(n536), .B(n537), .C(n538), .D(n539), .Y(n532) );
  nr4d1_hd U948 ( .A(n48), .B(n54), .C(n120), .D(n56), .Y(n539) );
  nr4d1_hd U949 ( .A(n46), .B(n60), .C(n61), .D(n64), .Y(n538) );
  nr4d1_hd U950 ( .A(n118), .B(n52), .C(n62), .D(n49), .Y(n537) );
  nr4d1_hd U951 ( .A(n55), .B(n53), .C(n50), .D(n58), .Y(n536) );
  ivd1_hd U952 ( .A(n401), .Y(n410) );
  nd4d1_hd U953 ( .A(n132), .B(n19), .C(n65), .D(n521), .Y(n401) );
  nr4d1_hd U954 ( .A(n583), .B(n582), .C(n449), .D(n540), .Y(n521) );
  nd4d1_hd U955 ( .A(n467), .B(n465), .C(n455), .D(n460), .Y(n540) );
  ivd1_hd U956 ( .A(n586), .Y(n460) );
  ivd1_hd U957 ( .A(n584), .Y(n455) );
  ivd1_hd U958 ( .A(n587), .Y(n465) );
  ivd1_hd U959 ( .A(n585), .Y(n467) );
  ivd1_hd U960 ( .A(n127), .Y(n449) );
  ivd1_hd U1 ( .A(i_RST), .Y(n1) );
  ivd1_hd U2 ( .A(i_RST), .Y(n2) );
  ivd1_hd U3 ( .A(i_RST), .Y(n3) );
  ivd1_hd U4 ( .A(i_RST), .Y(n4) );
  ivd1_hd U5 ( .A(i_RST), .Y(n5) );
  ivd1_hd U6 ( .A(i_RST), .Y(n12) );
  ivd6_hd U11 ( .A(n6) );
  ivd6_hd U12 ( .A(n11) );
  ivd6_hd U13 ( .A(n10) );
  ivd6_hd U14 ( .A(n7) );
  ivd6_hd U15 ( .A(n8) );
  ivd6_hd U16 ( .A(n9) );
  fds2eqd1_hd clk_r_REG136_S4 ( .CRN(n2), .D(state[2]), .E(N511), .CK(i_CLK), 
        .Q(n130) );
  fds2eqd1_hd clk_r_REG135_S4 ( .CRN(n12), .D(state[0]), .E(N511), .CK(i_CLK), 
        .Q(n605) );
  fds2eqd1_hd clk_r_REG125_S3 ( .CRN(n3), .D(state[3]), .E(N511), .CK(i_CLK), 
        .Q(n566) );
  fd1eqd1_hd clk_r_REG77_S13 ( .D(sticky), .E(N668), .CK(n754), .Q(n15) );
  fd1eqd1_hd clk_r_REG74_S10 ( .D(z_m[0]), .E(N664), .CK(n758), .Q(n22) );
  fd1eqd1_hd clk_r_REG145_S8 ( .D(b_m[0]), .E(n573), .CK(n753), .Q(n571) );
  fd1eqd1_hd clk_r_REG128_S4 ( .D(z_e[2]), .E(N629), .CK(n758), .Q(n124) );
  fd1eqd1_hd clk_r_REG127_S4 ( .D(z_e[1]), .E(N629), .CK(n758), .Q(n125) );
  fd1eqd1_hd clk_r_REG126_S4 ( .D(z_e[0]), .E(N629), .CK(n758), .Q(n126) );
  fd1eqd1_hd clk_r_REG151_S8 ( .D(a_m[0]), .E(n569), .CK(n752), .Q(n567) );
  fd1eqd1_hd clk_r_REG129_S4 ( .D(z_e[3]), .E(N629), .CK(n758), .Q(n123) );
  fd1eqd1_hd clk_r_REG130_S4 ( .D(z_e[4]), .E(N629), .CK(n758), .Q(n122) );
  fd1eqd1_hd clk_r_REG180_S5 ( .D(a_e[6]), .E(N574), .CK(n758), .Q(n576) );
  fd1eqd1_hd clk_r_REG179_S5 ( .D(a_e[5]), .E(N574), .CK(n758), .Q(n577) );
  fd1eqd1_hd clk_r_REG178_S5 ( .D(a_e[4]), .E(N574), .CK(n758), .Q(n578) );
  fd1eqd1_hd clk_r_REG177_S5 ( .D(a_e[3]), .E(N574), .CK(n758), .Q(n579) );
  fd1eqd1_hd clk_r_REG176_S5 ( .D(a_e[2]), .E(N574), .CK(n758), .Q(n580) );
  fd1eqd1_hd clk_r_REG175_S5 ( .D(a_e[1]), .E(N574), .CK(n758), .Q(n581) );
  fd1eqd1_hd clk_r_REG174_S5 ( .D(a_e[0]), .E(N574), .CK(n758), .Q(n66) );
  fd1eqd1_hd clk_r_REG138_S2 ( .D(a_e[8]), .E(N574), .CK(n758), .Q(n131) );
  fd1eqd1_hd clk_r_REG137_S5 ( .D(a_e[7]), .E(N574), .CK(n758), .Q(n128) );
  fd1eqd1_hd clk_r_REG187_S5 ( .D(b_e[6]), .E(N585), .CK(n758), .Q(n582) );
  fd1eqd1_hd clk_r_REG186_S5 ( .D(b_e[5]), .E(N585), .CK(n758), .Q(n583) );
  fd1eqd1_hd clk_r_REG181_S5 ( .D(b_e[0]), .E(N585), .CK(n758), .Q(n65) );
  fd1eqd1_hd clk_r_REG141_S6 ( .D(b_e[9]), .E(N585), .CK(n758), .Q(n19) );
  fd1eqd1_hd clk_r_REG140_S6 ( .D(b_e[8]), .E(N585), .CK(n758), .Q(n132) );
  fd1eqd1_hd clk_r_REG139_S5 ( .D(b_e[7]), .E(N585), .CK(n758), .Q(n127) );
  fd1eqd1_hd clk_r_REG131_S4 ( .D(z_e[5]), .E(N629), .CK(n758), .Q(n121) );
  fd1eqd1_hd clk_r_REG132_S4 ( .D(z_e[6]), .E(N629), .CK(n758), .Q(n114) );
  fd1eqd1_hd clk_r_REG133_S4 ( .D(z_e[7]), .E(N629), .CK(n758), .Q(n113) );
  fd1eqd1_hd clk_r_REG134_S4 ( .D(z_e[8]), .E(N629), .CK(n758), .Q(n112) );
  fd1eqd1_hd clk_r_REG124_S3 ( .D(z_e[9]), .E(N629), .CK(i_CLK), .Q(n111) );
  fd1eqd1_hd clk_r_REG19_S20 ( .D(z_m[23]), .E(N664), .CK(n758), .Q(n44) );
  oa21d2_hd U7 ( .A(n514), .B(n486), .C(n179), .Y(C3_Z_0) );
  or2d8_hd U9 ( .A(N220), .B(n185), .Y(n729) );
  mx2id1_hd U10 ( .D0(n419), .D1(n388), .S(n486), .YN(C2_Z_3) );
  clknd2d1_hd U17 ( .A(n566), .B(n427), .Y(n332) );
  nr2d4_hd U20 ( .A(n177), .B(n182), .Y(n541) );
  clknd2d1_hd U22 ( .A(n660), .B(C1_DATA1_8), .Y(n730) );
  clknd2d1_hd U23 ( .A(n660), .B(n560), .Y(n731) );
  ao22d1_hd U24 ( .A(n393), .B(C1_DATA2_3), .C(n660), .D(C1_DATA1_3), .Y(n732)
         );
  ao22d1_hd U25 ( .A(n393), .B(C1_DATA2_2), .C(n660), .D(C1_DATA1_2), .Y(n733)
         );
  ao22d1_hd U32 ( .A(n393), .B(C1_DATA2_1), .C(n660), .D(C1_DATA1_1), .Y(n734)
         );
  ao22d1_hd U33 ( .A(n393), .B(n548), .C(n660), .D(n558), .Y(n735) );
  ao22d1_hd U34 ( .A(n393), .B(n547), .C(n660), .D(n557), .Y(n736) );
  ao22d1_hd U35 ( .A(n393), .B(n546), .C(n660), .D(n556), .Y(n737) );
  ao22d1_hd U36 ( .A(n393), .B(n545), .C(n660), .D(n555), .Y(n738) );
  ao22d1_hd U37 ( .A(n393), .B(n544), .C(n660), .D(n554), .Y(n739) );
  ao22d1_hd U38 ( .A(n393), .B(n543), .C(n660), .D(n553), .Y(n740) );
  ivd4_hd U39 ( .A(n84), .Y(n660) );
  fd1qd1_hd clk_r_REG0_S1 ( .D(i_A[31]), .CK(n748), .Q(n686) );
  fd1qd1_hd clk_r_REG222_S1 ( .D(i_A[22]), .CK(n748), .Q(n685) );
  fd1qd1_hd clk_r_REG223_S1 ( .D(i_A[21]), .CK(n748), .Q(n684) );
  fd1qd1_hd clk_r_REG224_S1 ( .D(i_A[20]), .CK(n748), .Q(n683) );
  fd1qd1_hd clk_r_REG225_S1 ( .D(i_A[19]), .CK(n748), .Q(n682) );
  fd1qd1_hd clk_r_REG226_S1 ( .D(i_A[18]), .CK(n748), .Q(n681) );
  fd1qd1_hd clk_r_REG227_S1 ( .D(i_A[17]), .CK(n748), .Q(n680) );
  fd1qd1_hd clk_r_REG228_S1 ( .D(i_A[16]), .CK(n748), .Q(n679) );
  fd1qd1_hd clk_r_REG229_S1 ( .D(i_A[15]), .CK(n748), .Q(n678) );
  fd1qd1_hd clk_r_REG230_S1 ( .D(i_A[14]), .CK(n748), .Q(n677) );
  fd1qd1_hd clk_r_REG231_S1 ( .D(i_A[13]), .CK(n748), .Q(n676) );
  fd1qd1_hd clk_r_REG232_S1 ( .D(i_A[12]), .CK(n748), .Q(n675) );
  fd1qd1_hd clk_r_REG233_S1 ( .D(i_A[11]), .CK(n748), .Q(n674) );
  fd1qd1_hd clk_r_REG234_S1 ( .D(i_A[10]), .CK(n748), .Q(n673) );
  fd1qd1_hd clk_r_REG235_S1 ( .D(i_A[9]), .CK(n748), .Q(n672) );
  fd1qd1_hd clk_r_REG236_S1 ( .D(i_A[8]), .CK(n748), .Q(n671) );
  fd1qd1_hd clk_r_REG237_S1 ( .D(i_A[7]), .CK(n748), .Q(n670) );
  fd1qd1_hd clk_r_REG238_S1 ( .D(i_A[6]), .CK(n748), .Q(n669) );
  fd1qd1_hd clk_r_REG239_S1 ( .D(i_A[5]), .CK(n748), .Q(n668) );
  fd1qd1_hd clk_r_REG240_S1 ( .D(i_A[4]), .CK(n748), .Q(n667) );
  fd1qd1_hd clk_r_REG241_S1 ( .D(i_A[3]), .CK(n748), .Q(n666) );
  fd1qd1_hd clk_r_REG242_S1 ( .D(i_A[2]), .CK(n748), .Q(n665) );
  fd1qd1_hd clk_r_REG243_S1 ( .D(i_A[1]), .CK(n748), .Q(n664) );
  fd1qd1_hd clk_r_REG244_S1 ( .D(i_A[0]), .CK(n748), .Q(n663) );
  fd1qd1_hd clk_r_REG245_S1 ( .D(i_B[31]), .CK(n748), .Q(n662) );
  fd1qd1_hd clk_r_REG255_S1 ( .D(i_B[22]), .CK(n748), .Q(n659) );
  fd1qd1_hd clk_r_REG256_S1 ( .D(i_B[21]), .CK(n748), .Q(n658) );
  fd1qd1_hd clk_r_REG257_S1 ( .D(i_B[20]), .CK(n748), .Q(n657) );
  fd1qd1_hd clk_r_REG258_S1 ( .D(i_B[19]), .CK(n748), .Q(n656) );
  fd1qd1_hd clk_r_REG259_S1 ( .D(i_B[18]), .CK(n748), .Q(n655) );
  fd1qd1_hd clk_r_REG260_S1 ( .D(i_B[17]), .CK(n748), .Q(n654) );
  fd1qd1_hd clk_r_REG261_S1 ( .D(i_B[16]), .CK(n748), .Q(n653) );
  fd1qd1_hd clk_r_REG262_S1 ( .D(i_B[15]), .CK(n748), .Q(n652) );
  fd1qd1_hd clk_r_REG263_S1 ( .D(i_B[14]), .CK(n748), .Q(n651) );
  fd1qd1_hd clk_r_REG264_S1 ( .D(i_B[13]), .CK(n748), .Q(n650) );
  fd1qd1_hd clk_r_REG265_S1 ( .D(i_B[12]), .CK(n748), .Q(n649) );
  fd1qd1_hd clk_r_REG266_S1 ( .D(i_B[11]), .CK(n748), .Q(n648) );
  fd1qd1_hd clk_r_REG267_S1 ( .D(i_B[10]), .CK(n748), .Q(n647) );
  fd1qd1_hd clk_r_REG268_S1 ( .D(i_B[9]), .CK(n748), .Q(n646) );
  fd1qd1_hd clk_r_REG269_S1 ( .D(i_B[8]), .CK(n748), .Q(n645) );
  fd1qd1_hd clk_r_REG270_S1 ( .D(i_B[7]), .CK(n748), .Q(n644) );
  fd1qd1_hd clk_r_REG271_S1 ( .D(i_B[6]), .CK(n748), .Q(n643) );
  fd1qd1_hd clk_r_REG272_S1 ( .D(i_B[5]), .CK(n748), .Q(n642) );
  fd1qd1_hd clk_r_REG273_S1 ( .D(i_B[4]), .CK(n748), .Q(n641) );
  fd1qd1_hd clk_r_REG274_S1 ( .D(i_B[3]), .CK(n748), .Q(n640) );
  fd1qd1_hd clk_r_REG275_S1 ( .D(i_B[2]), .CK(n748), .Q(n639) );
  fd1qd1_hd clk_r_REG276_S1 ( .D(i_B[1]), .CK(n748), .Q(n638) );
  fd1qd1_hd clk_r_REG277_S1 ( .D(i_B[0]), .CK(n748), .Q(n637) );
  fd1qd1_hd clk_r_REG22_S21 ( .D(n697), .CK(n749), .Q(n589) );
  fd1qd1_hd clk_r_REG24_S21 ( .D(n698), .CK(n749), .Q(n591) );
  fd1qd1_hd clk_r_REG26_S21 ( .D(n699), .CK(n749), .Q(n593) );
  fd1qd1_hd clk_r_REG28_S21 ( .D(n700), .CK(n749), .Q(n595) );
  fd1qd1_hd clk_r_REG30_S21 ( .D(n701), .CK(n749), .Q(n597) );
  fd1qd1_hd clk_r_REG32_S21 ( .D(n702), .CK(n749), .Q(n599) );
  fd1qd1_hd clk_r_REG34_S21 ( .D(n703), .CK(n749), .Q(n601) );
  fd1qd1_hd clk_r_REG36_S21 ( .D(n704), .CK(n749), .Q(n603) );
  fd1qd1_hd clk_r_REG38_S20 ( .D(n705), .CK(n749), .Q(n17) );
  fd1qd1_hd clk_r_REG40_S19 ( .D(n706), .CK(n749), .Q(n562) );
  fd1qd1_hd clk_r_REG42_S18 ( .D(n707), .CK(n749), .Q(n187) );
  fd1qd1_hd clk_r_REG44_S17 ( .D(n708), .CK(n749), .Q(n172) );
  fd1qd1_hd clk_r_REG46_S16 ( .D(n709), .CK(n749), .Q(n170) );
  fd1qd1_hd clk_r_REG48_S15 ( .D(n710), .CK(n749), .Q(n168) );
  fd1qd1_hd clk_r_REG50_S14 ( .D(n711), .CK(n749), .Q(n166) );
  fd1qd1_hd clk_r_REG52_S13 ( .D(n712), .CK(n749), .Q(n164) );
  fd1qd1_hd clk_r_REG54_S12 ( .D(n713), .CK(n749), .Q(n162) );
  fd1qd1_hd clk_r_REG56_S11 ( .D(n714), .CK(n749), .Q(n160) );
  fd1qd1_hd clk_r_REG58_S10 ( .D(n715), .CK(n749), .Q(n158) );
  fd1qd1_hd clk_r_REG60_S9 ( .D(n716), .CK(n749), .Q(n156) );
  fd1qd1_hd clk_r_REG62_S8 ( .D(n717), .CK(n749), .Q(n154) );
  fd1qd1_hd clk_r_REG64_S7 ( .D(n718), .CK(n749), .Q(n152) );
  fd1qd1_hd clk_r_REG66_S6 ( .D(n719), .CK(n749), .Q(n150) );
  fd1qd1_hd clk_r_REG78_S11 ( .D(n727), .CK(n749), .Q(n134) );
  fd1qd1_hd clk_r_REG80_S10 ( .D(n726), .CK(n749), .Q(n136) );
  fd1qd1_hd clk_r_REG82_S9 ( .D(n725), .CK(n749), .Q(n138) );
  fd1qd1_hd clk_r_REG84_S8 ( .D(n724), .CK(n749), .Q(n140) );
  fd1qd1_hd clk_r_REG86_S7 ( .D(n723), .CK(n749), .Q(n142) );
  fd1qd1_hd clk_r_REG88_S6 ( .D(n722), .CK(n749), .Q(n144) );
  fd1qd1_hd clk_r_REG90_S5 ( .D(n721), .CK(n749), .Q(n146) );
  fd1qd1_hd clk_r_REG92_S5 ( .D(n720), .CK(n749), .Q(n148) );
  fd1qd1_hd clk_r_REG20_S21 ( .D(n696), .CK(n749), .Q(n21) );
  fd1qd1_hd clk_r_REG21_S22 ( .D(n21), .CK(n750), .Q(o_Z[31]) );
  fd1qd1_hd clk_r_REG23_S22 ( .D(n589), .CK(n750), .Q(o_Z[30]) );
  fd1qd1_hd clk_r_REG25_S22 ( .D(n591), .CK(n750), .Q(o_Z[29]) );
  fd1qd1_hd clk_r_REG27_S22 ( .D(n593), .CK(n750), .Q(o_Z[28]) );
  fd1qd1_hd clk_r_REG29_S22 ( .D(n595), .CK(n750), .Q(o_Z[27]) );
  fd1qd1_hd clk_r_REG31_S22 ( .D(n597), .CK(n750), .Q(o_Z[26]) );
  fd1qd1_hd clk_r_REG33_S22 ( .D(n599), .CK(n750), .Q(o_Z[25]) );
  fd1qd1_hd clk_r_REG35_S22 ( .D(n601), .CK(n750), .Q(o_Z[24]) );
  fd1qd1_hd clk_r_REG37_S22 ( .D(n603), .CK(n750), .Q(o_Z[23]) );
  fd1qd1_hd clk_r_REG39_S21 ( .D(n17), .CK(n750), .Q(o_Z[22]) );
  fd1qd1_hd clk_r_REG41_S20 ( .D(n562), .CK(n750), .Q(o_Z[21]) );
  fd1qd1_hd clk_r_REG43_S19 ( .D(n187), .CK(n750), .Q(o_Z[20]) );
  fd1qd1_hd clk_r_REG45_S18 ( .D(n172), .CK(n750), .Q(o_Z[19]) );
  fd1qd1_hd clk_r_REG47_S17 ( .D(n170), .CK(n750), .Q(o_Z[18]) );
  fd1qd1_hd clk_r_REG49_S16 ( .D(n168), .CK(n750), .Q(o_Z[17]) );
  fd1qd1_hd clk_r_REG51_S15 ( .D(n166), .CK(n750), .Q(o_Z[16]) );
  fd1qd1_hd clk_r_REG53_S14 ( .D(n164), .CK(n750), .Q(o_Z[15]) );
  fd1qd1_hd clk_r_REG55_S13 ( .D(n162), .CK(n750), .Q(o_Z[14]) );
  fd1qd1_hd clk_r_REG57_S12 ( .D(n160), .CK(n750), .Q(o_Z[13]) );
  fd1qd1_hd clk_r_REG59_S11 ( .D(n158), .CK(n750), .Q(o_Z[12]) );
  fd1qd1_hd clk_r_REG61_S10 ( .D(n156), .CK(n750), .Q(o_Z[11]) );
  fd1qd1_hd clk_r_REG63_S9 ( .D(n154), .CK(n750), .Q(o_Z[10]) );
  fd1qd1_hd clk_r_REG65_S8 ( .D(n152), .CK(n750), .Q(o_Z[9]) );
  fd1qd1_hd clk_r_REG67_S7 ( .D(n150), .CK(n750), .Q(o_Z[8]) );
  fd1qd1_hd clk_r_REG79_S12 ( .D(n134), .CK(n750), .Q(o_Z[0]) );
  fd1qd1_hd clk_r_REG81_S11 ( .D(n136), .CK(n750), .Q(o_Z[1]) );
  fd1qd1_hd clk_r_REG83_S10 ( .D(n138), .CK(n750), .Q(o_Z[2]) );
  fd1qd1_hd clk_r_REG85_S9 ( .D(n140), .CK(n750), .Q(o_Z[3]) );
  fd1qd1_hd clk_r_REG87_S8 ( .D(n142), .CK(n750), .Q(o_Z[4]) );
  fd1qd1_hd clk_r_REG89_S7 ( .D(n144), .CK(n750), .Q(o_Z[5]) );
  fd1qd1_hd clk_r_REG91_S6 ( .D(n146), .CK(n750), .Q(o_Z[6]) );
  fd1qd1_hd clk_r_REG93_S6 ( .D(n148), .CK(n750), .Q(o_Z[7]) );
  fd1qd1_hd clk_r_REG110_S3 ( .D(sum[27]), .CK(n751), .Q(n636) );
  fd1qd1_hd clk_r_REG109_S3 ( .D(sum[26]), .CK(n751), .Q(n634) );
  fd1qd1_hd clk_r_REG108_S3 ( .D(sum[25]), .CK(n751), .Q(n633) );
  fd1qd1_hd clk_r_REG107_S3 ( .D(sum[24]), .CK(n751), .Q(n632) );
  fd1qd1_hd clk_r_REG106_S3 ( .D(sum[23]), .CK(n751), .Q(n631) );
  fd1qd1_hd clk_r_REG105_S3 ( .D(sum[22]), .CK(n751), .Q(n630) );
  fd1qd1_hd clk_r_REG104_S3 ( .D(sum[21]), .CK(n751), .Q(n629) );
  fd1qd1_hd clk_r_REG103_S3 ( .D(sum[20]), .CK(n751), .Q(n628) );
  fd1qd1_hd clk_r_REG102_S3 ( .D(sum[19]), .CK(n751), .Q(n627) );
  fd1qd1_hd clk_r_REG101_S3 ( .D(sum[18]), .CK(n751), .Q(n626) );
  fd1qd1_hd clk_r_REG100_S3 ( .D(sum[17]), .CK(n751), .Q(n625) );
  fd1qd1_hd clk_r_REG99_S3 ( .D(sum[16]), .CK(n751), .Q(n624) );
  fd1qd1_hd clk_r_REG98_S3 ( .D(sum[15]), .CK(n751), .Q(n623) );
  fd1qd1_hd clk_r_REG97_S3 ( .D(sum[14]), .CK(n751), .Q(n622) );
  fd1qd1_hd clk_r_REG96_S3 ( .D(sum[13]), .CK(n751), .Q(n621) );
  fd1qd1_hd clk_r_REG95_S3 ( .D(sum[12]), .CK(n751), .Q(n620) );
  fd1qd1_hd clk_r_REG94_S3 ( .D(sum[11]), .CK(n751), .Q(n619) );
  fd1qd1_hd clk_r_REG2_S3 ( .D(sum[10]), .CK(n751), .Q(n618) );
  fd1qd1_hd clk_r_REG111_S3 ( .D(sum[9]), .CK(n751), .Q(n617) );
  fd1qd1_hd clk_r_REG112_S3 ( .D(sum[8]), .CK(n751), .Q(n616) );
  fd1qd1_hd clk_r_REG113_S3 ( .D(sum[7]), .CK(n751), .Q(n615) );
  fd1qd1_hd clk_r_REG116_S3 ( .D(sum[6]), .CK(n751), .Q(n614) );
  fd1qd1_hd clk_r_REG115_S3 ( .D(sum[5]), .CK(n751), .Q(n613) );
  fd1qd1_hd clk_r_REG118_S3 ( .D(sum[4]), .CK(n751), .Q(n612) );
  fd1qd1_hd clk_r_REG117_S3 ( .D(sum[3]), .CK(n751), .Q(n611) );
  fd1qd1_hd clk_r_REG121_S3 ( .D(sum[2]), .CK(n751), .Q(n610) );
  fd1qd1_hd clk_r_REG120_S3 ( .D(sum[1]), .CK(n751), .Q(n609) );
  fd1qd1_hd clk_r_REG119_S3 ( .D(sum[0]), .CK(n751), .Q(n608) );
  fd1qd1_hd clk_r_REG114_S3 ( .D(z_s), .CK(n751), .Q(n564) );
  fd1qd1_hd clk_r_REG123_S2 ( .D(n795), .CK(n752), .Q(n18) );
  fd1qd1_hd clk_r_REG148_S5 ( .D(a_m[3]), .CK(n752), .Q(n117) );
  fd1qd1_hd clk_r_REG149_S6 ( .D(a_m[2]), .CK(n752), .Q(n570) );
  fd1qd1_hd clk_r_REG150_S7 ( .D(a_m[1]), .CK(n752), .Q(n568) );
  fd1qd1_hd clk_r_REG152_S5 ( .D(a_m[4]), .CK(n752), .Q(n116) );
  fd1qd1_hd clk_r_REG153_S5 ( .D(a_m[5]), .CK(n752), .Q(n115) );
  fd1qd1_hd clk_r_REG154_S5 ( .D(a_m[6]), .CK(n752), .Q(n110) );
  fd1qd1_hd clk_r_REG155_S5 ( .D(a_m[7]), .CK(n752), .Q(n109) );
  fd1qd1_hd clk_r_REG156_S5 ( .D(a_m[8]), .CK(n752), .Q(n108) );
  fd1qd1_hd clk_r_REG157_S5 ( .D(a_m[9]), .CK(n752), .Q(n83) );
  fd1qd1_hd clk_r_REG158_S5 ( .D(a_m[10]), .CK(n752), .Q(n82) );
  fd1qd1_hd clk_r_REG159_S5 ( .D(a_m[11]), .CK(n752), .Q(n81) );
  fd1qd1_hd clk_r_REG160_S5 ( .D(a_m[12]), .CK(n752), .Q(n80) );
  fd1qd1_hd clk_r_REG161_S5 ( .D(a_m[13]), .CK(n752), .Q(n79) );
  fd1qd1_hd clk_r_REG162_S5 ( .D(a_m[14]), .CK(n752), .Q(n78) );
  fd1qd1_hd clk_r_REG163_S5 ( .D(a_m[15]), .CK(n752), .Q(n77) );
  fd1qd1_hd clk_r_REG164_S5 ( .D(a_m[16]), .CK(n752), .Q(n76) );
  fd1qd1_hd clk_r_REG165_S5 ( .D(a_m[17]), .CK(n752), .Q(n75) );
  fd1qd1_hd clk_r_REG166_S5 ( .D(a_m[18]), .CK(n752), .Q(n74) );
  fd1qd1_hd clk_r_REG167_S5 ( .D(a_m[19]), .CK(n752), .Q(n73) );
  fd1qd1_hd clk_r_REG168_S5 ( .D(a_m[20]), .CK(n752), .Q(n72) );
  fd1qd1_hd clk_r_REG169_S5 ( .D(a_m[21]), .CK(n752), .Q(n71) );
  fd1qd1_hd clk_r_REG170_S5 ( .D(a_m[22]), .CK(n752), .Q(n70) );
  fd1qd1_hd clk_r_REG172_S5 ( .D(a_m[24]), .CK(n752), .Q(n68) );
  fd1qd1_hd clk_r_REG173_S5 ( .D(a_m[25]), .CK(n752), .Q(n67) );
  fd1qd1_hd clk_r_REG142_S5 ( .D(b_m[3]), .CK(n753), .Q(n120) );
  fd1qd1_hd clk_r_REG143_S6 ( .D(b_m[2]), .CK(n753), .Q(n574) );
  fd1qd1_hd clk_r_REG144_S7 ( .D(b_m[1]), .CK(n753), .Q(n572) );
  fd1qd1_hd clk_r_REG146_S5 ( .D(b_m[4]), .CK(n753), .Q(n119) );
  fd1qd1_hd clk_r_REG147_S5 ( .D(b_m[5]), .CK(n753), .Q(n118) );
  fd1qd1_hd clk_r_REG188_S5 ( .D(b_m[6]), .CK(n753), .Q(n64) );
  fd1qd1_hd clk_r_REG189_S5 ( .D(b_m[7]), .CK(n753), .Q(n63) );
  fd1qd1_hd clk_r_REG190_S5 ( .D(b_m[8]), .CK(n753), .Q(n62) );
  fd1qd1_hd clk_r_REG191_S5 ( .D(b_m[9]), .CK(n753), .Q(n61) );
  fd1qd1_hd clk_r_REG192_S5 ( .D(b_m[10]), .CK(n753), .Q(n60) );
  fd1qd1_hd clk_r_REG193_S5 ( .D(b_m[11]), .CK(n753), .Q(n59) );
  fd1qd1_hd clk_r_REG194_S5 ( .D(b_m[12]), .CK(n753), .Q(n58) );
  fd1qd1_hd clk_r_REG195_S5 ( .D(b_m[13]), .CK(n753), .Q(n57) );
  fd1qd1_hd clk_r_REG196_S5 ( .D(b_m[14]), .CK(n753), .Q(n56) );
  fd1qd1_hd clk_r_REG197_S5 ( .D(b_m[15]), .CK(n753), .Q(n55) );
  fd1qd1_hd clk_r_REG198_S5 ( .D(b_m[16]), .CK(n753), .Q(n54) );
  fd1qd1_hd clk_r_REG199_S5 ( .D(b_m[17]), .CK(n753), .Q(n53) );
  fd1qd1_hd clk_r_REG200_S5 ( .D(b_m[18]), .CK(n753), .Q(n52) );
  fd1qd1_hd clk_r_REG201_S5 ( .D(b_m[19]), .CK(n753), .Q(n51) );
  fd1qd1_hd clk_r_REG202_S5 ( .D(b_m[20]), .CK(n753), .Q(n50) );
  fd1qd1_hd clk_r_REG203_S5 ( .D(b_m[21]), .CK(n753), .Q(n49) );
  fd1qd1_hd clk_r_REG204_S5 ( .D(b_m[22]), .CK(n753), .Q(n48) );
  fd1qd1_hd clk_r_REG205_S5 ( .D(b_m[23]), .CK(n753), .Q(n47) );
  fd1qd1_hd clk_r_REG206_S5 ( .D(b_m[24]), .CK(n753), .Q(n46) );
  fd1qd1_hd clk_r_REG207_S5 ( .D(b_m[25]), .CK(n753), .Q(n45) );
  fd1qd1_hd clk_r_REG18_S19 ( .D(z_m[22]), .CK(n754), .Q(n43) );
  fd1qd1_hd clk_r_REG17_S18 ( .D(z_m[21]), .CK(n754), .Q(n42) );
  fd1qd1_hd clk_r_REG16_S17 ( .D(z_m[20]), .CK(n754), .Q(n41) );
  fd1qd1_hd clk_r_REG15_S16 ( .D(z_m[19]), .CK(n754), .Q(n40) );
  fd1qd1_hd clk_r_REG14_S15 ( .D(z_m[18]), .CK(n754), .Q(n39) );
  fd1qd1_hd clk_r_REG13_S14 ( .D(z_m[17]), .CK(n754), .Q(n38) );
  fd1qd1_hd clk_r_REG12_S13 ( .D(z_m[16]), .CK(n754), .Q(n37) );
  fd1qd1_hd clk_r_REG11_S12 ( .D(z_m[15]), .CK(n754), .Q(n36) );
  fd1qd1_hd clk_r_REG10_S11 ( .D(z_m[14]), .CK(n754), .Q(n35) );
  fd1qd1_hd clk_r_REG9_S10 ( .D(z_m[13]), .CK(n754), .Q(n34) );
  fd1qd1_hd clk_r_REG8_S9 ( .D(z_m[12]), .CK(n754), .Q(n33) );
  fd1qd1_hd clk_r_REG7_S8 ( .D(z_m[11]), .CK(n754), .Q(n32) );
  fd1qd1_hd clk_r_REG72_S8 ( .D(z_m[2]), .CK(n754), .Q(n563) );
  fd1qd1_hd clk_r_REG73_S9 ( .D(z_m[1]), .CK(n754), .Q(n23) );
  fd1qd1_hd clk_r_REG3_S4 ( .D(z_m[7]), .CK(n754), .Q(n28) );
  fd1qd1_hd clk_r_REG5_S6 ( .D(z_m[9]), .CK(n754), .Q(n30) );
  fd1qd1_hd clk_r_REG70_S6 ( .D(z_m[4]), .CK(n754), .Q(n25) );
  fd1qd1_hd clk_r_REG4_S5 ( .D(z_m[8]), .CK(n754), .Q(n29) );
  fd1qd1_hd clk_r_REG6_S7 ( .D(z_m[10]), .CK(n754), .Q(n31) );
  fd1qd1_hd clk_r_REG68_S4 ( .D(z_m[6]), .CK(n754), .Q(n27) );
  fd1qd1_hd clk_r_REG69_S5 ( .D(z_m[5]), .CK(n754), .Q(n26) );
  fd1qd1_hd clk_r_REG71_S7 ( .D(z_m[3]), .CK(n754), .Q(n24) );
  fd1qd1_hd clk_r_REG182_S5 ( .D(b_e[1]), .CK(n755), .Q(n587) );
  fd1qd1_hd clk_r_REG183_S5 ( .D(b_e[2]), .CK(n755), .Q(n586) );
  fd1qd1_hd clk_r_REG184_S5 ( .D(b_e[3]), .CK(n755), .Q(n585) );
  fd1qd1_hd clk_r_REG185_S5 ( .D(b_e[4]), .CK(n755), .Q(n584) );
  fd1qd1_hd clk_r_REG209_S5 ( .D(N543), .CK(n756), .Q(n607) );
  fd1qd1_hd clk_r_REG210_S5 ( .D(n293), .CK(n756), .Q(n687) );
  fd1qd1_hd clk_r_REG211_S5 ( .D(n293), .CK(n757), .Q(n688) );
  fd1eqd1_hd clk_r_REG214_S5 ( .D(n763), .E(n782), .CK(i_CLK), .Q(n129) );
  fd1eqd1_hd clk_r_REG278_S1 ( .D(n761), .E(n785), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1eqd1_hd clk_r_REG279_S1 ( .D(n759), .E(n787), .CK(i_CLK), .Q(o_Z_STB) );
  fd1eqd1_hd clk_r_REG246_S2 ( .D(n662), .E(n660), .CK(n757), .Q(n661) );
  fd1eqd1_hd clk_r_REG1_S2 ( .D(n686), .E(n660), .CK(n757), .Q(n565) );
  fd1eqd1_hd clk_r_REG76_S12 ( .D(round_bit), .E(N667), .CK(n754), .Q(n14) );
  fd1eqd1_hd clk_r_REG75_S11 ( .D(guard), .E(N667), .CK(n754), .Q(n13) );
  float_adder_DW01_inc_0 add_x_6 ( .A({n44, n43, n42, n41, n40, n39, n38, n37, 
        n36, n35, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, n563, 
        n23, n22}), .SUM({N431, N430, N429, N428, N427, N426, N425, N424, N423, 
        N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, 
        N410, N409, N408}) );
  float_adder_DP_OP_131_125_8359_0 DP_OP_131_125_8359 ( .I1(i_B[30:23]), .O1({
        n560, n559, n558, n557, n556, n555, n554, n553, n552}), .U488_Y(1'b0), 
        .i_CLK(i_CLK), .IN0(n748) );
  float_adder_DP_OP_132_126_1283_0 DP_OP_132_126_1283 ( .I1({n19, n132, n127, 
        n582, n583, n584, n585, n586, n587, n65}), .O1({n551, n550, n549, n548, 
        n547, n546, n545, n544, n543, n542}) );
  float_adder_DP_OP_128_128_163_0 DP_OP_128_128_163 ( .I1(i_A[30:23]), .O1({
        C1_DATA1_8, C1_DATA1_7, C1_DATA1_6, C1_DATA1_5, C1_DATA1_4, C1_DATA1_3, 
        C1_DATA1_2, C1_DATA1_1, C1_DATA1_0}), .U488_Y(1'b0), .i_CLK(i_CLK), 
        .IN0(n748) );
  float_adder_DP_OP_129_129_1948_0 DP_OP_129_129_1948 ( .I1({n18, n131, n128, 
        n576, n577, n578, n579, n580, n581, n66}), .O1({C1_DATA2_9, C1_DATA2_8, 
        C1_DATA2_7, C1_DATA2_6, C1_DATA2_5, C1_DATA2_4, C1_DATA2_3, C1_DATA2_2, 
        C1_DATA2_1, C1_DATA2_0}) );
  float_adder_DP_OP_143_130_3257_0 DP_OP_143_130_3257 ( .I1({n111, n112, n113, 
        n114, n121, n122, n123, n124, n125, n126}), .I2(n92), .O1({C85_DATA2_9, 
        C85_DATA2_8, C85_DATA2_7, C85_DATA2_6, C85_DATA2_5, C85_DATA2_4, 
        C85_DATA2_3, C85_DATA2_2, C85_DATA2_1, C85_DATA2_0}) );
  float_adder_DP_OP_43_133_2142_0 DP_OP_43_133_2142 ( .I1({C2_Z_26, C2_Z_25, 
        C2_Z_24, C2_Z_23, C2_Z_22, C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, 
        C2_Z_16, C2_Z_15, C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, 
        C2_Z_8, C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0}), .I2({C3_Z_26, C3_Z_25, C3_Z_24, C3_Z_23, C3_Z_22, C3_Z_21, C3_Z_20, C3_Z_19, 
        C3_Z_18, C3_Z_17, C3_Z_16, C3_Z_15, C3_Z_14, C3_Z_13, C3_Z_12, C3_Z_11, 
        C3_Z_10, C3_Z_9, C3_Z_8, C3_Z_7, C3_Z_6, C3_Z_5, C3_Z_4, C3_Z_3, 
        C3_Z_2, C3_Z_1, C3_Z_0}), .I3(n541), .O1(sum) );
  float_adder_DW_cmp_6 gte_x_3 ( .A({1'b0, n67, n68, n69, n70, n71, n72, n73, 
        n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n108, n109, n110, 
        n115, n116, n117, n570, n568, n567}), .B({N543, n45, n46, n47, n48, 
        n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, 
        n63, n64, n118, n119, n120, n574, n572, n571}), .TC(1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b1), .GE_LT_GT_LE(N220), .U780_Y(1'b0), .i_CLK(i_CLK), .U786_Y(
        1'b0), .IN0(n757), .IN1(n756), .IN2(n743) );
  SNPS_CLOCK_GATE_HIGH_float_adder_12_0 clk_gate_clk_r_REG74_S10_0 ( .CLK(
        i_CLK), .EN(n789), .ENCLK(n758), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_10_0 clk_gate_clk_r_REG213_S5 ( .CLK(i_CLK), 
        .EN(N545), .ENCLK(n757), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_9_0 clk_gate_clk_r_REG212_S5 ( .CLK(i_CLK), 
        .EN(N573), .ENCLK(n756), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_7_0 clk_gate_clk_r_REG182_S5_0 ( .CLK(i_CLK), .EN(N585), .ENCLK(n755), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_6_0 clk_gate_clk_r_REG75_S11_0 ( .CLK(i_CLK), .EN(N664), .ENCLK(n754), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_5_0 clk_gate_clk_r_REG142_S5_0 ( .CLK(i_CLK), .EN(n573), .ENCLK(n753), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_4_0 clk_gate_clk_r_REG123_S2_0 ( .CLK(i_CLK), .EN(n569), .ENCLK(n752), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_3_0 clk_gate_clk_r_REG110_S3_0 ( .CLK(i_CLK), .EN(n741), .ENCLK(n751), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_2_0 clk_gate_clk_r_REG21_S22_0 ( .CLK(i_CLK), .EN(N87), .ENCLK(n750), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_1_0 clk_gate_clk_r_REG22_S21_0 ( .CLK(i_CLK), .EN(N596), .ENCLK(n749), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_adder_0_0 clk_gate_clk_r_REG247_S1 ( .CLK(i_CLK), 
        .EN(N516), .ENCLK(n748), .TE(1'b0) );
  fd1qd1_hd R_0_clk_r_REG208_S5 ( .D(N543), .CK(n757), .Q(n743) );
  fd1qd1_hd clk_r_REG171_S5 ( .D(a_m[23]), .CK(n752), .Q(n69) );
  ivd16_hd U8 ( .A(n729), .Y(n486) );
  clknd2d1_hd U18 ( .A(n443), .B(n19), .Y(n771) );
  nd2bd1_hd U19 ( .AN(n513), .B(n486), .Y(n179) );
  nr2bd1_hd U21 ( .AN(N47), .B(n695), .Y(N516) );
  oa21d1_hd U40 ( .A(n422), .B(n293), .C(n332), .Y(N596) );
  nr3d1_hd U41 ( .A(n130), .B(n440), .C(n439), .Y(N87) );
  nr4d2_hd U42 ( .A(n605), .B(n129), .C(n566), .D(n425), .Y(n741) );
  ivd1_hd U43 ( .A(n760), .Y(n759) );
  clknd2d1_hd U44 ( .A(n5), .B(n786), .Y(n760) );
  ivd1_hd U45 ( .A(n762), .Y(n761) );
  clknd2d1_hd U46 ( .A(n4), .B(n784), .Y(n762) );
  ivd1_hd U47 ( .A(n764), .Y(n763) );
  clknd2d1_hd U48 ( .A(n1), .B(n781), .Y(n764) );
  oa21d1_hd U49 ( .A(n401), .B(n402), .C(n403), .Y(N585) );
  ivd1_hd U50 ( .A(n409), .Y(n569) );
  ivd1_hd U51 ( .A(n403), .Y(n573) );
  nd2bd1_hd U52 ( .AN(N667), .B(n228), .Y(N664) );
  ao21d1_hd U58 ( .A(n129), .B(n765), .C(n766), .Y(n781) );
  oa211d1_hd U59 ( .A(n783), .B(n129), .C(n1), .D(n605), .Y(n766) );
  ao21d1_hd U60 ( .A(n566), .B(n425), .C(n767), .Y(n765) );
  ao211d1_hd U61 ( .A(n130), .B(n768), .C(n566), .D(n769), .Y(n767) );
  ad4d1_hd U62 ( .A(n445), .B(n770), .C(n771), .D(n772), .Y(n769) );
  ao211d1_hd U63 ( .A(n65), .B(n469), .C(n130), .D(n444), .Y(n772) );
  nr2d1_hd U64 ( .A(n471), .B(n773), .Y(n770) );
  nd3d1_hd U65 ( .A(n456), .B(n478), .C(n441), .Y(n773) );
  oa21d1_hd U66 ( .A(n774), .B(n436), .C(n111), .Y(n768) );
  scg12d1_hd U67 ( .A(n336), .B(n338), .C(n125), .Y(n774) );
  scg15d1_hd U68 ( .A(n605), .B(n783), .C(n1), .D(n775), .Y(n782) );
  nd3d1_hd U69 ( .A(n566), .B(n431), .C(n776), .Y(n775) );
  nr2d1_hd U70 ( .A(n130), .B(n605), .Y(n776) );
  nd2bd1_hd U71 ( .AN(n425), .B(n566), .Y(n783) );
  ad2d1_hd U72 ( .A(n695), .B(n4), .Y(n784) );
  nd2bd1_hd U73 ( .AN(N47), .B(n4), .Y(n785) );
  ad2d1_hd U74 ( .A(n728), .B(n5), .Y(n786) );
  nd2bd1_hd U75 ( .AN(N87), .B(n5), .Y(n787) );
  oa22ad1_hd U76 ( .A(n777), .B(n778), .C(n778), .D(n484), .Y(n789) );
  or2d1_hd U77 ( .A(n129), .B(n130), .Y(n778) );
  ao22d1_hd U78 ( .A(n566), .B(n434), .C(n605), .D(n484), .Y(n777) );
  oa21d1_hd U79 ( .A(n293), .B(n779), .C(n780), .Y(n795) );
  ao22d1_hd U80 ( .A(n660), .B(C1_DATA1_8), .C(C1_DATA2_9), .D(n393), .Y(n780)
         );
  nr2d1_hd U81 ( .A(n393), .B(n660), .Y(n779) );
endmodule


module float_multiplier_DW01_inc_0 ( A, SUM );
  input [23:0] A;
  output [23:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;

  had1_hd U2 ( .A(A[22]), .B(n2), .CO(n1), .S(SUM[22]) );
  had1_hd U3 ( .A(A[21]), .B(n3), .CO(n2), .S(SUM[21]) );
  had1_hd U4 ( .A(A[20]), .B(n4), .CO(n3), .S(SUM[20]) );
  had1_hd U5 ( .A(A[19]), .B(n5), .CO(n4), .S(SUM[19]) );
  had1_hd U6 ( .A(A[18]), .B(n6), .CO(n5), .S(SUM[18]) );
  had1_hd U7 ( .A(A[17]), .B(n7), .CO(n6), .S(SUM[17]) );
  had1_hd U8 ( .A(A[16]), .B(n8), .CO(n7), .S(SUM[16]) );
  had1_hd U9 ( .A(A[15]), .B(n9), .CO(n8), .S(SUM[15]) );
  had1_hd U10 ( .A(A[14]), .B(n10), .CO(n9), .S(SUM[14]) );
  had1_hd U11 ( .A(A[13]), .B(n11), .CO(n10), .S(SUM[13]) );
  had1_hd U12 ( .A(A[12]), .B(n12), .CO(n11), .S(SUM[12]) );
  had1_hd U13 ( .A(A[11]), .B(n13), .CO(n12), .S(SUM[11]) );
  had1_hd U14 ( .A(A[10]), .B(n14), .CO(n13), .S(SUM[10]) );
  had1_hd U15 ( .A(A[9]), .B(n15), .CO(n14), .S(SUM[9]) );
  had1_hd U16 ( .A(A[8]), .B(n16), .CO(n15), .S(SUM[8]) );
  had1_hd U17 ( .A(A[7]), .B(n17), .CO(n16), .S(SUM[7]) );
  had1_hd U18 ( .A(A[6]), .B(n18), .CO(n17), .S(SUM[6]) );
  had1_hd U19 ( .A(A[5]), .B(n19), .CO(n18), .S(SUM[5]) );
  had1_hd U20 ( .A(A[4]), .B(n20), .CO(n19), .S(SUM[4]) );
  had1_hd U21 ( .A(A[3]), .B(n21), .CO(n20), .S(SUM[3]) );
  had1_hd U22 ( .A(A[2]), .B(n22), .CO(n21), .S(SUM[2]) );
  had1_hd U23 ( .A(A[1]), .B(A[0]), .CO(n22), .S(SUM[1]) );
  xo2d1_hd U27 ( .A(n1), .B(A[23]), .Y(SUM[23]) );
  ivd1_hd U28 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module float_multiplier_DP_OP_114_130_61_0 ( I1, I2, I3, I4, I5, I6, O1 );
  input [9:0] I1;
  input [9:0] I2;
  input [9:0] I4;
  output [9:0] O1;
  input I3, I5, I6;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n87, n88;

  fad1_hd U3 ( .A(n32), .B(I6), .CI(n3), .CO(n2), .S(O1[8]) );
  fad1_hd U4 ( .A(n31), .B(I6), .CI(n4), .CO(n3), .S(O1[7]) );
  fad1_hd U5 ( .A(n30), .B(I6), .CI(n5), .CO(n4), .S(O1[6]) );
  fad1_hd U6 ( .A(n29), .B(I6), .CI(n6), .CO(n5), .S(O1[5]) );
  fad1_hd U7 ( .A(n28), .B(I6), .CI(n7), .CO(n6), .S(O1[4]) );
  fad1_hd U8 ( .A(n27), .B(I6), .CI(n8), .CO(n7), .S(O1[3]) );
  fad1_hd U9 ( .A(n26), .B(I6), .CI(n9), .CO(n8), .S(O1[2]) );
  fad1_hd U10 ( .A(n10), .B(I6), .CI(n25), .CO(n9), .S(O1[1]) );
  fad1_hd U24 ( .A(I1[8]), .B(I2[8]), .CI(n13), .CO(n12), .S(n42) );
  fad1_hd U25 ( .A(I1[7]), .B(I2[7]), .CI(n14), .CO(n13), .S(n41) );
  fad1_hd U26 ( .A(I1[6]), .B(I2[6]), .CI(n15), .CO(n14), .S(n40) );
  fad1_hd U27 ( .A(I1[5]), .B(I2[5]), .CI(n16), .CO(n15), .S(n39) );
  fad1_hd U28 ( .A(I1[4]), .B(I2[4]), .CI(n17), .CO(n16), .S(n38) );
  fad1_hd U29 ( .A(I1[3]), .B(I2[3]), .CI(n18), .CO(n17), .S(n37) );
  fad1_hd U30 ( .A(I1[2]), .B(I2[2]), .CI(n19), .CO(n18), .S(n36) );
  fad1_hd U31 ( .A(I1[1]), .B(I2[1]), .CI(n20), .CO(n19), .S(n35) );
  had1_hd U32 ( .A(I2[0]), .B(I1[0]), .CO(n20), .S(n34) );
  scg2d1_hd U35 ( .A(I5), .B(I4[8]), .C(I3), .D(n42), .Y(n32) );
  scg2d1_hd U36 ( .A(I5), .B(I4[7]), .C(I3), .D(n41), .Y(n31) );
  scg2d1_hd U37 ( .A(I5), .B(I4[6]), .C(I3), .D(n40), .Y(n30) );
  scg2d1_hd U38 ( .A(I4[9]), .B(I5), .C(n88), .D(I3), .Y(n87) );
  scg2d1_hd U39 ( .A(I5), .B(I4[1]), .C(I3), .D(n35), .Y(n25) );
  scg2d1_hd U40 ( .A(I5), .B(I4[2]), .C(I3), .D(n36), .Y(n26) );
  scg2d1_hd U41 ( .A(I5), .B(I4[3]), .C(I3), .D(n37), .Y(n27) );
  scg2d1_hd U42 ( .A(I5), .B(I4[4]), .C(I3), .D(n38), .Y(n28) );
  scg2d1_hd U43 ( .A(I5), .B(I4[5]), .C(I3), .D(n39), .Y(n29) );
  xo3d1_hd U44 ( .A(I6), .B(n2), .C(n87), .Y(O1[9]) );
  xo3d1_hd U45 ( .A(n12), .B(I1[9]), .C(I2[9]), .Y(n88) );
  ivd1_hd U46 ( .A(O1[0]), .Y(n10) );
  ao22d1_hd U47 ( .A(I5), .B(I4[0]), .C(I3), .D(n34), .Y(O1[0]) );
endmodule


module float_multiplier_DW_mult_uns_2 ( a, b, product );
  input [23:0] a;
  input [23:0] b;
  output [47:0] product;
  wire   n1, n3, n5, n9, n11, n13, n15, n19, n21, n23, n25, n29, n31, n33, n35,
         n39, n41, n43, n45, n49, n51, n53, n55, n59, n61, n63, n65, n69, n71,
         n73, n75, n79, n81, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n179, n180, n181, n182, n183, n185, n187,
         n188, n189, n190, n191, n193, n195, n196, n197, n198, n199, n201,
         n203, n204, n205, n206, n207, n209, n211, n212, n213, n214, n215,
         n217, n219, n220, n221, n222, n223, n225, n227, n228, n229, n230,
         n231, n233, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n297, n299, n300, n301, n302,
         n304, n307, n308, n309, n310, n312, n314, n315, n316, n317, n318,
         n319, n320, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n339, n341, n342, n343,
         n344, n345, n346, n347, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n366, n368,
         n369, n371, n373, n374, n375, n377, n379, n380, n381, n382, n383,
         n385, n387, n388, n389, n390, n391, n393, n395, n396, n398, n399,
         n400, n401, n403, n405, n407, n409, n411, n413, n415, n417, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n431,
         n433, n434, n435, n436, n438, n439, n440, n441, n445, n447, n450,
         n451, n452, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n866, n869, n872, n875, n878, n881, n884, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n971, n972, n973, n974, n975, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n993, n994, n995, n996, n997, n998, n999, n1000, n1003, n1004,
         n1005, n1006, n1007, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1083, n1085, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1761, n1762,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030;

  fad2_hd U606 ( .A(n1295), .B(n669), .CI(n1223), .CO(n653), .S(n654) );
  ivd1_hd U1732 ( .A(n943), .Y(n941) );
  clknd2d1_hd U1733 ( .A(n965), .B(n951), .Y(n945) );
  ivd1_hd U1734 ( .A(n945), .Y(n947) );
  ao21d1_hd U1735 ( .A(n966), .B(n951), .C(n952), .Y(n946) );
  ivd1_hd U1736 ( .A(n946), .Y(n948) );
  ivd1_hd U1737 ( .A(n942), .Y(n940) );
  xn2d1_hd U1738 ( .A(n901), .B(n1044), .Y(n2006) );
  clknd2d1_hd U1739 ( .A(n1056), .B(n1048), .Y(n1046) );
  nr2d1_hd U1740 ( .A(n1063), .B(n1058), .Y(n1056) );
  nr2bd2_hd U1741 ( .AN(n1817), .B(n1825), .Y(n35) );
  nr2d2_hd U1742 ( .A(n1833), .B(n1817), .Y(n33) );
  ivd1_hd U1743 ( .A(n1066), .Y(n1065) );
  xo2d1_hd U1744 ( .A(n1052), .B(n902), .Y(n2005) );
  ivd1_hd U1746 ( .A(a[23]), .Y(n918) );
  xo2d1_hd U1749 ( .A(b[20]), .B(b[19]), .Y(n1830) );
  nr2bd2_hd U1750 ( .AN(n1814), .B(n1822), .Y(n65) );
  xn2d1_hd U1751 ( .A(b[19]), .B(b[18]), .Y(n1822) );
  fad1_hd U1752 ( .A(n1175), .B(n1199), .CI(n656), .CO(n651), .S(n652) );
  fad1_hd U1753 ( .A(n627), .B(n1148), .CI(n614), .CO(n609), .S(n610) );
  xo2d1_hd U1754 ( .A(b[14]), .B(n1492), .Y(n1202) );
  xo2d1_hd U1755 ( .A(n985), .B(n894), .Y(n2013) );
  fad1_hd U1756 ( .A(n696), .B(n1226), .CI(n1298), .CO(n691), .S(n692) );
  xo2d1_hd U1757 ( .A(b[5]), .B(n1646), .Y(n1281) );
  xo2d1_hd U1758 ( .A(b[2]), .B(n1694), .Y(n1304) );
  xo2d1_hd U1759 ( .A(b[11]), .B(n1550), .Y(n1235) );
  xo2d1_hd U1760 ( .A(b[2]), .B(n1697), .Y(n1307) );
  xo2d1_hd U1761 ( .A(b[5]), .B(n1648), .Y(n1283) );
  nr2d2_hd U1762 ( .A(n1835), .B(n1819), .Y(n13) );
  xo2d1_hd U1763 ( .A(b[5]), .B(b[4]), .Y(n1835) );
  xn2d1_hd U1764 ( .A(b[2]), .B(b[3]), .Y(n1819) );
  nr2bd2_hd U1765 ( .AN(n1819), .B(n1827), .Y(n15) );
  xn2d1_hd U1766 ( .A(n907), .B(n1074), .Y(n2000) );
  oa21d1_hd U1767 ( .A(n1076), .B(n1078), .C(n1077), .Y(n1075) );
  fad1_hd U1768 ( .A(n1262), .B(n814), .CI(n1286), .CO(n811), .S(n812) );
  xo2d1_hd U1769 ( .A(b[11]), .B(n1553), .Y(n1238) );
  xn2d1_hd U1770 ( .A(n903), .B(n1055), .Y(n2004) );
  ivd1_hd U1771 ( .A(n1075), .Y(n1074) );
  clknd2d1_hd U1772 ( .A(n2023), .B(n1078), .Y(n1761) );
  nr2d2_hd U1774 ( .A(n1836), .B(n1820), .Y(n3) );
  xn2d1_hd U1775 ( .A(n1078), .B(n908), .Y(n1999) );
  nr2d1_hd U1777 ( .A(n924), .B(n918), .Y(n916) );
  nr2d1_hd U1778 ( .A(n974), .B(n971), .Y(n965) );
  ivd1_hd U1779 ( .A(n1028), .Y(n1094) );
  nr2d1_hd U1780 ( .A(n1013), .B(n979), .Y(n977) );
  clknd2d1_hd U1781 ( .A(n947), .B(n940), .Y(n938) );
  oa21d1_hd U1783 ( .A(n2018), .B(n29), .C(n1610), .Y(n1584) );
  oa21d1_hd U1784 ( .A(n1999), .B(n49), .C(n1526), .Y(n1500) );
  ao21d1_hd U1785 ( .A(n1065), .B(n1056), .C(n1057), .Y(n1055) );
  xo2d1_hd U1786 ( .A(n919), .B(n918), .Y(n2020) );
  xo2d1_hd U1787 ( .A(n944), .B(n889), .Y(n2017) );
  xo2d1_hd U1788 ( .A(b[17]), .B(n1440), .Y(n1175) );
  fad1_hd U1789 ( .A(n1154), .B(n698), .CI(n1178), .CO(n695), .S(n696) );
  oa21d1_hd U1790 ( .A(n2007), .B(n39), .C(n1570), .Y(n1544) );
  xo2d1_hd U1791 ( .A(n1023), .B(n898), .Y(n2009) );
  xo2d1_hd U1792 ( .A(n1041), .B(n900), .Y(n2007) );
  fad1_hd U1793 ( .A(n1146), .B(n1170), .CI(n585), .CO(n582), .S(n583) );
  xo2d1_hd U1794 ( .A(b[8]), .B(n1596), .Y(n1256) );
  xn2d1_hd U1795 ( .A(n904), .B(n1060), .Y(n2003) );
  xo2d1_hd U1796 ( .A(n1071), .B(n906), .Y(n2001) );
  fad1_hd U1797 ( .A(n1281), .B(n1305), .CI(n783), .CO(n771), .S(n772) );
  fad1_hd U1798 ( .A(n1235), .B(n794), .CI(n1259), .CO(n791), .S(n792) );
  ad3d2_hd U1799 ( .A(n1836), .B(n1828), .C(n1820), .Y(n11) );
  or2bd2_hd U1800 ( .B(n1820), .AN(n1836), .Y(n9) );
  clknd2d1_hd U1801 ( .A(n399), .B(n401), .Y(n398) );
  nr2d1_hd U1802 ( .A(a[14]), .B(a[15]), .Y(n990) );
  nr2d1_hd U1803 ( .A(n942), .B(n935), .Y(n933) );
  oa21d1_hd U1804 ( .A(n971), .B(n975), .C(n972), .Y(n966) );
  nr2d1_hd U1805 ( .A(n1042), .B(n1039), .Y(n1033) );
  oa21d1_hd U1806 ( .A(n1014), .B(n979), .C(n980), .Y(n978) );
  ao21d1_hd U1807 ( .A(n948), .B(n940), .C(n941), .Y(n939) );
  xn2d1_hd U1808 ( .A(b[12]), .B(b[11]), .Y(n1816) );
  oa21d1_hd U1809 ( .A(n2004), .B(n69), .C(n1417), .Y(n1391) );
  oa21d1_hd U1810 ( .A(n1999), .B(n69), .C(n1422), .Y(n1396) );
  clknd2d1_hd U1811 ( .A(n1033), .B(n1094), .Y(n1024) );
  ao21d2_hd U1812 ( .A(n1045), .B(n977), .C(n978), .Y(n1) );
  nr2bd2_hd U1813 ( .AN(n1813), .B(n1821), .Y(n75) );
  or2bd2_hd U1814 ( .B(n1814), .AN(n1830), .Y(n69) );
  oa21d1_hd U1816 ( .A(n1970), .B(n19), .C(n1659), .Y(n1633) );
  oa21d1_hd U1817 ( .A(n1970), .B(n9), .C(n1711), .Y(n1685) );
  oa21d1_hd U1818 ( .A(n2018), .B(n19), .C(n1662), .Y(n1636) );
  xo2d1_hd U1819 ( .A(n973), .B(n892), .Y(n2014) );
  xo2d1_hd U1820 ( .A(n962), .B(n891), .Y(n2015) );
  xo2d1_hd U1821 ( .A(n1005), .B(n896), .Y(n2011) );
  or2bd2_hd U1822 ( .B(n1817), .AN(n1833), .Y(n39) );
  or2bd2_hd U1824 ( .B(n1818), .AN(n1834), .Y(n29) );
  scg9d1_hd U1825 ( .A(n1), .B(n1972), .C(n2024), .Y(n1970) );
  xo2d1_hd U1826 ( .A(n937), .B(n888), .Y(n2018) );
  fad1_hd U1827 ( .A(n599), .B(n586), .CI(n1122), .CO(n584), .S(n585) );
  fad1_hd U1828 ( .A(n858), .B(b[2]), .CI(n1124), .CO(n613), .S(n614) );
  fad1_hd U1829 ( .A(n859), .B(b[2]), .CI(n1149), .CO(n627), .S(n628) );
  xo2d1_hd U1830 ( .A(b[2]), .B(n1688), .Y(n1298) );
  had1_hd U1831 ( .A(n1156), .B(n735), .CO(n723), .S(n724) );
  oa21d1_hd U1832 ( .A(n2007), .B(n29), .C(n1622), .Y(n1596) );
  oa21d1_hd U1833 ( .A(n2007), .B(n19), .C(n1674), .Y(n1648) );
  oa21d1_hd U1834 ( .A(n2006), .B(n19), .C(n1675), .Y(n1649) );
  fad1_hd U1835 ( .A(n559), .B(n548), .CI(n1119), .CO(n546), .S(n547) );
  fad1_hd U1836 ( .A(n1121), .B(n1145), .CI(n584), .CO(n569), .S(n570) );
  fad1_hd U1837 ( .A(n1181), .B(n736), .CI(n1205), .CO(n733), .S(n734) );
  fad1_hd U1838 ( .A(n1208), .B(n768), .CI(n1232), .CO(n765), .S(n766) );
  had1_hd U1839 ( .A(n819), .B(n1238), .CO(n813), .S(n814) );
  xo2d1_hd U1840 ( .A(n1065), .B(n905), .Y(n2002) );
  fad1_hd U1841 ( .A(n1304), .B(n775), .CI(n1256), .CO(n763), .S(n764) );
  fad1_hd U1842 ( .A(n1307), .B(n799), .CI(n1283), .CO(n789), .S(n790) );
  had1_hd U1843 ( .A(n831), .B(n1265), .CO(n827), .S(n828) );
  nr2bd2_hd U1844 ( .AN(n1820), .B(n1828), .Y(n5) );
  had1_hd U1845 ( .A(n837), .B(n1292), .CO(n835), .S(n836) );
  clknd2d1_hd U1846 ( .A(n629), .B(n616), .Y(n265) );
  nr2d1_hd U1848 ( .A(n398), .B(n1983), .Y(n396) );
  ao21d2_hd U1852 ( .A(n196), .B(n2027), .C(n193), .Y(n191) );
  had1_hd U1861 ( .A(n711), .B(n1130), .CO(n697), .S(n698) );
  xo2d1_hd U1862 ( .A(b[23]), .B(n1345), .Y(n1130) );
  oa21d1_hd U1863 ( .A(n79), .B(n1761), .C(n1974), .Y(n1345) );
  had1_hd U1864 ( .A(b[20]), .B(n1158), .CO(n747), .S(n748) );
  xo2d1_hd U1865 ( .A(b[20]), .B(n1398), .Y(n1158) );
  oa21d1_hd U1866 ( .A(n69), .B(n1762), .C(n1997), .Y(n1398) );
  had1_hd U1868 ( .A(b[14]), .B(n1212), .CO(n801), .S(n802) );
  xo2d1_hd U1869 ( .A(b[14]), .B(n1502), .Y(n1212) );
  oa21d1_hd U1870 ( .A(n49), .B(n1762), .C(n1995), .Y(n1502) );
  oa21d1_hd U1871 ( .A(n1058), .B(n1064), .C(n1059), .Y(n1057) );
  oa21d1_hd U1872 ( .A(n2001), .B(n79), .C(n1368), .Y(n1342) );
  ao222d1_hd U1873 ( .A(n73), .B(a[4]), .C(n75), .D(a[3]), .E(n81), .F(a[2]), 
        .Y(n1368) );
  ao222d1_hd U1874 ( .A(n63), .B(a[7]), .C(n65), .D(a[6]), .E(n71), .F(a[5]), 
        .Y(n1417) );
  ivd1_hd U1875 ( .A(n856), .Y(n586) );
  xo2d1_hd U1876 ( .A(b[23]), .B(n1337), .Y(n1122) );
  oa21d1_hd U1877 ( .A(n2006), .B(n79), .C(n1363), .Y(n1337) );
  ad2d1_hd U1878 ( .A(b[23]), .B(a[4]), .Y(n858) );
  xo2d1_hd U1879 ( .A(b[23]), .B(n1339), .Y(n1124) );
  oa21d1_hd U1880 ( .A(n2004), .B(n79), .C(n1365), .Y(n1339) );
  clknd2d1_hd U1881 ( .A(n21), .B(a[23]), .Y(n1659) );
  ao222d1_hd U1882 ( .A(n23), .B(a[22]), .C(n25), .D(a[21]), .E(n31), .F(a[20]), .Y(n1610) );
  ad2d1_hd U1883 ( .A(b[23]), .B(a[3]), .Y(n859) );
  xo2d1_hd U1884 ( .A(b[20]), .B(n1389), .Y(n1149) );
  oa21d1_hd U1885 ( .A(n2006), .B(n69), .C(n1415), .Y(n1389) );
  ao222d1_hd U1886 ( .A(n13), .B(a[22]), .C(n15), .D(a[21]), .E(n21), .F(a[20]), .Y(n1662) );
  xo2d1_hd U1887 ( .A(b[17]), .B(n1443), .Y(n1178) );
  xo2d1_hd U1888 ( .A(b[20]), .B(n1394), .Y(n1154) );
  oa21d1_hd U1889 ( .A(n2004), .B(n59), .C(n1469), .Y(n1443) );
  xo2d1_hd U1890 ( .A(b[20]), .B(n1396), .Y(n1156) );
  ao222d1_hd U1891 ( .A(n63), .B(a[2]), .C(n65), .D(a[1]), .E(n71), .F(a[0]), 
        .Y(n1422) );
  oa21d1_hd U1892 ( .A(n2001), .B(n59), .C(n1472), .Y(n1446) );
  ao222d1_hd U1893 ( .A(n53), .B(a[4]), .C(n55), .D(a[3]), .E(n61), .F(a[2]), 
        .Y(n1472) );
  had1_hd U1894 ( .A(n777), .B(n1184), .CO(n767), .S(n768) );
  xo2d1_hd U1895 ( .A(b[17]), .B(n1449), .Y(n1184) );
  oa21d1_hd U1896 ( .A(n59), .B(n1761), .C(n1989), .Y(n1449) );
  oa21d1_hd U1897 ( .A(n2001), .B(n49), .C(n1524), .Y(n1498) );
  ao222d1_hd U1898 ( .A(n43), .B(a[4]), .C(n45), .D(a[3]), .E(n51), .F(a[2]), 
        .Y(n1524) );
  oa21d1_hd U1899 ( .A(n1043), .B(n1039), .C(n1040), .Y(n1034) );
  nr2d1_hd U1901 ( .A(a[20]), .B(a[21]), .Y(n942) );
  ao21d1_hd U1902 ( .A(n1057), .B(n1048), .C(n1049), .Y(n1047) );
  oa21d1_hd U1903 ( .A(n1050), .B(n1054), .C(n1051), .Y(n1049) );
  fad1_hd U1905 ( .A(n573), .B(n856), .CI(n1241), .CO(n571), .S(n572) );
  ivd1_hd U1906 ( .A(n855), .Y(n573) );
  xo2d1_hd U1907 ( .A(b[8]), .B(n1581), .Y(n1241) );
  oa21d1_hd U1908 ( .A(n1970), .B(n29), .C(n1607), .Y(n1581) );
  xo2d1_hd U1909 ( .A(b[2]), .B(n1685), .Y(n1295) );
  xo2d1_hd U1910 ( .A(b[11]), .B(n1538), .Y(n1223) );
  xo2d1_hd U1912 ( .A(b[14]), .B(n1500), .Y(n1210) );
  ao222d1_hd U1913 ( .A(n43), .B(a[2]), .C(n45), .D(a[1]), .E(n51), .F(a[0]), 
        .Y(n1526) );
  oa21d1_hd U1914 ( .A(n2001), .B(n39), .C(n1576), .Y(n1550) );
  ao222d1_hd U1915 ( .A(n33), .B(a[4]), .C(n35), .D(a[3]), .E(n41), .F(a[2]), 
        .Y(n1576) );
  oa21d1_hd U1916 ( .A(n39), .B(n1761), .C(n1987), .Y(n1553) );
  oa21d1_hd U1917 ( .A(n2001), .B(n29), .C(n1628), .Y(n1602) );
  ao222d1_hd U1918 ( .A(n23), .B(a[4]), .C(n25), .D(a[3]), .E(n31), .F(a[2]), 
        .Y(n1628) );
  oa21d1_hd U1919 ( .A(n2006), .B(n59), .C(n1467), .Y(n1441) );
  ao222d1_hd U1920 ( .A(n53), .B(a[9]), .C(n55), .D(a[8]), .E(n61), .F(a[7]), 
        .Y(n1467) );
  oa21d1_hd U1921 ( .A(n2001), .B(n69), .C(n1420), .Y(n1394) );
  ao222d1_hd U1922 ( .A(n63), .B(a[4]), .C(n65), .D(a[3]), .E(n71), .F(a[2]), 
        .Y(n1420) );
  oa21d1_hd U1923 ( .A(n2018), .B(n49), .C(n1506), .Y(n1480) );
  ao222d1_hd U1924 ( .A(n43), .B(a[22]), .C(n45), .D(a[21]), .E(n51), .F(a[20]), .Y(n1506) );
  oa21d1_hd U1926 ( .A(n2018), .B(n39), .C(n1558), .Y(n1532) );
  ao222d1_hd U1927 ( .A(n33), .B(a[22]), .C(n35), .D(a[21]), .E(n41), .F(a[20]), .Y(n1558) );
  oa21d1_hd U1928 ( .A(n2009), .B(n59), .C(n1464), .Y(n1438) );
  ao222d1_hd U1929 ( .A(n53), .B(a[12]), .C(n55), .D(a[11]), .E(n61), .F(a[10]), .Y(n1464) );
  oa21d1_hd U1930 ( .A(n2009), .B(n49), .C(n1516), .Y(n1490) );
  ao222d1_hd U1931 ( .A(n43), .B(a[12]), .C(n45), .D(a[11]), .E(n51), .F(a[10]), .Y(n1516) );
  oa21d1_hd U1932 ( .A(n2006), .B(n49), .C(n1519), .Y(n1493) );
  ao222d1_hd U1933 ( .A(n43), .B(a[9]), .C(n45), .D(a[8]), .E(n51), .F(a[7]), 
        .Y(n1519) );
  oa21d1_hd U1934 ( .A(n2009), .B(n39), .C(n1568), .Y(n1542) );
  ao222d1_hd U1935 ( .A(n33), .B(a[12]), .C(n35), .D(a[11]), .E(n41), .F(a[10]), .Y(n1568) );
  oa21d1_hd U1936 ( .A(n2006), .B(n39), .C(n1571), .Y(n1545) );
  ao222d1_hd U1937 ( .A(n33), .B(a[9]), .C(n35), .D(a[8]), .E(n41), .F(a[7]), 
        .Y(n1571) );
  oa21d1_hd U1938 ( .A(n2009), .B(n29), .C(n1620), .Y(n1594) );
  ao222d1_hd U1939 ( .A(n23), .B(a[12]), .C(n25), .D(a[11]), .E(n31), .F(a[10]), .Y(n1620) );
  nr2d1_hd U1940 ( .A(a[23]), .B(a[22]), .Y(n924) );
  oa21d1_hd U1941 ( .A(n943), .B(n935), .C(n936), .Y(n934) );
  nr2d1_hd U1942 ( .A(a[21]), .B(a[22]), .Y(n935) );
  clknd2d1_hd U1943 ( .A(a[21]), .B(a[22]), .Y(n936) );
  oa21d1_hd U1944 ( .A(n2018), .B(n69), .C(n1402), .Y(n1376) );
  ao222d1_hd U1945 ( .A(n63), .B(a[22]), .C(n65), .D(a[21]), .E(n71), .F(a[20]), .Y(n1402) );
  oa21d1_hd U1946 ( .A(n2018), .B(n59), .C(n1454), .Y(n1428) );
  ao222d1_hd U1947 ( .A(n53), .B(a[22]), .C(n55), .D(a[21]), .E(n61), .F(a[20]), .Y(n1454) );
  fad1_hd U1948 ( .A(n516), .B(n849), .CI(n1187), .CO(n505), .S(n506) );
  ad2d1_hd U1949 ( .A(b[23]), .B(a[13]), .Y(n849) );
  xo2d1_hd U1950 ( .A(b[14]), .B(n1477), .Y(n1187) );
  oa21d1_hd U1951 ( .A(n1970), .B(n49), .C(n1503), .Y(n1477) );
  fad1_hd U1952 ( .A(n548), .B(n852), .CI(n1214), .CO(n535), .S(n536) );
  ad2d1_hd U1953 ( .A(b[23]), .B(a[10]), .Y(n852) );
  xo2d1_hd U1954 ( .A(b[11]), .B(n1529), .Y(n1214) );
  oa21d1_hd U1955 ( .A(n1970), .B(n39), .C(n1555), .Y(n1529) );
  xo2d1_hd U1956 ( .A(b[23]), .B(n1334), .Y(n1119) );
  oa21d1_hd U1957 ( .A(n2009), .B(n79), .C(n1360), .Y(n1334) );
  ao222d1_hd U1958 ( .A(n73), .B(a[12]), .C(n75), .D(a[11]), .E(n81), .F(a[10]), .Y(n1360) );
  xo2d1_hd U1959 ( .A(b[23]), .B(n1336), .Y(n1121) );
  xo2d1_hd U1960 ( .A(b[20]), .B(n1385), .Y(n1145) );
  oa21d1_hd U1961 ( .A(n2007), .B(n79), .C(n1362), .Y(n1336) );
  xo2d1_hd U1962 ( .A(b[20]), .B(n1386), .Y(n1146) );
  xo2d1_hd U1963 ( .A(b[17]), .B(n1435), .Y(n1170) );
  oa21d1_hd U1964 ( .A(n2009), .B(n69), .C(n1412), .Y(n1386) );
  xo2d1_hd U1965 ( .A(b[20]), .B(n1388), .Y(n1148) );
  oa21d1_hd U1966 ( .A(n2007), .B(n69), .C(n1414), .Y(n1388) );
  ao222d1_hd U1967 ( .A(n63), .B(a[10]), .C(n65), .D(a[9]), .E(n71), .F(a[8]), 
        .Y(n1414) );
  xo2d1_hd U1968 ( .A(b[14]), .B(n1489), .Y(n1199) );
  oa21d1_hd U1969 ( .A(n2007), .B(n59), .C(n1466), .Y(n1440) );
  xo2d1_hd U1970 ( .A(b[11]), .B(n1541), .Y(n1226) );
  oa21d1_hd U1971 ( .A(n2018), .B(n9), .C(n1714), .Y(n1688) );
  xo2d1_hd U1972 ( .A(b[8]), .B(n1590), .Y(n1250) );
  oa21d1_hd U1973 ( .A(n2007), .B(n49), .C(n1518), .Y(n1492) );
  xo2d1_hd U1974 ( .A(b[14]), .B(n1495), .Y(n1205) );
  xo2d1_hd U1975 ( .A(b[17]), .B(n1446), .Y(n1181) );
  oa21d1_hd U1976 ( .A(n2004), .B(n49), .C(n1521), .Y(n1495) );
  ao222d1_hd U1977 ( .A(n33), .B(a[10]), .C(n35), .D(a[9]), .E(n41), .F(a[8]), 
        .Y(n1570) );
  xo2d1_hd U1978 ( .A(b[11]), .B(n1547), .Y(n1232) );
  xo2d1_hd U1979 ( .A(b[14]), .B(n1498), .Y(n1208) );
  oa21d1_hd U1980 ( .A(n2004), .B(n39), .C(n1573), .Y(n1547) );
  oa21d1_hd U1981 ( .A(n2006), .B(n29), .C(n1623), .Y(n1597) );
  ao222d1_hd U1982 ( .A(n23), .B(a[9]), .C(n25), .D(a[8]), .E(n31), .F(a[7]), 
        .Y(n1623) );
  ao222d1_hd U1983 ( .A(n13), .B(a[9]), .C(n15), .D(a[8]), .E(n21), .F(a[7]), 
        .Y(n1675) );
  nr2d1_hd U1984 ( .A(a[11]), .B(a[12]), .Y(n1021) );
  ao21d1_hd U1985 ( .A(n1034), .B(n1094), .C(n1027), .Y(n1025) );
  ivd1_hd U1986 ( .A(n1029), .Y(n1027) );
  clknd2d1_hd U1987 ( .A(a[11]), .B(a[12]), .Y(n1022) );
  clknd2d1_hd U1989 ( .A(a[8]), .B(a[9]), .Y(n1043) );
  nr2d1_hd U1990 ( .A(a[8]), .B(a[9]), .Y(n1042) );
  clknd2d1_hd U1991 ( .A(a[9]), .B(a[10]), .Y(n1040) );
  nr2d1_hd U1992 ( .A(a[6]), .B(a[7]), .Y(n1053) );
  clknd2d1_hd U1993 ( .A(a[6]), .B(a[7]), .Y(n1054) );
  nr2d1_hd U1994 ( .A(a[3]), .B(a[4]), .Y(n1069) );
  clknd2d1_hd U1995 ( .A(a[3]), .B(a[4]), .Y(n1070) );
  nr2d1_hd U1996 ( .A(a[2]), .B(a[3]), .Y(n1072) );
  clknd2d1_hd U1997 ( .A(a[2]), .B(a[3]), .Y(n1073) );
  oa21d1_hd U1999 ( .A(n953), .B(n961), .C(n954), .Y(n952) );
  ao21d1_hd U2000 ( .A(n916), .B(n934), .C(n917), .Y(n915) );
  nr2d1_hd U2001 ( .A(n925), .B(n918), .Y(n917) );
  xo2d1_hd U2002 ( .A(b[2]), .B(n1695), .Y(n1305) );
  oa21d1_hd U2003 ( .A(n2009), .B(n19), .C(n1672), .Y(n1646) );
  xo2d1_hd U2004 ( .A(b[8]), .B(n1599), .Y(n1259) );
  oa21d1_hd U2005 ( .A(n2004), .B(n29), .C(n1625), .Y(n1599) );
  xo2d1_hd U2006 ( .A(b[5]), .B(n1651), .Y(n1286) );
  xo2d1_hd U2007 ( .A(b[8]), .B(n1602), .Y(n1262) );
  oa21d1_hd U2008 ( .A(n2004), .B(n19), .C(n1677), .Y(n1651) );
  xo2d1_hd U2009 ( .A(b[8]), .B(n1605), .Y(n1265) );
  oa21d1_hd U2010 ( .A(n29), .B(n1761), .C(n1986), .Y(n1605) );
  oa21d1_hd U2011 ( .A(n2001), .B(n19), .C(n1680), .Y(n1654) );
  ao222d1_hd U2012 ( .A(n13), .B(a[4]), .C(n15), .D(a[3]), .E(n21), .F(a[2]), 
        .Y(n1680) );
  xo2d1_hd U2014 ( .A(b[5]), .B(n1657), .Y(n1292) );
  oa21d1_hd U2015 ( .A(n19), .B(n1761), .C(n1985), .Y(n1657) );
  clknd2d1_hd U2016 ( .A(n1103), .B(n1077), .Y(n908) );
  ivd1_hd U2017 ( .A(n1076), .Y(n1103) );
  nr2d1_hd U2018 ( .A(n999), .B(n990), .Y(n988) );
  ivd1_hd U2019 ( .A(n997), .Y(n999) );
  ad2d1_hd U2020 ( .A(b[23]), .B(a[9]), .Y(n853) );
  ao222d1_hd U2021 ( .A(n73), .B(a[9]), .C(n75), .D(a[8]), .E(n81), .F(a[7]), 
        .Y(n1363) );
  ao222d1_hd U2022 ( .A(n73), .B(a[7]), .C(n75), .D(a[6]), .E(n81), .F(a[5]), 
        .Y(n1365) );
  ao222d1_hd U2023 ( .A(n73), .B(a[6]), .C(n75), .D(a[5]), .E(n81), .F(a[4]), 
        .Y(n1366) );
  oa21d1_hd U2024 ( .A(n2012), .B(n49), .C(n1513), .Y(n1487) );
  ao222d1_hd U2025 ( .A(n43), .B(a[15]), .C(n45), .D(a[14]), .E(n51), .F(a[13]), .Y(n1513) );
  ao222d1_hd U2026 ( .A(n73), .B(a[5]), .C(n75), .D(a[4]), .E(n81), .F(a[3]), 
        .Y(n1367) );
  ao222d1_hd U2027 ( .A(n63), .B(a[9]), .C(n65), .D(a[8]), .E(n71), .F(a[7]), 
        .Y(n1415) );
  ao222d1_hd U2028 ( .A(n73), .B(a[3]), .C(n75), .D(a[2]), .E(n81), .F(a[1]), 
        .Y(n1369) );
  ao222d1_hd U2029 ( .A(n63), .B(a[6]), .C(n65), .D(a[5]), .E(n71), .F(a[4]), 
        .Y(n1418) );
  ao222d1_hd U2030 ( .A(n53), .B(a[7]), .C(n55), .D(a[6]), .E(n61), .F(a[5]), 
        .Y(n1469) );
  had1_hd U2031 ( .A(b[23]), .B(n1131), .CO(n711), .S(n712) );
  xo2d1_hd U2032 ( .A(b[23]), .B(n1346), .Y(n1131) );
  oa21d1_hd U2033 ( .A(n79), .B(n1762), .C(n1975), .Y(n1346) );
  ivd1_hd U2034 ( .A(n1014), .Y(n1016) );
  ivd1_hd U2035 ( .A(n1013), .Y(n1015) );
  ao21d1_hd U2036 ( .A(n1016), .B(n988), .C(n989), .Y(n987) );
  oa21d1_hd U2037 ( .A(n1000), .B(n990), .C(n993), .Y(n989) );
  ivd1_hd U2038 ( .A(n998), .Y(n1000) );
  clknd2d1_hd U2039 ( .A(n988), .B(n1015), .Y(n986) );
  ao21d1_hd U2040 ( .A(n1016), .B(n997), .C(n998), .Y(n996) );
  clknd2d1_hd U2041 ( .A(n1015), .B(n997), .Y(n995) );
  nr2d1_hd U2042 ( .A(a[11]), .B(a[10]), .Y(n1028) );
  xn2d1_hd U2043 ( .A(b[9]), .B(b[10]), .Y(n1825) );
  nr2d1_hd U2044 ( .A(a[12]), .B(a[13]), .Y(n1010) );
  nr2d1_hd U2045 ( .A(n1028), .B(n1021), .Y(n1019) );
  oa21d1_hd U2046 ( .A(n1003), .B(n1011), .C(n1004), .Y(n998) );
  clknd2d1_hd U2047 ( .A(a[14]), .B(a[15]), .Y(n993) );
  nr2d1_hd U2048 ( .A(a[15]), .B(a[16]), .Y(n983) );
  clknd2d1_hd U2049 ( .A(a[15]), .B(a[16]), .Y(n984) );
  nr2d1_hd U2050 ( .A(n1050), .B(n1053), .Y(n1048) );
  nr2d1_hd U2051 ( .A(a[18]), .B(a[19]), .Y(n960) );
  ivd1_hd U2052 ( .A(n933), .Y(n931) );
  clknd2d1_hd U2053 ( .A(n61), .B(a[23]), .Y(n1451) );
  ad2d1_hd U2054 ( .A(b[23]), .B(a[12]), .Y(n850) );
  ad2d1_hd U2055 ( .A(b[23]), .B(a[15]), .Y(n847) );
  ivd1_hd U2056 ( .A(n850), .Y(n516) );
  clknd2d1_hd U2057 ( .A(n51), .B(a[23]), .Y(n1503) );
  clknd2d1_hd U2058 ( .A(n41), .B(a[23]), .Y(n1555) );
  xn2d1_hd U2059 ( .A(b[15]), .B(b[16]), .Y(n1823) );
  ao222d1_hd U2060 ( .A(n63), .B(a[17]), .C(n65), .D(a[16]), .E(n71), .F(a[15]), .Y(n1407) );
  fad1_hd U2061 ( .A(n851), .B(n1213), .CI(n853), .CO(n525), .S(n526) );
  ivd1_hd U2062 ( .A(b[11]), .Y(n1213) );
  ad2d1_hd U2063 ( .A(b[23]), .B(a[11]), .Y(n851) );
  oa21d1_hd U2064 ( .A(n2011), .B(n79), .C(n1358), .Y(n1332) );
  ao222d1_hd U2065 ( .A(n73), .B(a[14]), .C(n75), .D(a[13]), .E(n81), .F(a[12]), .Y(n1358) );
  ivd1_hd U2066 ( .A(n853), .Y(n548) );
  oa21d1_hd U2067 ( .A(n2013), .B(n69), .C(n1408), .Y(n1382) );
  ao222d1_hd U2068 ( .A(n63), .B(a[16]), .C(n65), .D(a[15]), .E(n71), .F(a[14]), .Y(n1408) );
  oa21d1_hd U2069 ( .A(n2010), .B(n79), .C(n1359), .Y(n1333) );
  ao222d1_hd U2070 ( .A(n73), .B(a[13]), .C(n75), .D(a[12]), .E(n81), .F(a[11]), .Y(n1359) );
  ao222d1_hd U2071 ( .A(n53), .B(a[17]), .C(n55), .D(a[16]), .E(n61), .F(a[15]), .Y(n1459) );
  oa21d1_hd U2072 ( .A(n2011), .B(n69), .C(n1410), .Y(n1384) );
  ao222d1_hd U2073 ( .A(n63), .B(a[14]), .C(n65), .D(a[13]), .E(n71), .F(a[12]), .Y(n1410) );
  fad1_hd U2074 ( .A(n855), .B(n1240), .CI(n854), .CO(n559), .S(n560) );
  ivd1_hd U2075 ( .A(b[8]), .Y(n1240) );
  ad2d1_hd U2076 ( .A(b[23]), .B(a[8]), .Y(n854) );
  oa21d1_hd U2077 ( .A(n2014), .B(n59), .C(n1458), .Y(n1432) );
  ao222d1_hd U2078 ( .A(n53), .B(a[18]), .C(n55), .D(a[17]), .E(n61), .F(a[16]), .Y(n1458) );
  oa21d1_hd U2079 ( .A(n2020), .B(n39), .C(n1556), .Y(n1530) );
  ao21d1_hd U2080 ( .A(n41), .B(a[22]), .C(n875), .Y(n1556) );
  ad2d1_hd U2081 ( .A(n35), .B(a[23]), .Y(n875) );
  oa21d1_hd U2082 ( .A(n2012), .B(n69), .C(n1409), .Y(n1383) );
  ao222d1_hd U2083 ( .A(n63), .B(a[15]), .C(n65), .D(a[14]), .E(n71), .F(a[13]), .Y(n1409) );
  ao222d1_hd U2084 ( .A(n73), .B(a[10]), .C(n75), .D(a[9]), .E(n81), .F(a[8]), 
        .Y(n1362) );
  oa21d1_hd U2085 ( .A(n2010), .B(n69), .C(n1411), .Y(n1385) );
  ao222d1_hd U2086 ( .A(n63), .B(a[13]), .C(n65), .D(a[12]), .E(n71), .F(a[11]), .Y(n1411) );
  ad2d1_hd U2087 ( .A(b[23]), .B(a[6]), .Y(n856) );
  clknd2d1_hd U2088 ( .A(n31), .B(a[23]), .Y(n1607) );
  ad2d1_hd U2089 ( .A(b[23]), .B(a[7]), .Y(n855) );
  ao222d1_hd U2090 ( .A(n73), .B(a[11]), .C(n75), .D(a[10]), .E(n81), .F(a[9]), 
        .Y(n1361) );
  oa21d1_hd U2091 ( .A(n2019), .B(n39), .C(n1557), .Y(n1531) );
  ao222d1_hd U2092 ( .A(n33), .B(a[23]), .C(n35), .D(a[22]), .E(n41), .F(a[21]), .Y(n1557) );
  ao222d1_hd U2093 ( .A(n43), .B(a[17]), .C(n45), .D(a[16]), .E(n51), .F(a[15]), .Y(n1511) );
  oa21d1_hd U2094 ( .A(n2011), .B(n59), .C(n1462), .Y(n1436) );
  ao222d1_hd U2095 ( .A(n53), .B(a[14]), .C(n55), .D(a[13]), .E(n61), .F(a[12]), .Y(n1462) );
  fad1_hd U2096 ( .A(n1294), .B(n1267), .CI(n857), .CO(n599), .S(n600) );
  ad2d1_hd U2097 ( .A(b[23]), .B(a[5]), .Y(n857) );
  ivd1_hd U2098 ( .A(b[2]), .Y(n1294) );
  ivd1_hd U2099 ( .A(b[5]), .Y(n1267) );
  ao222d1_hd U2100 ( .A(n63), .B(a[12]), .C(n65), .D(a[11]), .E(n71), .F(a[10]), .Y(n1412) );
  oa21d1_hd U2101 ( .A(n2012), .B(n59), .C(n1461), .Y(n1435) );
  ao222d1_hd U2102 ( .A(n53), .B(a[15]), .C(n55), .D(a[14]), .E(n61), .F(a[13]), .Y(n1461) );
  oa21d1_hd U2103 ( .A(n2013), .B(n59), .C(n1460), .Y(n1434) );
  ao222d1_hd U2104 ( .A(n53), .B(a[16]), .C(n55), .D(a[15]), .E(n61), .F(a[14]), .Y(n1460) );
  oa21d1_hd U2105 ( .A(n2015), .B(n49), .C(n1509), .Y(n1483) );
  ao222d1_hd U2106 ( .A(n43), .B(a[19]), .C(n45), .D(a[18]), .E(n51), .F(a[17]), .Y(n1509) );
  oa21d1_hd U2107 ( .A(n2014), .B(n49), .C(n1510), .Y(n1484) );
  ao222d1_hd U2108 ( .A(n43), .B(a[18]), .C(n45), .D(a[17]), .E(n51), .F(a[16]), .Y(n1510) );
  oa21d1_hd U2109 ( .A(n2017), .B(n39), .C(n1559), .Y(n1533) );
  ao222d1_hd U2110 ( .A(n33), .B(a[21]), .C(n35), .D(a[20]), .E(n41), .F(a[19]), .Y(n1559) );
  oa21d1_hd U2111 ( .A(n2020), .B(n29), .C(n1608), .Y(n1582) );
  ao21d1_hd U2112 ( .A(n31), .B(a[22]), .C(n878), .Y(n1608) );
  ad2d1_hd U2113 ( .A(n25), .B(a[23]), .Y(n878) );
  ao222d1_hd U2114 ( .A(n73), .B(a[8]), .C(n75), .D(a[7]), .E(n81), .F(a[6]), 
        .Y(n1364) );
  oa21d1_hd U2115 ( .A(n2008), .B(n69), .C(n1413), .Y(n1387) );
  ao222d1_hd U2116 ( .A(n63), .B(a[11]), .C(n65), .D(a[10]), .E(n71), .F(a[9]), 
        .Y(n1413) );
  oa21d1_hd U2117 ( .A(n2010), .B(n59), .C(n1463), .Y(n1437) );
  ao222d1_hd U2118 ( .A(n53), .B(a[13]), .C(n55), .D(a[12]), .E(n61), .F(a[11]), .Y(n1463) );
  oa21d1_hd U2119 ( .A(n2013), .B(n49), .C(n1512), .Y(n1486) );
  ao222d1_hd U2120 ( .A(n43), .B(a[16]), .C(n45), .D(a[15]), .E(n51), .F(a[14]), .Y(n1512) );
  ao222d1_hd U2121 ( .A(n33), .B(a[20]), .C(n35), .D(a[19]), .E(n41), .F(a[18]), .Y(n1560) );
  oa21d1_hd U2122 ( .A(n2019), .B(n29), .C(n1609), .Y(n1583) );
  ao222d1_hd U2123 ( .A(n23), .B(a[23]), .C(n25), .D(a[22]), .E(n31), .F(a[21]), .Y(n1609) );
  ao222d1_hd U2124 ( .A(n33), .B(a[19]), .C(n35), .D(a[18]), .E(n41), .F(a[17]), .Y(n1561) );
  ao222d1_hd U2125 ( .A(n23), .B(a[21]), .C(n25), .D(a[20]), .E(n31), .F(a[19]), .Y(n1611) );
  oa21d1_hd U2126 ( .A(n2020), .B(n19), .C(n1660), .Y(n1634) );
  ao21d1_hd U2127 ( .A(n21), .B(a[22]), .C(n881), .Y(n1660) );
  ad2d1_hd U2128 ( .A(n15), .B(a[23]), .Y(n881) );
  fad1_hd U2129 ( .A(n641), .B(n1125), .CI(n1197), .CO(n625), .S(n626) );
  xo2d1_hd U2130 ( .A(b[23]), .B(n1340), .Y(n1125) );
  xo2d1_hd U2131 ( .A(b[14]), .B(n1487), .Y(n1197) );
  oa21d1_hd U2132 ( .A(n2003), .B(n79), .C(n1366), .Y(n1340) );
  oa21d1_hd U2133 ( .A(n2008), .B(n59), .C(n1465), .Y(n1439) );
  ao222d1_hd U2134 ( .A(n53), .B(a[11]), .C(n55), .D(a[10]), .E(n61), .F(a[9]), 
        .Y(n1465) );
  oa21d1_hd U2135 ( .A(n2011), .B(n49), .C(n1514), .Y(n1488) );
  ao222d1_hd U2136 ( .A(n43), .B(a[14]), .C(n45), .D(a[13]), .E(n51), .F(a[12]), .Y(n1514) );
  oa21d1_hd U2137 ( .A(n1998), .B(n39), .C(n1563), .Y(n1537) );
  ao222d1_hd U2138 ( .A(n33), .B(a[17]), .C(n35), .D(a[16]), .E(n41), .F(a[15]), .Y(n1563) );
  fad1_hd U2139 ( .A(n860), .B(b[2]), .CI(n1126), .CO(n641), .S(n642) );
  ad2d1_hd U2140 ( .A(b[23]), .B(a[2]), .Y(n860) );
  xo2d1_hd U2141 ( .A(b[23]), .B(n1341), .Y(n1126) );
  oa21d1_hd U2142 ( .A(n2002), .B(n79), .C(n1367), .Y(n1341) );
  ao222d1_hd U2143 ( .A(n33), .B(a[18]), .C(n35), .D(a[17]), .E(n41), .F(a[16]), .Y(n1562) );
  clknd2d1_hd U2144 ( .A(n11), .B(a[23]), .Y(n1711) );
  oa21d1_hd U2145 ( .A(n2013), .B(n39), .C(n1564), .Y(n1538) );
  ao222d1_hd U2146 ( .A(n33), .B(a[16]), .C(n35), .D(a[15]), .E(n41), .F(a[14]), .Y(n1564) );
  fad1_hd U2147 ( .A(n1128), .B(n862), .CI(n683), .CO(n669), .S(n670) );
  ad2d1_hd U2148 ( .A(b[23]), .B(a[0]), .Y(n862) );
  xo2d1_hd U2149 ( .A(b[23]), .B(n1343), .Y(n1128) );
  oa21d1_hd U2150 ( .A(n2000), .B(n79), .C(n1369), .Y(n1343) );
  ao222d1_hd U2151 ( .A(n53), .B(a[10]), .C(n55), .D(a[9]), .E(n61), .F(a[8]), 
        .Y(n1466) );
  oa21d1_hd U2152 ( .A(n2010), .B(n49), .C(n1515), .Y(n1489) );
  ao222d1_hd U2153 ( .A(n43), .B(a[13]), .C(n45), .D(a[12]), .E(n51), .F(a[11]), .Y(n1515) );
  fad1_hd U2154 ( .A(n1127), .B(n861), .CI(n1151), .CO(n655), .S(n656) );
  ad2d1_hd U2155 ( .A(b[23]), .B(a[1]), .Y(n861) );
  xo2d1_hd U2156 ( .A(b[20]), .B(n1391), .Y(n1151) );
  xo2d1_hd U2157 ( .A(b[23]), .B(n1342), .Y(n1127) );
  ao222d1_hd U2158 ( .A(n23), .B(a[20]), .C(n25), .D(a[19]), .E(n31), .F(a[18]), .Y(n1612) );
  oa21d1_hd U2159 ( .A(n2019), .B(n19), .C(n1661), .Y(n1635) );
  ao222d1_hd U2160 ( .A(n13), .B(a[23]), .C(n15), .D(a[22]), .E(n21), .F(a[21]), .Y(n1661) );
  ao222d1_hd U2161 ( .A(n23), .B(a[19]), .C(n25), .D(a[18]), .E(n31), .F(a[17]), .Y(n1613) );
  ao222d1_hd U2162 ( .A(n13), .B(a[21]), .C(n15), .D(a[20]), .E(n21), .F(a[19]), .Y(n1663) );
  oa21d1_hd U2163 ( .A(n2020), .B(n9), .C(n1712), .Y(n1686) );
  ao21d1_hd U2164 ( .A(n11), .B(a[22]), .C(n884), .Y(n1712) );
  ad2d1_hd U2165 ( .A(n5), .B(a[23]), .Y(n884) );
  fad1_hd U2166 ( .A(n1152), .B(n1176), .CI(n670), .CO(n667), .S(n668) );
  xo2d1_hd U2167 ( .A(b[20]), .B(n1392), .Y(n1152) );
  xo2d1_hd U2168 ( .A(b[17]), .B(n1441), .Y(n1176) );
  oa21d1_hd U2169 ( .A(n2003), .B(n69), .C(n1418), .Y(n1392) );
  oa21d1_hd U2170 ( .A(n2012), .B(n39), .C(n1565), .Y(n1539) );
  ao222d1_hd U2171 ( .A(n33), .B(a[15]), .C(n35), .D(a[14]), .E(n41), .F(a[13]), .Y(n1565) );
  oa21d1_hd U2172 ( .A(n2014), .B(n29), .C(n1614), .Y(n1588) );
  ao222d1_hd U2173 ( .A(n23), .B(a[18]), .C(n25), .D(a[17]), .E(n31), .F(a[16]), .Y(n1614) );
  ao222d1_hd U2174 ( .A(n53), .B(a[8]), .C(n55), .D(a[7]), .E(n61), .F(a[6]), 
        .Y(n1468) );
  oa21d1_hd U2175 ( .A(n2008), .B(n49), .C(n1517), .Y(n1491) );
  ao222d1_hd U2176 ( .A(n43), .B(a[11]), .C(n45), .D(a[10]), .E(n51), .F(a[9]), 
        .Y(n1517) );
  had1_hd U2177 ( .A(n1129), .B(n697), .CO(n683), .S(n684) );
  xo2d1_hd U2178 ( .A(b[23]), .B(n1344), .Y(n1129) );
  oa21d1_hd U2179 ( .A(n1999), .B(n79), .C(n1370), .Y(n1344) );
  ao222d1_hd U2180 ( .A(n73), .B(a[2]), .C(n75), .D(a[1]), .E(n81), .F(a[0]), 
        .Y(n1370) );
  ao222d1_hd U2181 ( .A(n23), .B(a[17]), .C(n25), .D(a[16]), .E(n31), .F(a[15]), .Y(n1615) );
  oa21d1_hd U2182 ( .A(n2002), .B(n69), .C(n1419), .Y(n1393) );
  ao222d1_hd U2183 ( .A(n63), .B(a[5]), .C(n65), .D(a[4]), .E(n71), .F(a[3]), 
        .Y(n1419) );
  oa21d1_hd U2184 ( .A(n2019), .B(n9), .C(n1713), .Y(n1687) );
  ao222d1_hd U2185 ( .A(n3), .B(a[23]), .C(n5), .D(a[22]), .E(n11), .F(a[21]), 
        .Y(n1713) );
  oa21d1_hd U2186 ( .A(n2011), .B(n39), .C(n1566), .Y(n1540) );
  ao222d1_hd U2187 ( .A(n33), .B(a[14]), .C(n35), .D(a[13]), .E(n41), .F(a[12]), .Y(n1566) );
  oa21d1_hd U2188 ( .A(n2016), .B(n19), .C(n1664), .Y(n1638) );
  ao222d1_hd U2189 ( .A(n13), .B(a[20]), .C(n15), .D(a[19]), .E(n21), .F(a[18]), .Y(n1664) );
  ao222d1_hd U2190 ( .A(n3), .B(a[22]), .C(n5), .D(a[21]), .E(n11), .F(a[20]), 
        .Y(n1714) );
  oa21d1_hd U2191 ( .A(n2010), .B(n39), .C(n1567), .Y(n1541) );
  ao222d1_hd U2192 ( .A(n33), .B(a[13]), .C(n35), .D(a[12]), .E(n41), .F(a[11]), .Y(n1567) );
  ao222d1_hd U2193 ( .A(n43), .B(a[10]), .C(n45), .D(a[9]), .E(n51), .F(a[8]), 
        .Y(n1518) );
  oa21d1_hd U2194 ( .A(n2013), .B(n29), .C(n1616), .Y(n1590) );
  ao222d1_hd U2195 ( .A(n23), .B(a[16]), .C(n25), .D(a[15]), .E(n31), .F(a[14]), .Y(n1616) );
  ao222d1_hd U2196 ( .A(n53), .B(a[6]), .C(n55), .D(a[5]), .E(n61), .F(a[4]), 
        .Y(n1470) );
  fad1_hd U2197 ( .A(n1155), .B(n712), .CI(n723), .CO(n709), .S(n710) );
  xo2d1_hd U2198 ( .A(b[20]), .B(n1395), .Y(n1155) );
  oa21d1_hd U2199 ( .A(n2000), .B(n69), .C(n1421), .Y(n1395) );
  ao222d1_hd U2200 ( .A(n63), .B(a[3]), .C(n65), .D(a[2]), .E(n71), .F(a[1]), 
        .Y(n1421) );
  nr2d1_hd U2201 ( .A(a[17]), .B(a[18]), .Y(n971) );
  nr2d1_hd U2202 ( .A(a[17]), .B(a[16]), .Y(n974) );
  clknd2d1_hd U2203 ( .A(a[17]), .B(a[16]), .Y(n975) );
  clknd2d1_hd U2204 ( .A(a[17]), .B(a[18]), .Y(n972) );
  oa21d1_hd U2205 ( .A(n2012), .B(n29), .C(n1617), .Y(n1591) );
  ao222d1_hd U2206 ( .A(n23), .B(a[15]), .C(n25), .D(a[14]), .E(n31), .F(a[13]), .Y(n1617) );
  oa21d1_hd U2207 ( .A(n2017), .B(n9), .C(n1715), .Y(n1689) );
  ao222d1_hd U2208 ( .A(n3), .B(a[21]), .C(n5), .D(a[20]), .E(n11), .F(a[19]), 
        .Y(n1715) );
  ao222d1_hd U2209 ( .A(n13), .B(a[17]), .C(n15), .D(a[16]), .E(n21), .F(a[15]), .Y(n1667) );
  oa21d1_hd U2210 ( .A(n2002), .B(n59), .C(n1471), .Y(n1445) );
  ao222d1_hd U2211 ( .A(n53), .B(a[5]), .C(n55), .D(a[4]), .E(n61), .F(a[3]), 
        .Y(n1471) );
  nr2d1_hd U2212 ( .A(a[14]), .B(a[13]), .Y(n1003) );
  ao21d1_hd U2213 ( .A(n1016), .B(n1092), .C(n1009), .Y(n1007) );
  ivd1_hd U2214 ( .A(n1011), .Y(n1009) );
  clknd2d1_hd U2215 ( .A(n1015), .B(n1092), .Y(n1006) );
  clknd2d1_hd U2216 ( .A(a[14]), .B(a[13]), .Y(n1004) );
  ao222d1_hd U2217 ( .A(n43), .B(a[8]), .C(n45), .D(a[7]), .E(n51), .F(a[6]), 
        .Y(n1520) );
  oa21d1_hd U2218 ( .A(n2008), .B(n39), .C(n1569), .Y(n1543) );
  ao222d1_hd U2219 ( .A(n33), .B(a[11]), .C(n35), .D(a[10]), .E(n41), .F(a[9]), 
        .Y(n1569) );
  had1_hd U2220 ( .A(n747), .B(n1157), .CO(n735), .S(n736) );
  xo2d1_hd U2221 ( .A(b[20]), .B(n1397), .Y(n1157) );
  oa21d1_hd U2222 ( .A(n69), .B(n1761), .C(n1990), .Y(n1397) );
  ao222d1_hd U2223 ( .A(n43), .B(a[7]), .C(n45), .D(a[6]), .E(n51), .F(a[5]), 
        .Y(n1521) );
  ivd1_hd U2224 ( .A(n960), .Y(n958) );
  ivd1_hd U2225 ( .A(n965), .Y(n963) );
  ao222d1_hd U2226 ( .A(n13), .B(a[16]), .C(n15), .D(a[15]), .E(n21), .F(a[14]), .Y(n1668) );
  oa21d1_hd U2227 ( .A(n2010), .B(n29), .C(n1619), .Y(n1593) );
  ao222d1_hd U2228 ( .A(n23), .B(a[13]), .C(n25), .D(a[12]), .E(n31), .F(a[11]), .Y(n1619) );
  ao222d1_hd U2229 ( .A(n43), .B(a[6]), .C(n45), .D(a[5]), .E(n51), .F(a[4]), 
        .Y(n1522) );
  fad1_hd U2230 ( .A(n1182), .B(n748), .CI(n757), .CO(n745), .S(n746) );
  xo2d1_hd U2231 ( .A(b[17]), .B(n1447), .Y(n1182) );
  oa21d1_hd U2232 ( .A(n2000), .B(n59), .C(n1473), .Y(n1447) );
  ao222d1_hd U2233 ( .A(n53), .B(a[3]), .C(n55), .D(a[2]), .E(n61), .F(a[1]), 
        .Y(n1473) );
  oa21d1_hd U2234 ( .A(n2014), .B(n9), .C(n1718), .Y(n1692) );
  ao222d1_hd U2235 ( .A(n3), .B(a[18]), .C(n5), .D(a[17]), .E(n11), .F(a[16]), 
        .Y(n1718) );
  oa21d1_hd U2236 ( .A(n2012), .B(n19), .C(n1669), .Y(n1643) );
  ao222d1_hd U2237 ( .A(n13), .B(a[15]), .C(n15), .D(a[14]), .E(n21), .F(a[13]), .Y(n1669) );
  ao222d1_hd U2238 ( .A(n3), .B(a[17]), .C(n5), .D(a[16]), .E(n11), .F(a[15]), 
        .Y(n1719) );
  had1_hd U2239 ( .A(n1183), .B(n767), .CO(n757), .S(n758) );
  xo2d1_hd U2240 ( .A(b[17]), .B(n1448), .Y(n1183) );
  oa21d1_hd U2241 ( .A(n1999), .B(n59), .C(n1474), .Y(n1448) );
  ao222d1_hd U2242 ( .A(n53), .B(a[2]), .C(n55), .D(a[1]), .E(n61), .F(a[0]), 
        .Y(n1474) );
  oa21d1_hd U2243 ( .A(n2002), .B(n49), .C(n1523), .Y(n1497) );
  ao222d1_hd U2244 ( .A(n43), .B(a[5]), .C(n45), .D(a[4]), .E(n51), .F(a[3]), 
        .Y(n1523) );
  xn2d1_hd U2245 ( .A(n893), .B(n1), .Y(n1998) );
  clknd2d1_hd U2246 ( .A(n1088), .B(n975), .Y(n893) );
  ivd1_hd U2247 ( .A(n974), .Y(n1088) );
  ivd1_hd U2248 ( .A(n1033), .Y(n1031) );
  clknd2d1_hd U2249 ( .A(n1089), .B(n984), .Y(n894) );
  oa21d1_hd U2250 ( .A(n1044), .B(n986), .C(n987), .Y(n985) );
  ivd1_hd U2251 ( .A(n983), .Y(n1089) );
  ao222d1_hd U2252 ( .A(n33), .B(a[7]), .C(n35), .D(a[6]), .E(n41), .F(a[5]), 
        .Y(n1573) );
  clknd2d1_hd U2253 ( .A(a[12]), .B(a[13]), .Y(n1011) );
  ivd1_hd U2254 ( .A(n1010), .Y(n1092) );
  had1_hd U2255 ( .A(b[17]), .B(n1185), .CO(n777), .S(n778) );
  xo2d1_hd U2256 ( .A(b[17]), .B(n1450), .Y(n1185) );
  oa21d1_hd U2257 ( .A(n59), .B(n1762), .C(n1996), .Y(n1450) );
  clknd2d1_hd U2259 ( .A(n1090), .B(n993), .Y(n895) );
  oa21d1_hd U2260 ( .A(n1044), .B(n995), .C(n996), .Y(n994) );
  ivd1_hd U2261 ( .A(n990), .Y(n1090) );
  clknd2d1_hd U2262 ( .A(a[11]), .B(a[10]), .Y(n1029) );
  ad3d2_hd U2263 ( .A(n1833), .B(n1825), .C(n1817), .Y(n41) );
  xn2d1_hd U2264 ( .A(b[6]), .B(b[7]), .Y(n1826) );
  ao21d1_hd U2265 ( .A(n1075), .B(n1067), .C(n1068), .Y(n1066) );
  nr2d1_hd U2266 ( .A(n1072), .B(n1069), .Y(n1067) );
  oa21d1_hd U2267 ( .A(n1073), .B(n1069), .C(n1070), .Y(n1068) );
  nr2d1_hd U2268 ( .A(a[5]), .B(a[4]), .Y(n1063) );
  clknd2d1_hd U2269 ( .A(n1019), .B(n1033), .Y(n1013) );
  nr2d1_hd U2271 ( .A(n990), .B(n983), .Y(n981) );
  ao21d1_hd U2272 ( .A(n1019), .B(n1034), .C(n1020), .Y(n1014) );
  oa21d1_hd U2273 ( .A(n1021), .B(n1029), .C(n1022), .Y(n1020) );
  ao21d1_hd U2274 ( .A(n998), .B(n981), .C(n982), .Y(n980) );
  oa21d1_hd U2275 ( .A(n993), .B(n983), .C(n984), .Y(n982) );
  clknd2d1_hd U2276 ( .A(a[18]), .B(a[19]), .Y(n961) );
  ivd1_hd U2277 ( .A(n925), .Y(n923) );
  nr2d1_hd U2278 ( .A(n945), .B(n931), .Y(n929) );
  ivd1_hd U2279 ( .A(n929), .Y(n927) );
  clknd2d1_hd U2280 ( .A(a[23]), .B(a[22]), .Y(n925) );
  oa21d1_hd U2281 ( .A(n946), .B(n931), .C(n932), .Y(n930) );
  ivd1_hd U2282 ( .A(n934), .Y(n932) );
  ivd1_hd U2283 ( .A(n924), .Y(n922) );
  ad2d1_hd U2284 ( .A(b[23]), .B(a[18]), .Y(n844) );
  clknd2d1_hd U2285 ( .A(n71), .B(a[23]), .Y(n1399) );
  clknd2d1_hd U2286 ( .A(a[20]), .B(a[21]), .Y(n943) );
  ad2d1_hd U2287 ( .A(n65), .B(a[23]), .Y(n866) );
  ivd1_hd U2288 ( .A(n844), .Y(n470) );
  nr2d1_hd U2289 ( .A(a[20]), .B(a[19]), .Y(n953) );
  ao21d1_hd U2290 ( .A(n966), .B(n958), .C(n959), .Y(n957) );
  ivd1_hd U2291 ( .A(n961), .Y(n959) );
  clknd2d1_hd U2292 ( .A(n965), .B(n958), .Y(n956) );
  clknd2d1_hd U2293 ( .A(a[20]), .B(a[19]), .Y(n954) );
  ad3d2_hd U2295 ( .A(n1830), .B(n1822), .C(n1814), .Y(n71) );
  fad1_hd U2296 ( .A(n847), .B(n1159), .CI(n845), .CO(n475), .S(n476) );
  ivd1_hd U2297 ( .A(b[17]), .Y(n1159) );
  ad2d1_hd U2298 ( .A(b[23]), .B(a[17]), .Y(n845) );
  xn2d1_hd U2299 ( .A(b[21]), .B(b[22]), .Y(n1821) );
  ao222d1_hd U2300 ( .A(n73), .B(a[19]), .C(n75), .D(a[18]), .E(n81), .F(a[17]), .Y(n1353) );
  fad1_hd U2301 ( .A(n490), .B(n846), .CI(n1160), .CO(n481), .S(n482) );
  ad2d1_hd U2302 ( .A(b[23]), .B(a[16]), .Y(n846) );
  xo2d1_hd U2303 ( .A(b[17]), .B(n1425), .Y(n1160) );
  oa21d1_hd U2304 ( .A(n1970), .B(n59), .C(n1451), .Y(n1425) );
  fad1_hd U2305 ( .A(n850), .B(n1186), .CI(n848), .CO(n497), .S(n498) );
  ivd1_hd U2306 ( .A(b[14]), .Y(n1186) );
  ad2d1_hd U2307 ( .A(b[23]), .B(a[14]), .Y(n848) );
  ad2d1_hd U2308 ( .A(n55), .B(a[23]), .Y(n869) );
  ivd1_hd U2309 ( .A(n847), .Y(n490) );
  ao222d1_hd U2310 ( .A(n73), .B(a[18]), .C(n75), .D(a[17]), .E(n81), .F(a[16]), .Y(n1354) );
  oa21d1_hd U2311 ( .A(n2017), .B(n69), .C(n1403), .Y(n1377) );
  ao222d1_hd U2312 ( .A(n63), .B(a[21]), .C(n65), .D(a[20]), .E(n71), .F(a[19]), .Y(n1403) );
  oa21d1_hd U2313 ( .A(n2013), .B(n79), .C(n1356), .Y(n1330) );
  ao222d1_hd U2314 ( .A(n73), .B(a[16]), .C(n75), .D(a[15]), .E(n81), .F(a[14]), .Y(n1356) );
  oa21d1_hd U2315 ( .A(n2015), .B(n69), .C(n1405), .Y(n1379) );
  ao222d1_hd U2316 ( .A(n63), .B(a[19]), .C(n65), .D(a[18]), .E(n71), .F(a[17]), .Y(n1405) );
  ao222d1_hd U2317 ( .A(n63), .B(a[20]), .C(n65), .D(a[19]), .E(n71), .F(a[18]), .Y(n1404) );
  oa21d1_hd U2318 ( .A(n2019), .B(n59), .C(n1453), .Y(n1427) );
  ao222d1_hd U2319 ( .A(n53), .B(a[23]), .C(n55), .D(a[22]), .E(n61), .F(a[21]), .Y(n1453) );
  fad1_hd U2320 ( .A(n1114), .B(n498), .CI(n505), .CO(n495), .S(n496) );
  xo2d1_hd U2321 ( .A(b[23]), .B(n1329), .Y(n1114) );
  oa21d1_hd U2322 ( .A(n1998), .B(n79), .C(n1355), .Y(n1329) );
  ao222d1_hd U2323 ( .A(n73), .B(a[17]), .C(n75), .D(a[16]), .E(n81), .F(a[15]), .Y(n1355) );
  ao222d1_hd U2324 ( .A(n53), .B(a[21]), .C(n55), .D(a[20]), .E(n61), .F(a[19]), .Y(n1455) );
  oa21d1_hd U2325 ( .A(n2014), .B(n69), .C(n1406), .Y(n1380) );
  ao222d1_hd U2326 ( .A(n63), .B(a[18]), .C(n65), .D(a[17]), .E(n71), .F(a[16]), .Y(n1406) );
  fad1_hd U2327 ( .A(n525), .B(n516), .CI(n1116), .CO(n514), .S(n515) );
  xo2d1_hd U2328 ( .A(b[23]), .B(n1331), .Y(n1116) );
  oa21d1_hd U2329 ( .A(n2012), .B(n79), .C(n1357), .Y(n1331) );
  ao222d1_hd U2330 ( .A(n73), .B(a[15]), .C(n75), .D(a[14]), .E(n81), .F(a[13]), .Y(n1357) );
  ao222d1_hd U2331 ( .A(n43), .B(a[23]), .C(n45), .D(a[22]), .E(n51), .F(a[21]), .Y(n1505) );
  oa21d1_hd U2332 ( .A(n2016), .B(n59), .C(n1456), .Y(n1430) );
  ao222d1_hd U2333 ( .A(n53), .B(a[20]), .C(n55), .D(a[19]), .E(n61), .F(a[18]), .Y(n1456) );
  ad2d1_hd U2334 ( .A(n45), .B(a[23]), .Y(n872) );
  ad3d2_hd U2337 ( .A(n1831), .B(n1815), .C(n1823), .Y(n61) );
  fad1_hd U2338 ( .A(n1141), .B(n526), .CI(n1117), .CO(n523), .S(n524) );
  xo2d1_hd U2339 ( .A(b[20]), .B(n1381), .Y(n1141) );
  xo2d1_hd U2340 ( .A(b[23]), .B(n1332), .Y(n1117) );
  oa21d1_hd U2341 ( .A(n1998), .B(n69), .C(n1407), .Y(n1381) );
  fad1_hd U2342 ( .A(n1118), .B(n1142), .CI(n1190), .CO(n533), .S(n534) );
  xo2d1_hd U2343 ( .A(b[23]), .B(n1333), .Y(n1118) );
  xo2d1_hd U2344 ( .A(b[14]), .B(n1480), .Y(n1190) );
  xo2d1_hd U2345 ( .A(b[20]), .B(n1382), .Y(n1142) );
  fad1_hd U2346 ( .A(n1168), .B(n560), .CI(n1144), .CO(n557), .S(n558) );
  xo2d1_hd U2347 ( .A(b[17]), .B(n1433), .Y(n1168) );
  xo2d1_hd U2348 ( .A(b[20]), .B(n1384), .Y(n1144) );
  oa21d1_hd U2349 ( .A(n1998), .B(n59), .C(n1459), .Y(n1433) );
  ad3d2_hd U2350 ( .A(n1832), .B(n1824), .C(n1816), .Y(n51) );
  fad1_hd U2351 ( .A(n1167), .B(n1143), .CI(n1215), .CO(n544), .S(n545) );
  xo2d1_hd U2352 ( .A(b[20]), .B(n1383), .Y(n1143) );
  xo2d1_hd U2353 ( .A(b[11]), .B(n1530), .Y(n1215) );
  xo2d1_hd U2354 ( .A(b[17]), .B(n1432), .Y(n1167) );
  fad1_hd U2355 ( .A(n571), .B(n1120), .CI(n1216), .CO(n555), .S(n556) );
  xo2d1_hd U2356 ( .A(b[23]), .B(n1335), .Y(n1120) );
  xo2d1_hd U2357 ( .A(b[11]), .B(n1531), .Y(n1216) );
  oa21d1_hd U2358 ( .A(n2008), .B(n79), .C(n1361), .Y(n1335) );
  fad1_hd U2359 ( .A(n1195), .B(n600), .CI(n1171), .CO(n597), .S(n598) );
  xo2d1_hd U2360 ( .A(b[14]), .B(n1485), .Y(n1195) );
  xo2d1_hd U2361 ( .A(b[17]), .B(n1436), .Y(n1171) );
  oa21d1_hd U2362 ( .A(n1998), .B(n49), .C(n1511), .Y(n1485) );
  fad1_hd U2363 ( .A(n1217), .B(n1169), .CI(n1193), .CO(n567), .S(n568) );
  xo2d1_hd U2364 ( .A(b[14]), .B(n1483), .Y(n1193) );
  xo2d1_hd U2365 ( .A(b[17]), .B(n1434), .Y(n1169) );
  xo2d1_hd U2366 ( .A(b[11]), .B(n1532), .Y(n1217) );
  fad1_hd U2367 ( .A(n1218), .B(n1194), .CI(n1242), .CO(n580), .S(n581) );
  xo2d1_hd U2368 ( .A(b[8]), .B(n1582), .Y(n1242) );
  xo2d1_hd U2369 ( .A(b[11]), .B(n1533), .Y(n1218) );
  xo2d1_hd U2370 ( .A(b[14]), .B(n1484), .Y(n1194) );
  fad1_hd U2371 ( .A(n1123), .B(n1147), .CI(n613), .CO(n595), .S(n596) );
  xo2d1_hd U2372 ( .A(b[23]), .B(n1338), .Y(n1123) );
  xo2d1_hd U2373 ( .A(b[20]), .B(n1387), .Y(n1147) );
  oa21d1_hd U2374 ( .A(n2005), .B(n79), .C(n1364), .Y(n1338) );
  fad1_hd U2375 ( .A(n1172), .B(n1268), .CI(n1196), .CO(n611), .S(n612) );
  xo2d1_hd U2376 ( .A(b[5]), .B(n1633), .Y(n1268) );
  xo2d1_hd U2377 ( .A(b[14]), .B(n1486), .Y(n1196) );
  xo2d1_hd U2378 ( .A(b[17]), .B(n1437), .Y(n1172) );
  fad1_hd U2379 ( .A(n1219), .B(n1243), .CI(n598), .CO(n593), .S(n594) );
  xo2d1_hd U2380 ( .A(b[11]), .B(n1534), .Y(n1219) );
  xo2d1_hd U2381 ( .A(b[8]), .B(n1583), .Y(n1243) );
  oa21d1_hd U2382 ( .A(n2016), .B(n39), .C(n1560), .Y(n1534) );
  fad1_hd U2383 ( .A(n1220), .B(n1244), .CI(n625), .CO(n607), .S(n608) );
  xo2d1_hd U2384 ( .A(b[11]), .B(n1535), .Y(n1220) );
  xo2d1_hd U2385 ( .A(b[8]), .B(n1584), .Y(n1244) );
  oa21d1_hd U2386 ( .A(n2015), .B(n39), .C(n1561), .Y(n1535) );
  fad1_hd U2387 ( .A(n1245), .B(n1269), .CI(n626), .CO(n621), .S(n622) );
  xo2d1_hd U2388 ( .A(b[8]), .B(n1585), .Y(n1245) );
  xo2d1_hd U2389 ( .A(b[5]), .B(n1634), .Y(n1269) );
  oa21d1_hd U2390 ( .A(n2017), .B(n29), .C(n1611), .Y(n1585) );
  fad1_hd U2391 ( .A(n1174), .B(n1222), .CI(n1198), .CO(n637), .S(n638) );
  xo2d1_hd U2392 ( .A(b[11]), .B(n1537), .Y(n1222) );
  xo2d1_hd U2393 ( .A(b[14]), .B(n1488), .Y(n1198) );
  xo2d1_hd U2394 ( .A(b[17]), .B(n1439), .Y(n1174) );
  fad1_hd U2395 ( .A(n1150), .B(n642), .CI(n655), .CO(n639), .S(n640) );
  xo2d1_hd U2396 ( .A(b[20]), .B(n1390), .Y(n1150) );
  oa21d1_hd U2397 ( .A(n2005), .B(n69), .C(n1416), .Y(n1390) );
  ao222d1_hd U2398 ( .A(n63), .B(a[8]), .C(n65), .D(a[7]), .E(n71), .F(a[6]), 
        .Y(n1416) );
  fad1_hd U2399 ( .A(n628), .B(n1173), .CI(n1221), .CO(n623), .S(n624) );
  xo2d1_hd U2400 ( .A(b[11]), .B(n1536), .Y(n1221) );
  xo2d1_hd U2401 ( .A(b[17]), .B(n1438), .Y(n1173) );
  oa21d1_hd U2402 ( .A(n2014), .B(n39), .C(n1562), .Y(n1536) );
  fad1_hd U2403 ( .A(n1246), .B(n1270), .CI(n653), .CO(n635), .S(n636) );
  xo2d1_hd U2404 ( .A(b[8]), .B(n1586), .Y(n1246) );
  xo2d1_hd U2405 ( .A(b[5]), .B(n1635), .Y(n1270) );
  oa21d1_hd U2406 ( .A(n2016), .B(n29), .C(n1612), .Y(n1586) );
  fad1_hd U2407 ( .A(n638), .B(n640), .CI(n651), .CO(n633), .S(n634) );
  fad1_hd U2408 ( .A(n1247), .B(n1271), .CI(n667), .CO(n649), .S(n650) );
  xo2d1_hd U2409 ( .A(b[8]), .B(n1587), .Y(n1247) );
  xo2d1_hd U2410 ( .A(b[5]), .B(n1636), .Y(n1271) );
  oa21d1_hd U2411 ( .A(n2015), .B(n29), .C(n1613), .Y(n1587) );
  fad1_hd U2412 ( .A(n1272), .B(n1296), .CI(n668), .CO(n663), .S(n664) );
  xo2d1_hd U2413 ( .A(b[5]), .B(n1637), .Y(n1272) );
  xo2d1_hd U2414 ( .A(b[2]), .B(n1686), .Y(n1296) );
  oa21d1_hd U2415 ( .A(n2017), .B(n19), .C(n1663), .Y(n1637) );
  fad1_hd U2416 ( .A(n1200), .B(n1224), .CI(n1248), .CO(n665), .S(n666) );
  xo2d1_hd U2417 ( .A(b[8]), .B(n1588), .Y(n1248) );
  xo2d1_hd U2418 ( .A(b[14]), .B(n1490), .Y(n1200) );
  xo2d1_hd U2419 ( .A(b[11]), .B(n1539), .Y(n1224) );
  fad1_hd U2420 ( .A(n1177), .B(n1201), .CI(n695), .CO(n679), .S(n680) );
  xo2d1_hd U2421 ( .A(b[17]), .B(n1442), .Y(n1177) );
  xo2d1_hd U2422 ( .A(b[14]), .B(n1491), .Y(n1201) );
  oa21d1_hd U2423 ( .A(n2005), .B(n59), .C(n1468), .Y(n1442) );
  fad1_hd U2424 ( .A(n684), .B(n1153), .CI(n1249), .CO(n681), .S(n682) );
  xo2d1_hd U2425 ( .A(b[8]), .B(n1589), .Y(n1249) );
  xo2d1_hd U2426 ( .A(b[20]), .B(n1393), .Y(n1153) );
  oa21d1_hd U2427 ( .A(n1998), .B(n29), .C(n1615), .Y(n1589) );
  fad1_hd U2428 ( .A(n1297), .B(n1225), .CI(n1273), .CO(n677), .S(n678) );
  xo2d1_hd U2429 ( .A(b[5]), .B(n1638), .Y(n1273) );
  xo2d1_hd U2430 ( .A(b[11]), .B(n1540), .Y(n1225) );
  xo2d1_hd U2431 ( .A(b[2]), .B(n1687), .Y(n1297) );
  fad1_hd U2432 ( .A(n1179), .B(n1203), .CI(n710), .CO(n707), .S(n708) );
  xo2d1_hd U2433 ( .A(b[17]), .B(n1444), .Y(n1179) );
  xo2d1_hd U2434 ( .A(b[14]), .B(n1493), .Y(n1203) );
  oa21d1_hd U2435 ( .A(n2003), .B(n59), .C(n1470), .Y(n1444) );
  clknd2d1_hd U2436 ( .A(n1087), .B(n972), .Y(n892) );
  oa21d1_hd U2437 ( .A(n1), .B(n974), .C(n975), .Y(n973) );
  ivd1_hd U2438 ( .A(n971), .Y(n1087) );
  fad1_hd U2439 ( .A(n1227), .B(n1251), .CI(n1299), .CO(n705), .S(n706) );
  xo2d1_hd U2440 ( .A(b[11]), .B(n1542), .Y(n1227) );
  xo2d1_hd U2441 ( .A(b[2]), .B(n1689), .Y(n1299) );
  xo2d1_hd U2442 ( .A(b[8]), .B(n1591), .Y(n1251) );
  ao222d1_hd U2443 ( .A(n23), .B(a[14]), .C(n25), .D(a[13]), .E(n31), .F(a[12]), .Y(n1618) );
  oa21d1_hd U2444 ( .A(n2016), .B(n9), .C(n1716), .Y(n1690) );
  ao222d1_hd U2445 ( .A(n3), .B(a[20]), .C(n5), .D(a[19]), .E(n11), .F(a[18]), 
        .Y(n1716) );
  fad1_hd U2446 ( .A(n724), .B(n1180), .CI(n1276), .CO(n721), .S(n722) );
  xo2d1_hd U2447 ( .A(b[5]), .B(n1641), .Y(n1276) );
  xo2d1_hd U2448 ( .A(b[17]), .B(n1445), .Y(n1180) );
  oa21d1_hd U2449 ( .A(n1998), .B(n19), .C(n1667), .Y(n1641) );
  clknd2d1_hd U2450 ( .A(n1091), .B(n1004), .Y(n896) );
  oa21d1_hd U2451 ( .A(n1044), .B(n1006), .C(n1007), .Y(n1005) );
  ivd1_hd U2452 ( .A(n1003), .Y(n1091) );
  fad1_hd U2453 ( .A(n1204), .B(n1228), .CI(n733), .CO(n719), .S(n720) );
  xo2d1_hd U2454 ( .A(b[14]), .B(n1494), .Y(n1204) );
  xo2d1_hd U2455 ( .A(b[11]), .B(n1543), .Y(n1228) );
  oa21d1_hd U2456 ( .A(n2005), .B(n49), .C(n1520), .Y(n1494) );
  ao222d1_hd U2457 ( .A(n3), .B(a[19]), .C(n5), .D(a[18]), .E(n11), .F(a[17]), 
        .Y(n1717) );
  clknd2d1_hd U2458 ( .A(n958), .B(n961), .Y(n891) );
  oa21d1_hd U2459 ( .A(n1), .B(n963), .C(n964), .Y(n962) );
  ivd1_hd U2460 ( .A(n966), .Y(n964) );
  fad1_hd U2461 ( .A(n1253), .B(n745), .CI(n1277), .CO(n731), .S(n732) );
  xo2d1_hd U2462 ( .A(b[5]), .B(n1642), .Y(n1277) );
  xo2d1_hd U2463 ( .A(b[8]), .B(n1593), .Y(n1253) );
  oa21d1_hd U2464 ( .A(n2013), .B(n19), .C(n1668), .Y(n1642) );
  fad1_hd U2465 ( .A(n1206), .B(n1230), .CI(n746), .CO(n743), .S(n744) );
  xo2d1_hd U2466 ( .A(b[14]), .B(n1496), .Y(n1206) );
  xo2d1_hd U2467 ( .A(b[11]), .B(n1545), .Y(n1230) );
  oa21d1_hd U2468 ( .A(n2003), .B(n49), .C(n1522), .Y(n1496) );
  fad1_hd U2469 ( .A(n1278), .B(n1254), .CI(n1302), .CO(n741), .S(n742) );
  xo2d1_hd U2470 ( .A(b[5]), .B(n1643), .Y(n1278) );
  xo2d1_hd U2471 ( .A(b[2]), .B(n1692), .Y(n1302) );
  xo2d1_hd U2472 ( .A(b[8]), .B(n1594), .Y(n1254) );
  fad1_hd U2473 ( .A(n758), .B(n1207), .CI(n1303), .CO(n755), .S(n756) );
  xo2d1_hd U2474 ( .A(b[2]), .B(n1693), .Y(n1303) );
  xo2d1_hd U2475 ( .A(b[14]), .B(n1497), .Y(n1207) );
  oa21d1_hd U2476 ( .A(n1998), .B(n9), .C(n1719), .Y(n1693) );
  clknd2d1_hd U2478 ( .A(n1094), .B(n1029), .Y(n899) );
  oa21d1_hd U2479 ( .A(n1044), .B(n1031), .C(n1032), .Y(n1030) );
  ivd1_hd U2480 ( .A(n1034), .Y(n1032) );
  ao222d1_hd U2481 ( .A(n33), .B(a[8]), .C(n35), .D(a[7]), .E(n41), .F(a[6]), 
        .Y(n1572) );
  oa21d1_hd U2482 ( .A(n2011), .B(n19), .C(n1670), .Y(n1644) );
  ao222d1_hd U2483 ( .A(n13), .B(a[14]), .C(n15), .D(a[13]), .E(n21), .F(a[12]), .Y(n1670) );
  ao222d1_hd U2484 ( .A(n23), .B(a[10]), .C(n25), .D(a[9]), .E(n31), .F(a[8]), 
        .Y(n1622) );
  oa21d1_hd U2485 ( .A(n2013), .B(n9), .C(n1720), .Y(n1694) );
  ao222d1_hd U2486 ( .A(n3), .B(a[16]), .C(n5), .D(a[15]), .E(n11), .F(a[14]), 
        .Y(n1720) );
  clknd2d1_hd U2488 ( .A(n1092), .B(n1011), .Y(n897) );
  oa21d1_hd U2489 ( .A(n1044), .B(n1013), .C(n1014), .Y(n1012) );
  ao222d1_hd U2490 ( .A(n33), .B(a[6]), .C(n35), .D(a[5]), .E(n41), .F(a[4]), 
        .Y(n1574) );
  fad1_hd U2491 ( .A(n1209), .B(n778), .CI(n785), .CO(n775), .S(n776) );
  xo2d1_hd U2492 ( .A(b[14]), .B(n1499), .Y(n1209) );
  oa21d1_hd U2493 ( .A(n2000), .B(n49), .C(n1525), .Y(n1499) );
  ao222d1_hd U2494 ( .A(n43), .B(a[3]), .C(n45), .D(a[2]), .E(n51), .F(a[1]), 
        .Y(n1525) );
  ao222d1_hd U2495 ( .A(n13), .B(a[12]), .C(n15), .D(a[11]), .E(n21), .F(a[10]), .Y(n1672) );
  oa21d1_hd U2496 ( .A(n2012), .B(n9), .C(n1721), .Y(n1695) );
  ao222d1_hd U2497 ( .A(n3), .B(a[15]), .C(n5), .D(a[14]), .E(n11), .F(a[13]), 
        .Y(n1721) );
  ao222d1_hd U2498 ( .A(n33), .B(a[5]), .C(n35), .D(a[4]), .E(n41), .F(a[3]), 
        .Y(n1575) );
  oa21d1_hd U2499 ( .A(n2011), .B(n9), .C(n1722), .Y(n1696) );
  ao222d1_hd U2500 ( .A(n3), .B(a[14]), .C(n5), .D(a[13]), .E(n11), .F(a[12]), 
        .Y(n1722) );
  ao222d1_hd U2501 ( .A(n23), .B(a[8]), .C(n25), .D(a[7]), .E(n31), .F(a[6]), 
        .Y(n1624) );
  oa21d1_hd U2502 ( .A(n2008), .B(n19), .C(n1673), .Y(n1647) );
  ao222d1_hd U2503 ( .A(n13), .B(a[11]), .C(n15), .D(a[10]), .E(n21), .F(a[9]), 
        .Y(n1673) );
  ao222d1_hd U2504 ( .A(n13), .B(a[10]), .C(n15), .D(a[9]), .E(n21), .F(a[8]), 
        .Y(n1674) );
  oa21d1_hd U2505 ( .A(n2010), .B(n9), .C(n1723), .Y(n1697) );
  ao222d1_hd U2506 ( .A(n3), .B(a[13]), .C(n5), .D(a[12]), .E(n11), .F(a[11]), 
        .Y(n1723) );
  ao222d1_hd U2507 ( .A(n23), .B(a[7]), .C(n25), .D(a[6]), .E(n31), .F(a[5]), 
        .Y(n1625) );
  had1_hd U2508 ( .A(n801), .B(n1211), .CO(n793), .S(n794) );
  xo2d1_hd U2509 ( .A(b[14]), .B(n1501), .Y(n1211) );
  oa21d1_hd U2510 ( .A(n49), .B(n1761), .C(n1988), .Y(n1501) );
  ao222d1_hd U2511 ( .A(n23), .B(a[6]), .C(n25), .D(a[5]), .E(n31), .F(a[4]), 
        .Y(n1626) );
  fad1_hd U2512 ( .A(n1236), .B(n802), .CI(n807), .CO(n799), .S(n800) );
  xo2d1_hd U2513 ( .A(b[11]), .B(n1551), .Y(n1236) );
  oa21d1_hd U2514 ( .A(n2000), .B(n39), .C(n1577), .Y(n1551) );
  ao222d1_hd U2515 ( .A(n33), .B(a[3]), .C(n35), .D(a[2]), .E(n41), .F(a[1]), 
        .Y(n1577) );
  ao222d1_hd U2516 ( .A(n23), .B(a[5]), .C(n25), .D(a[4]), .E(n31), .F(a[3]), 
        .Y(n1627) );
  oa21d1_hd U2517 ( .A(n2008), .B(n9), .C(n1725), .Y(n1699) );
  ao222d1_hd U2518 ( .A(n3), .B(a[11]), .C(n5), .D(a[10]), .E(n11), .F(a[9]), 
        .Y(n1725) );
  had1_hd U2519 ( .A(n1237), .B(n813), .CO(n807), .S(n808) );
  xo2d1_hd U2520 ( .A(b[11]), .B(n1552), .Y(n1237) );
  oa21d1_hd U2521 ( .A(n1999), .B(n39), .C(n1578), .Y(n1552) );
  ao222d1_hd U2522 ( .A(n33), .B(a[2]), .C(n35), .D(a[1]), .E(n41), .F(a[0]), 
        .Y(n1578) );
  nr2d1_hd U2523 ( .A(a[8]), .B(a[7]), .Y(n1050) );
  clknd2d1_hd U2524 ( .A(a[8]), .B(a[7]), .Y(n1051) );
  ao222d1_hd U2525 ( .A(n13), .B(a[7]), .C(n15), .D(a[6]), .E(n21), .F(a[5]), 
        .Y(n1677) );
  had1_hd U2526 ( .A(b[11]), .B(n1239), .CO(n819), .S(n820) );
  xo2d1_hd U2527 ( .A(b[11]), .B(n1554), .Y(n1239) );
  oa21d1_hd U2528 ( .A(n39), .B(n1762), .C(n1994), .Y(n1554) );
  clknd2d1_hd U2529 ( .A(n1096), .B(n1043), .Y(n901) );
  ivd1_hd U2530 ( .A(n1042), .Y(n1096) );
  ad3d2_hd U2531 ( .A(n1834), .B(n1826), .C(n1818), .Y(n31) );
  nr2d1_hd U2533 ( .A(a[5]), .B(a[6]), .Y(n1058) );
  ivd1_hd U2534 ( .A(n1064), .Y(n1062) );
  clknd2d1_hd U2535 ( .A(a[5]), .B(a[6]), .Y(n1059) );
  clknd2d1_hd U2536 ( .A(a[5]), .B(a[4]), .Y(n1064) );
  ivd1_hd U2537 ( .A(n1063), .Y(n1100) );
  xn2d1_hd U2538 ( .A(b[4]), .B(b[3]), .Y(n1827) );
  xo2d1_hd U2539 ( .A(b[22]), .B(b[23]), .Y(n1829) );
  ad2d1_hd U2540 ( .A(n75), .B(a[23]), .Y(n863) );
  oa21d1_hd U2541 ( .A(n1), .B(n920), .C(n921), .Y(n919) );
  clknd2d1_hd U2542 ( .A(n929), .B(n922), .Y(n920) );
  ao21d1_hd U2543 ( .A(n930), .B(n922), .C(n923), .Y(n921) );
  clknd2d1_hd U2545 ( .A(n922), .B(n925), .Y(n887) );
  oa21d1_hd U2546 ( .A(n1), .B(n927), .C(n928), .Y(n926) );
  ivd1_hd U2547 ( .A(n930), .Y(n928) );
  fad1_hd U2548 ( .A(n842), .B(n1132), .CI(n844), .CO(n459), .S(n460) );
  ivd1_hd U2549 ( .A(b[20]), .Y(n1132) );
  ad2d1_hd U2550 ( .A(b[23]), .B(a[20]), .Y(n842) );
  clknd2d1_hd U2551 ( .A(n1083), .B(n936), .Y(n888) );
  oa21d1_hd U2552 ( .A(n1), .B(n938), .C(n939), .Y(n937) );
  ivd1_hd U2553 ( .A(n935), .Y(n1083) );
  fad1_hd U2554 ( .A(n470), .B(n843), .CI(n1133), .CO(n463), .S(n464) );
  ad2d1_hd U2555 ( .A(b[23]), .B(a[19]), .Y(n843) );
  xo2d1_hd U2556 ( .A(b[20]), .B(n1373), .Y(n1133) );
  oa21d1_hd U2557 ( .A(n1970), .B(n69), .C(n1399), .Y(n1373) );
  clknd2d1_hd U2558 ( .A(n940), .B(n943), .Y(n889) );
  oa21d1_hd U2559 ( .A(n1), .B(n945), .C(n946), .Y(n944) );
  fad1_hd U2560 ( .A(n475), .B(n470), .CI(n1134), .CO(n468), .S(n469) );
  xo2d1_hd U2561 ( .A(b[20]), .B(n1374), .Y(n1134) );
  oa21d1_hd U2562 ( .A(n2020), .B(n69), .C(n1400), .Y(n1374) );
  ao21d1_hd U2563 ( .A(n71), .B(a[22]), .C(n866), .Y(n1400) );
  clknd2d1_hd U2565 ( .A(n1085), .B(n954), .Y(n890) );
  oa21d1_hd U2566 ( .A(n1), .B(n956), .C(n957), .Y(n955) );
  ivd1_hd U2567 ( .A(n953), .Y(n1085) );
  fad1_hd U2568 ( .A(n481), .B(n476), .CI(n1135), .CO(n473), .S(n474) );
  xo2d1_hd U2569 ( .A(b[20]), .B(n1375), .Y(n1135) );
  oa21d1_hd U2570 ( .A(n2019), .B(n69), .C(n1401), .Y(n1375) );
  ao222d1_hd U2571 ( .A(n63), .B(a[23]), .C(n65), .D(a[22]), .E(n71), .F(a[21]), .Y(n1401) );
  ad3d2_hd U2572 ( .A(n1829), .B(n1813), .C(n1821), .Y(n81) );
  fad1_hd U2573 ( .A(n1112), .B(n1136), .CI(n482), .CO(n479), .S(n480) );
  xo2d1_hd U2574 ( .A(b[23]), .B(n1327), .Y(n1112) );
  xo2d1_hd U2575 ( .A(b[20]), .B(n1376), .Y(n1136) );
  oa21d1_hd U2576 ( .A(n2015), .B(n79), .C(n1353), .Y(n1327) );
  fad1_hd U2577 ( .A(n497), .B(n490), .CI(n1161), .CO(n488), .S(n489) );
  xo2d1_hd U2578 ( .A(b[17]), .B(n1426), .Y(n1161) );
  oa21d1_hd U2579 ( .A(n2020), .B(n59), .C(n1452), .Y(n1426) );
  ao21d1_hd U2580 ( .A(n61), .B(a[22]), .C(n869), .Y(n1452) );
  fad1_hd U2581 ( .A(n1113), .B(n1137), .CI(n495), .CO(n486), .S(n487) );
  xo2d1_hd U2582 ( .A(b[23]), .B(n1328), .Y(n1113) );
  xo2d1_hd U2583 ( .A(b[20]), .B(n1377), .Y(n1137) );
  oa21d1_hd U2584 ( .A(n2014), .B(n79), .C(n1354), .Y(n1328) );
  fad1_hd U2585 ( .A(n1163), .B(n1115), .CI(n1139), .CO(n503), .S(n504) );
  xo2d1_hd U2586 ( .A(b[20]), .B(n1379), .Y(n1139) );
  xo2d1_hd U2587 ( .A(b[23]), .B(n1330), .Y(n1115) );
  xo2d1_hd U2588 ( .A(b[17]), .B(n1428), .Y(n1163) );
  fad1_hd U2589 ( .A(n1138), .B(n1162), .CI(n496), .CO(n493), .S(n494) );
  xo2d1_hd U2590 ( .A(b[20]), .B(n1378), .Y(n1138) );
  xo2d1_hd U2591 ( .A(b[17]), .B(n1427), .Y(n1162) );
  oa21d1_hd U2592 ( .A(n2016), .B(n69), .C(n1404), .Y(n1378) );
  fad1_hd U2593 ( .A(n1164), .B(n1140), .CI(n515), .CO(n512), .S(n513) );
  xo2d1_hd U2594 ( .A(b[17]), .B(n1429), .Y(n1164) );
  xo2d1_hd U2595 ( .A(b[20]), .B(n1380), .Y(n1140) );
  oa21d1_hd U2596 ( .A(n2017), .B(n59), .C(n1455), .Y(n1429) );
  fad1_hd U2597 ( .A(n514), .B(n506), .CI(n504), .CO(n501), .S(n502) );
  fad1_hd U2598 ( .A(n1165), .B(n535), .CI(n1189), .CO(n521), .S(n522) );
  xo2d1_hd U2599 ( .A(b[14]), .B(n1479), .Y(n1189) );
  xo2d1_hd U2600 ( .A(b[17]), .B(n1430), .Y(n1165) );
  oa21d1_hd U2601 ( .A(n2019), .B(n49), .C(n1505), .Y(n1479) );
  fad1_hd U2602 ( .A(n523), .B(n1188), .CI(n513), .CO(n510), .S(n511) );
  xo2d1_hd U2603 ( .A(b[14]), .B(n1478), .Y(n1188) );
  oa21d1_hd U2604 ( .A(n2020), .B(n49), .C(n1504), .Y(n1478) );
  ao21d1_hd U2605 ( .A(n51), .B(a[22]), .C(n872), .Y(n1504) );
  fad1_hd U2606 ( .A(n536), .B(n1166), .CI(n546), .CO(n531), .S(n532) );
  xo2d1_hd U2607 ( .A(b[17]), .B(n1431), .Y(n1166) );
  oa21d1_hd U2608 ( .A(n2015), .B(n59), .C(n1457), .Y(n1431) );
  ao222d1_hd U2609 ( .A(n53), .B(a[19]), .C(n55), .D(a[18]), .E(n61), .F(a[17]), .Y(n1457) );
  fad1_hd U2610 ( .A(n533), .B(n524), .CI(n522), .CO(n519), .S(n520) );
  fad1_hd U2611 ( .A(n547), .B(n1191), .CI(n557), .CO(n542), .S(n543) );
  xo2d1_hd U2612 ( .A(b[14]), .B(n1481), .Y(n1191) );
  oa21d1_hd U2613 ( .A(n2017), .B(n49), .C(n1507), .Y(n1481) );
  ao222d1_hd U2614 ( .A(n43), .B(a[21]), .C(n45), .D(a[20]), .E(n51), .F(a[19]), .Y(n1507) );
  fad1_hd U2615 ( .A(n544), .B(n534), .CI(n532), .CO(n529), .S(n530) );
  fad1_hd U2616 ( .A(n558), .B(n1192), .CI(n569), .CO(n553), .S(n554) );
  xo2d1_hd U2617 ( .A(b[14]), .B(n1482), .Y(n1192) );
  oa21d1_hd U2618 ( .A(n2016), .B(n49), .C(n1508), .Y(n1482) );
  ao222d1_hd U2619 ( .A(n43), .B(a[20]), .C(n45), .D(a[19]), .E(n51), .F(a[18]), .Y(n1508) );
  fad1_hd U2620 ( .A(n555), .B(n545), .CI(n543), .CO(n540), .S(n541) );
  fad1_hd U2621 ( .A(n570), .B(n572), .CI(n582), .CO(n565), .S(n566) );
  fad1_hd U2622 ( .A(n567), .B(n556), .CI(n554), .CO(n551), .S(n552) );
  fad1_hd U2623 ( .A(n583), .B(n597), .CI(n595), .CO(n578), .S(n579) );
  fad1_hd U2624 ( .A(n580), .B(n568), .CI(n566), .CO(n563), .S(n564) );
  fad1_hd U2625 ( .A(n593), .B(n581), .CI(n579), .CO(n576), .S(n577) );
  fad1_hd U2626 ( .A(n596), .B(n611), .CI(n609), .CO(n591), .S(n592) );
  fad1_hd U2627 ( .A(n610), .B(n612), .CI(n623), .CO(n605), .S(n606) );
  fad1_hd U2628 ( .A(n594), .B(n607), .CI(n592), .CO(n589), .S(n590) );
  fad1_hd U2629 ( .A(n621), .B(n608), .CI(n606), .CO(n603), .S(n604) );
  nr2d1_hd U2630 ( .A(n272), .B(n275), .Y(n270) );
  fad1_hd U2631 ( .A(n635), .B(n622), .CI(n633), .CO(n617), .S(n618) );
  fad1_hd U2632 ( .A(n637), .B(n639), .CI(n624), .CO(n619), .S(n620) );
  fad1_hd U2633 ( .A(n652), .B(n654), .CI(n665), .CO(n647), .S(n648) );
  fad1_hd U2634 ( .A(n636), .B(n649), .CI(n634), .CO(n631), .S(n632) );
  fad1_hd U2635 ( .A(n663), .B(n650), .CI(n648), .CO(n645), .S(n646) );
  fad1_hd U2636 ( .A(n664), .B(n677), .CI(n675), .CO(n659), .S(n660) );
  fad1_hd U2637 ( .A(n666), .B(n681), .CI(n679), .CO(n661), .S(n662) );
  fad1_hd U2638 ( .A(n693), .B(n682), .CI(n680), .CO(n675), .S(n676) );
  fad1_hd U2639 ( .A(n678), .B(n691), .CI(n689), .CO(n673), .S(n674) );
  fad1_hd U2640 ( .A(n692), .B(n705), .CI(n703), .CO(n687), .S(n688) );
  fad1_hd U2641 ( .A(n707), .B(n1274), .CI(n694), .CO(n689), .S(n690) );
  xo2d1_hd U2642 ( .A(b[5]), .B(n1639), .Y(n1274) );
  oa21d1_hd U2643 ( .A(n2015), .B(n19), .C(n1665), .Y(n1639) );
  ao222d1_hd U2644 ( .A(n13), .B(a[19]), .C(n15), .D(a[18]), .E(n21), .F(a[17]), .Y(n1665) );
  fad1_hd U2645 ( .A(n721), .B(n1275), .CI(n708), .CO(n703), .S(n704) );
  xo2d1_hd U2646 ( .A(b[5]), .B(n1640), .Y(n1275) );
  oa21d1_hd U2647 ( .A(n2014), .B(n19), .C(n1666), .Y(n1640) );
  ao222d1_hd U2648 ( .A(n13), .B(a[18]), .C(n15), .D(a[17]), .E(n21), .F(a[16]), .Y(n1666) );
  fad1_hd U2649 ( .A(n719), .B(n706), .CI(n717), .CO(n701), .S(n702) );
  fad1_hd U2650 ( .A(n1300), .B(n1252), .CI(n722), .CO(n717), .S(n718) );
  xo2d1_hd U2651 ( .A(b[8]), .B(n1592), .Y(n1252) );
  xo2d1_hd U2652 ( .A(b[2]), .B(n1690), .Y(n1300) );
  oa21d1_hd U2653 ( .A(n2011), .B(n29), .C(n1618), .Y(n1592) );
  fad1_hd U2654 ( .A(n720), .B(n731), .CI(n729), .CO(n715), .S(n716) );
  fad1_hd U2655 ( .A(n734), .B(n1229), .CI(n1301), .CO(n729), .S(n730) );
  xo2d1_hd U2656 ( .A(b[2]), .B(n1691), .Y(n1301) );
  xo2d1_hd U2657 ( .A(b[11]), .B(n1544), .Y(n1229) );
  oa21d1_hd U2658 ( .A(n2015), .B(n9), .C(n1717), .Y(n1691) );
  fad1_hd U2659 ( .A(n732), .B(n743), .CI(n741), .CO(n727), .S(n728) );
  fad1_hd U2660 ( .A(n744), .B(n755), .CI(n742), .CO(n739), .S(n740) );
  fad1_hd U2661 ( .A(n756), .B(n1255), .CI(n763), .CO(n751), .S(n752) );
  xo2d1_hd U2662 ( .A(b[8]), .B(n1595), .Y(n1255) );
  oa21d1_hd U2663 ( .A(n2008), .B(n29), .C(n1621), .Y(n1595) );
  ao222d1_hd U2664 ( .A(n23), .B(a[11]), .C(n25), .D(a[10]), .E(n31), .F(a[9]), 
        .Y(n1621) );
  fad1_hd U2665 ( .A(n1231), .B(n1279), .CI(n765), .CO(n753), .S(n754) );
  xo2d1_hd U2666 ( .A(b[11]), .B(n1546), .Y(n1231) );
  xo2d1_hd U2667 ( .A(b[5]), .B(n1644), .Y(n1279) );
  oa21d1_hd U2668 ( .A(n2005), .B(n39), .C(n1572), .Y(n1546) );
  fad1_hd U2669 ( .A(n766), .B(n1280), .CI(n773), .CO(n761), .S(n762) );
  xo2d1_hd U2670 ( .A(b[5]), .B(n1645), .Y(n1280) );
  oa21d1_hd U2671 ( .A(n2010), .B(n19), .C(n1671), .Y(n1645) );
  ao222d1_hd U2672 ( .A(n13), .B(a[13]), .C(n15), .D(a[12]), .E(n21), .F(a[11]), .Y(n1671) );
  fad1_hd U2673 ( .A(n1233), .B(n1257), .CI(n776), .CO(n773), .S(n774) );
  xo2d1_hd U2674 ( .A(b[11]), .B(n1548), .Y(n1233) );
  xo2d1_hd U2675 ( .A(b[8]), .B(n1597), .Y(n1257) );
  oa21d1_hd U2676 ( .A(n2003), .B(n39), .C(n1574), .Y(n1548) );
  fad1_hd U2677 ( .A(n786), .B(n1234), .CI(n1306), .CO(n783), .S(n784) );
  xo2d1_hd U2678 ( .A(b[11]), .B(n1549), .Y(n1234) );
  xo2d1_hd U2679 ( .A(b[2]), .B(n1696), .Y(n1306) );
  oa21d1_hd U2680 ( .A(n2002), .B(n39), .C(n1575), .Y(n1549) );
  fad1_hd U2681 ( .A(n1258), .B(n1282), .CI(n791), .CO(n781), .S(n782) );
  xo2d1_hd U2682 ( .A(b[8]), .B(n1598), .Y(n1258) );
  xo2d1_hd U2683 ( .A(b[5]), .B(n1647), .Y(n1282) );
  oa21d1_hd U2684 ( .A(n2005), .B(n29), .C(n1624), .Y(n1598) );
  fad1_hd U2685 ( .A(n1260), .B(n1284), .CI(n800), .CO(n797), .S(n798) );
  xo2d1_hd U2686 ( .A(b[8]), .B(n1600), .Y(n1260) );
  xo2d1_hd U2687 ( .A(b[5]), .B(n1649), .Y(n1284) );
  oa21d1_hd U2688 ( .A(n2003), .B(n29), .C(n1626), .Y(n1600) );
  clknd2d1_hd U2689 ( .A(n1093), .B(n1022), .Y(n898) );
  oa21d1_hd U2690 ( .A(n1044), .B(n1024), .C(n1025), .Y(n1023) );
  ivd1_hd U2691 ( .A(n1021), .Y(n1093) );
  fad1_hd U2692 ( .A(n808), .B(n1261), .CI(n1309), .CO(n805), .S(n806) );
  xo2d1_hd U2693 ( .A(b[8]), .B(n1601), .Y(n1261) );
  xo2d1_hd U2694 ( .A(b[2]), .B(n1699), .Y(n1309) );
  oa21d1_hd U2695 ( .A(n2002), .B(n29), .C(n1627), .Y(n1601) );
  clknd2d1_hd U2696 ( .A(n1097), .B(n1051), .Y(n902) );
  oa21d1_hd U2697 ( .A(n1055), .B(n1053), .C(n1054), .Y(n1052) );
  ivd1_hd U2698 ( .A(n1050), .Y(n1097) );
  clknd2d1_hd U2699 ( .A(n1095), .B(n1040), .Y(n900) );
  oa21d1_hd U2700 ( .A(n1044), .B(n1042), .C(n1043), .Y(n1041) );
  ivd1_hd U2701 ( .A(n1039), .Y(n1095) );
  ao222d1_hd U2702 ( .A(n13), .B(a[6]), .C(n15), .D(a[5]), .E(n21), .F(a[4]), 
        .Y(n1678) );
  fad1_hd U2703 ( .A(n1263), .B(n820), .CI(n823), .CO(n817), .S(n818) );
  xo2d1_hd U2704 ( .A(b[8]), .B(n1603), .Y(n1263) );
  oa21d1_hd U2705 ( .A(n2000), .B(n29), .C(n1629), .Y(n1603) );
  ao222d1_hd U2706 ( .A(n23), .B(a[3]), .C(n25), .D(a[2]), .E(n31), .F(a[1]), 
        .Y(n1629) );
  oa21d1_hd U2707 ( .A(n2006), .B(n9), .C(n1727), .Y(n1701) );
  ao222d1_hd U2708 ( .A(n3), .B(a[9]), .C(n5), .D(a[8]), .E(n11), .F(a[7]), 
        .Y(n1727) );
  ao222d1_hd U2709 ( .A(n13), .B(a[5]), .C(n15), .D(a[4]), .E(n21), .F(a[3]), 
        .Y(n1679) );
  oa21d1_hd U2710 ( .A(n2005), .B(n9), .C(n1728), .Y(n1702) );
  ao222d1_hd U2711 ( .A(n3), .B(a[8]), .C(n5), .D(a[7]), .E(n11), .F(a[6]), 
        .Y(n1728) );
  had1_hd U2712 ( .A(n1264), .B(n827), .CO(n823), .S(n824) );
  xo2d1_hd U2713 ( .A(b[8]), .B(n1604), .Y(n1264) );
  oa21d1_hd U2714 ( .A(n1999), .B(n29), .C(n1630), .Y(n1604) );
  ao222d1_hd U2715 ( .A(n23), .B(a[2]), .C(n25), .D(a[1]), .E(n31), .F(a[0]), 
        .Y(n1630) );
  ao222d1_hd U2716 ( .A(n3), .B(a[7]), .C(n5), .D(a[6]), .E(n11), .F(a[5]), 
        .Y(n1729) );
  clknd2d1_hd U2717 ( .A(n1098), .B(n1054), .Y(n903) );
  ivd1_hd U2718 ( .A(n1053), .Y(n1098) );
  clknd2d1_hd U2719 ( .A(n1099), .B(n1059), .Y(n904) );
  ao21d1_hd U2720 ( .A(n1065), .B(n1100), .C(n1062), .Y(n1060) );
  ivd1_hd U2721 ( .A(n1058), .Y(n1099) );
  had1_hd U2722 ( .A(b[8]), .B(n1266), .CO(n831), .S(n832) );
  xo2d1_hd U2723 ( .A(b[8]), .B(n1606), .Y(n1266) );
  oa21d1_hd U2724 ( .A(n29), .B(n1762), .C(n1993), .Y(n1606) );
  clknd2d1_hd U2725 ( .A(n1100), .B(n1064), .Y(n905) );
  ad3d2_hd U2726 ( .A(n1835), .B(n1819), .C(n1827), .Y(n21) );
  clknd2d1_hd U2727 ( .A(n1101), .B(n1070), .Y(n906) );
  oa21d1_hd U2728 ( .A(n1074), .B(n1072), .C(n1073), .Y(n1071) );
  ivd1_hd U2729 ( .A(n1069), .Y(n1101) );
  clknd2d1_hd U2730 ( .A(n1102), .B(n1073), .Y(n907) );
  ivd1_hd U2731 ( .A(n1072), .Y(n1102) );
  nr2d1_hd U2732 ( .A(a[2]), .B(a[1]), .Y(n1076) );
  clknd2d1_hd U2733 ( .A(a[2]), .B(a[1]), .Y(n1077) );
  xn2d1_hd U2734 ( .A(b[1]), .B(b[0]), .Y(n1828) );
  ivd1_hd U2735 ( .A(b[0]), .Y(n1820) );
  ad2d1_hd U2736 ( .A(b[23]), .B(a[21]), .Y(n841) );
  clknd2d1_hd U2737 ( .A(n916), .B(n933), .Y(n914) );
  clknd2d1_hd U2738 ( .A(n81), .B(a[23]), .Y(n1347) );
  ivd1_hd U2739 ( .A(n841), .Y(n456) );
  fad1_hd U2740 ( .A(n459), .B(n456), .CI(n1107), .CO(n454), .S(n455) );
  xo2d1_hd U2741 ( .A(b[23]), .B(n1322), .Y(n1107) );
  oa21d1_hd U2742 ( .A(n2020), .B(n79), .C(n1348), .Y(n1322) );
  ao21d1_hd U2743 ( .A(n81), .B(a[22]), .C(n863), .Y(n1348) );
  fad1_hd U2744 ( .A(n463), .B(n460), .CI(n1108), .CO(n457), .S(n458) );
  xo2d1_hd U2745 ( .A(b[23]), .B(n1323), .Y(n1108) );
  oa21d1_hd U2746 ( .A(n2019), .B(n79), .C(n1349), .Y(n1323) );
  ao222d1_hd U2747 ( .A(n73), .B(a[23]), .C(n75), .D(a[22]), .E(n81), .F(a[21]), .Y(n1349) );
  fad1_hd U2748 ( .A(n464), .B(n1109), .CI(n468), .CO(n461), .S(n462) );
  xo2d1_hd U2749 ( .A(b[23]), .B(n1324), .Y(n1109) );
  oa21d1_hd U2750 ( .A(n2018), .B(n79), .C(n1350), .Y(n1324) );
  ao222d1_hd U2751 ( .A(n73), .B(a[22]), .C(n75), .D(a[21]), .E(n81), .F(a[20]), .Y(n1350) );
  fad1_hd U2752 ( .A(n469), .B(n1110), .CI(n473), .CO(n466), .S(n467) );
  xo2d1_hd U2753 ( .A(b[23]), .B(n1325), .Y(n1110) );
  oa21d1_hd U2754 ( .A(n2017), .B(n79), .C(n1351), .Y(n1325) );
  ao222d1_hd U2755 ( .A(n73), .B(a[21]), .C(n75), .D(a[20]), .E(n81), .F(a[19]), .Y(n1351) );
  fad1_hd U2756 ( .A(n474), .B(n1111), .CI(n479), .CO(n471), .S(n472) );
  xo2d1_hd U2757 ( .A(b[23]), .B(n1326), .Y(n1111) );
  oa21d1_hd U2758 ( .A(n2016), .B(n79), .C(n1352), .Y(n1326) );
  ao222d1_hd U2759 ( .A(n73), .B(a[20]), .C(n75), .D(a[19]), .E(n81), .F(a[18]), .Y(n1352) );
  fad1_hd U2760 ( .A(n480), .B(n488), .CI(n486), .CO(n477), .S(n478) );
  fad1_hd U2761 ( .A(n493), .B(n489), .CI(n487), .CO(n484), .S(n485) );
  fad1_hd U2762 ( .A(n494), .B(n503), .CI(n501), .CO(n491), .S(n492) );
  fad1_hd U2763 ( .A(n502), .B(n512), .CI(n510), .CO(n499), .S(n500) );
  fad1_hd U2764 ( .A(n519), .B(n521), .CI(n511), .CO(n508), .S(n509) );
  fad1_hd U2765 ( .A(n520), .B(n531), .CI(n529), .CO(n517), .S(n518) );
  fad1_hd U2766 ( .A(n530), .B(n542), .CI(n540), .CO(n527), .S(n528) );
  fad1_hd U2767 ( .A(n541), .B(n553), .CI(n551), .CO(n538), .S(n539) );
  fad1_hd U2768 ( .A(n552), .B(n565), .CI(n563), .CO(n549), .S(n550) );
  nr2d1_hd U2769 ( .A(n254), .B(n249), .Y(n247) );
  fad1_hd U2770 ( .A(n576), .B(n578), .CI(n564), .CO(n561), .S(n562) );
  fad1_hd U2771 ( .A(n589), .B(n591), .CI(n577), .CO(n574), .S(n575) );
  fad1_hd U2772 ( .A(n603), .B(n605), .CI(n590), .CO(n587), .S(n588) );
  oa21d1_hd U2773 ( .A(n261), .B(n265), .C(n262), .Y(n260) );
  nr2d1_hd U2774 ( .A(n261), .B(n264), .Y(n259) );
  nr2d1_hd U2775 ( .A(n601), .B(n588), .Y(n254) );
  fad1_hd U2776 ( .A(n617), .B(n619), .CI(n604), .CO(n601), .S(n602) );
  ao21d1_hd U2778 ( .A(n270), .B(n279), .C(n271), .Y(n269) );
  clknd2d1_hd U2779 ( .A(n270), .B(n278), .Y(n268) );
  oa21d1_hd U2780 ( .A(n272), .B(n276), .C(n273), .Y(n271) );
  fad1_hd U2781 ( .A(n631), .B(n620), .CI(n618), .CO(n615), .S(n616) );
  fad1_hd U2782 ( .A(n645), .B(n647), .CI(n632), .CO(n629), .S(n630) );
  nr2d1_hd U2783 ( .A(n280), .B(n285), .Y(n278) );
  oa21d1_hd U2784 ( .A(n280), .B(n286), .C(n281), .Y(n279) );
  fad1_hd U2785 ( .A(n659), .B(n661), .CI(n646), .CO(n643), .S(n644) );
  fad1_hd U2786 ( .A(n673), .B(n662), .CI(n660), .CO(n657), .S(n658) );
  fad1_hd U2787 ( .A(n687), .B(n676), .CI(n674), .CO(n671), .S(n672) );
  ao21d1_hd U2788 ( .A(n289), .B(n308), .C(n290), .Y(n288) );
  nr2d1_hd U2789 ( .A(n294), .B(n291), .Y(n289) );
  oa21d1_hd U2790 ( .A(n295), .B(n291), .C(n292), .Y(n290) );
  nr2d1_hd U2791 ( .A(n685), .B(n672), .Y(n285) );
  fad1_hd U2792 ( .A(n701), .B(n690), .CI(n688), .CO(n685), .S(n686) );
  fad1_hd U2793 ( .A(n715), .B(n704), .CI(n702), .CO(n699), .S(n700) );
  fad1_hd U2794 ( .A(n727), .B(n718), .CI(n716), .CO(n713), .S(n714) );
  ao21d1_hd U2796 ( .A(n317), .B(n1977), .C(n312), .Y(n310) );
  clknd2d1_hd U2797 ( .A(n316), .B(n1977), .Y(n309) );
  ivd1_hd U2798 ( .A(n314), .Y(n312) );
  fad1_hd U2799 ( .A(n739), .B(n730), .CI(n728), .CO(n725), .S(n726) );
  fad1_hd U2800 ( .A(n751), .B(n753), .CI(n740), .CO(n737), .S(n738) );
  fad1_hd U2801 ( .A(n761), .B(n754), .CI(n752), .CO(n749), .S(n750) );
  ao21d1_hd U2802 ( .A(n335), .B(n327), .C(n328), .Y(n326) );
  nr2d1_hd U2803 ( .A(n329), .B(n332), .Y(n327) );
  oa21d1_hd U2804 ( .A(n329), .B(n333), .C(n330), .Y(n328) );
  nr2d1_hd U2805 ( .A(n750), .B(n759), .Y(n323) );
  fad1_hd U2806 ( .A(n771), .B(n764), .CI(n762), .CO(n759), .S(n760) );
  oa21d1_hd U2807 ( .A(n336), .B(n353), .C(n337), .Y(n335) );
  ao21d1_hd U2808 ( .A(n344), .B(n1976), .C(n339), .Y(n337) );
  clknd2d1_hd U2809 ( .A(n343), .B(n1976), .Y(n336) );
  ivd1_hd U2810 ( .A(n341), .Y(n339) );
  fad1_hd U2811 ( .A(n781), .B(n774), .CI(n772), .CO(n769), .S(n770) );
  fad1_hd U2812 ( .A(n789), .B(n784), .CI(n782), .CO(n779), .S(n780) );
  fad1_hd U2813 ( .A(n797), .B(n792), .CI(n790), .CO(n787), .S(n788) );
  fad1_hd U2814 ( .A(n805), .B(n1308), .CI(n798), .CO(n795), .S(n796) );
  xo2d1_hd U2815 ( .A(b[2]), .B(n1698), .Y(n1308) );
  oa21d1_hd U2816 ( .A(n2009), .B(n9), .C(n1724), .Y(n1698) );
  ao222d1_hd U2817 ( .A(n3), .B(a[12]), .C(n5), .D(a[11]), .E(n11), .F(a[10]), 
        .Y(n1724) );
  ao21d1_hd U2818 ( .A(n354), .B(n362), .C(n355), .Y(n353) );
  nr2d1_hd U2819 ( .A(n356), .B(n359), .Y(n354) );
  oa21d1_hd U2820 ( .A(n356), .B(n360), .C(n357), .Y(n355) );
  nr2d1_hd U2821 ( .A(n796), .B(n803), .Y(n350) );
  fad1_hd U2822 ( .A(n811), .B(n1285), .CI(n806), .CO(n803), .S(n804) );
  xo2d1_hd U2823 ( .A(b[5]), .B(n1650), .Y(n1285) );
  oa21d1_hd U2824 ( .A(n2005), .B(n19), .C(n1676), .Y(n1650) );
  ao222d1_hd U2825 ( .A(n13), .B(a[8]), .C(n15), .D(a[7]), .E(n21), .F(a[6]), 
        .Y(n1676) );
  oa21d1_hd U2826 ( .A(n363), .B(n375), .C(n364), .Y(n362) );
  clknd2d1_hd U2827 ( .A(n1971), .B(n1978), .Y(n363) );
  ao21d1_hd U2828 ( .A(n1978), .B(n371), .C(n366), .Y(n364) );
  ivd1_hd U2829 ( .A(n368), .Y(n366) );
  fad1_hd U2830 ( .A(n1310), .B(n817), .CI(n812), .CO(n809), .S(n810) );
  xo2d1_hd U2831 ( .A(b[2]), .B(n1700), .Y(n1310) );
  oa21d1_hd U2832 ( .A(n2007), .B(n9), .C(n1726), .Y(n1700) );
  ao222d1_hd U2833 ( .A(n3), .B(a[10]), .C(n5), .D(a[9]), .E(n11), .F(a[8]), 
        .Y(n1726) );
  fad1_hd U2834 ( .A(n1287), .B(n1311), .CI(n818), .CO(n815), .S(n816) );
  xo2d1_hd U2835 ( .A(b[5]), .B(n1652), .Y(n1287) );
  xo2d1_hd U2836 ( .A(b[2]), .B(n1701), .Y(n1311) );
  oa21d1_hd U2837 ( .A(n2003), .B(n19), .C(n1678), .Y(n1652) );
  fad1_hd U2838 ( .A(n824), .B(n1288), .CI(n1312), .CO(n821), .S(n822) );
  xo2d1_hd U2839 ( .A(b[5]), .B(n1653), .Y(n1288) );
  xo2d1_hd U2840 ( .A(b[2]), .B(n1702), .Y(n1312) );
  oa21d1_hd U2841 ( .A(n2002), .B(n19), .C(n1679), .Y(n1653) );
  ao21d1_hd U2842 ( .A(n380), .B(n1979), .C(n377), .Y(n375) );
  ivd1_hd U2843 ( .A(n379), .Y(n377) );
  fad1_hd U2844 ( .A(n1289), .B(n828), .CI(n1313), .CO(n825), .S(n826) );
  xo2d1_hd U2845 ( .A(b[2]), .B(n1703), .Y(n1313) );
  xo2d1_hd U2846 ( .A(b[5]), .B(n1654), .Y(n1289) );
  oa21d1_hd U2847 ( .A(n2004), .B(n9), .C(n1729), .Y(n1703) );
  xo2d1_hd U2848 ( .A(b[2]), .B(n1704), .Y(n1314) );
  oa21d1_hd U2849 ( .A(n2003), .B(n9), .C(n1730), .Y(n1704) );
  ao222d1_hd U2850 ( .A(n3), .B(a[6]), .C(n5), .D(a[5]), .E(n11), .F(a[4]), 
        .Y(n1730) );
  fad1_hd U2851 ( .A(n1290), .B(n832), .CI(n833), .CO(n829), .S(n830) );
  xo2d1_hd U2852 ( .A(b[5]), .B(n1655), .Y(n1290) );
  oa21d1_hd U2853 ( .A(n2000), .B(n19), .C(n1681), .Y(n1655) );
  ao222d1_hd U2854 ( .A(n13), .B(a[3]), .C(n15), .D(a[2]), .E(n21), .F(a[1]), 
        .Y(n1681) );
  xo2d1_hd U2855 ( .A(b[2]), .B(n1705), .Y(n1315) );
  oa21d1_hd U2856 ( .A(n2002), .B(n9), .C(n1731), .Y(n1705) );
  ao222d1_hd U2857 ( .A(n3), .B(a[5]), .C(n5), .D(a[4]), .E(n11), .F(a[3]), 
        .Y(n1731) );
  had1_hd U2858 ( .A(n1291), .B(n835), .CO(n833), .S(n834) );
  xo2d1_hd U2859 ( .A(b[5]), .B(n1656), .Y(n1291) );
  oa21d1_hd U2860 ( .A(n1999), .B(n19), .C(n1682), .Y(n1656) );
  ao222d1_hd U2861 ( .A(n13), .B(a[2]), .C(n15), .D(a[1]), .E(n21), .F(a[0]), 
        .Y(n1682) );
  xo2d1_hd U2862 ( .A(b[2]), .B(n1706), .Y(n1316) );
  oa21d1_hd U2863 ( .A(n2001), .B(n9), .C(n1732), .Y(n1706) );
  ao222d1_hd U2864 ( .A(n3), .B(a[4]), .C(n5), .D(a[3]), .E(n11), .F(a[2]), 
        .Y(n1732) );
  xo2d1_hd U2865 ( .A(b[2]), .B(n1707), .Y(n1317) );
  oa21d1_hd U2866 ( .A(n2000), .B(n9), .C(n1733), .Y(n1707) );
  ao222d1_hd U2867 ( .A(n3), .B(a[3]), .C(n5), .D(a[2]), .E(n11), .F(a[1]), 
        .Y(n1733) );
  had1_hd U2868 ( .A(b[5]), .B(n1293), .CO(n837), .S(n838) );
  xo2d1_hd U2869 ( .A(b[5]), .B(n1658), .Y(n1293) );
  oa21d1_hd U2870 ( .A(n19), .B(n1762), .C(n1992), .Y(n1658) );
  xo3d1_hd U2871 ( .A(n839), .B(n841), .C(n1105), .Y(n450) );
  ad2d1_hd U2872 ( .A(a[23]), .B(b[23]), .Y(n839) );
  ivd1_hd U2873 ( .A(b[23]), .Y(n1105) );
  fad1_hd U2874 ( .A(n456), .B(n840), .CI(n1106), .CO(n451), .S(n452) );
  ad2d1_hd U2875 ( .A(b[23]), .B(a[22]), .Y(n840) );
  xo2d1_hd U2876 ( .A(b[23]), .B(n1321), .Y(n1106) );
  oa21d1_hd U2877 ( .A(n1970), .B(n79), .C(n1347), .Y(n1321) );
  ivd1_hd U2878 ( .A(n187), .Y(n185) );
  nr2d1_hd U2879 ( .A(n454), .B(n452), .Y(n181) );
  clknd2d1_hd U2880 ( .A(n454), .B(n452), .Y(n182) );
  clknd2d1_hd U2881 ( .A(n457), .B(n455), .Y(n187) );
  ivd1_hd U2882 ( .A(n195), .Y(n193) );
  nr2d1_hd U2883 ( .A(n461), .B(n458), .Y(n189) );
  clknd2d1_hd U2884 ( .A(n461), .B(n458), .Y(n190) );
  clknd2d1_hd U2885 ( .A(n466), .B(n462), .Y(n195) );
  ivd1_hd U2886 ( .A(n203), .Y(n201) );
  nr2d1_hd U2887 ( .A(n471), .B(n467), .Y(n197) );
  clknd2d1_hd U2888 ( .A(n471), .B(n467), .Y(n198) );
  clknd2d1_hd U2889 ( .A(n477), .B(n472), .Y(n203) );
  ivd1_hd U2890 ( .A(n211), .Y(n209) );
  nr2d1_hd U2891 ( .A(n484), .B(n478), .Y(n205) );
  clknd2d1_hd U2892 ( .A(n484), .B(n478), .Y(n206) );
  clknd2d1_hd U2893 ( .A(n491), .B(n485), .Y(n211) );
  ivd1_hd U2894 ( .A(n219), .Y(n217) );
  nr2d1_hd U2895 ( .A(n499), .B(n492), .Y(n213) );
  clknd2d1_hd U2896 ( .A(n499), .B(n492), .Y(n214) );
  clknd2d1_hd U2897 ( .A(n508), .B(n500), .Y(n219) );
  ivd1_hd U2898 ( .A(n227), .Y(n225) );
  nr2d1_hd U2899 ( .A(n517), .B(n509), .Y(n221) );
  clknd2d1_hd U2900 ( .A(n517), .B(n509), .Y(n222) );
  clknd2d1_hd U2901 ( .A(n527), .B(n518), .Y(n227) );
  ivd1_hd U2902 ( .A(n235), .Y(n233) );
  nr2d1_hd U2903 ( .A(n538), .B(n528), .Y(n229) );
  clknd2d1_hd U2904 ( .A(n538), .B(n528), .Y(n230) );
  clknd2d1_hd U2905 ( .A(n549), .B(n539), .Y(n235) );
  nr2d1_hd U2908 ( .A(n245), .B(n242), .Y(n240) );
  nr2d1_hd U2910 ( .A(n561), .B(n550), .Y(n237) );
  clknd2d1_hd U2911 ( .A(n561), .B(n550), .Y(n238) );
  nr2d1_hd U2912 ( .A(n574), .B(n562), .Y(n242) );
  ao21d1_hd U2913 ( .A(n247), .B(n260), .C(n248), .Y(n246) );
  oa21d1_hd U2914 ( .A(n249), .B(n255), .C(n250), .Y(n248) );
  clknd2d1_hd U2915 ( .A(n247), .B(n259), .Y(n245) );
  clknd2d1_hd U2916 ( .A(n574), .B(n562), .Y(n243) );
  nr2d1_hd U2917 ( .A(n587), .B(n575), .Y(n249) );
  ivd1_hd U2918 ( .A(n255), .Y(n253) );
  clknd2d1_hd U2919 ( .A(n587), .B(n575), .Y(n250) );
  clknd2d1_hd U2920 ( .A(n601), .B(n588), .Y(n255) );
  oa21d1_hd U2921 ( .A(n266), .B(n257), .C(n258), .Y(n256) );
  ivd1_hd U2922 ( .A(n260), .Y(n258) );
  ivd1_hd U2923 ( .A(n259), .Y(n257) );
  ivd1_hd U2924 ( .A(n254), .Y(n422) );
  nr2d1_hd U2925 ( .A(n602), .B(n615), .Y(n261) );
  clknd2d1_hd U2926 ( .A(n602), .B(n615), .Y(n262) );
  nr2d1_hd U2927 ( .A(n629), .B(n616), .Y(n264) );
  ivd1_hd U2928 ( .A(n267), .Y(n266) );
  nr2d1_hd U2929 ( .A(n643), .B(n630), .Y(n272) );
  clknd2d1_hd U2930 ( .A(n643), .B(n630), .Y(n273) );
  nr2d1_hd U2931 ( .A(n644), .B(n657), .Y(n275) );
  ao21d1_hd U2932 ( .A(n287), .B(n278), .C(n279), .Y(n277) );
  clknd2d1_hd U2933 ( .A(n644), .B(n657), .Y(n276) );
  nr2d1_hd U2934 ( .A(n658), .B(n671), .Y(n280) );
  ivd1_hd U2935 ( .A(n286), .Y(n284) );
  clknd2d1_hd U2936 ( .A(n658), .B(n671), .Y(n281) );
  clknd2d1_hd U2937 ( .A(n685), .B(n672), .Y(n286) );
  ivd1_hd U2938 ( .A(n288), .Y(n287) );
  ivd1_hd U2939 ( .A(n285), .Y(n428) );
  nr2d1_hd U2940 ( .A(n686), .B(n699), .Y(n291) );
  ao21d1_hd U2941 ( .A(n1973), .B(n304), .C(n297), .Y(n295) );
  ivd1_hd U2942 ( .A(n299), .Y(n297) );
  ivd1_hd U2943 ( .A(n302), .Y(n304) );
  clknd2d1_hd U2944 ( .A(n1973), .B(n431), .Y(n294) );
  clknd2d1_hd U2945 ( .A(n686), .B(n699), .Y(n292) );
  clknd2d1_hd U2946 ( .A(n700), .B(n713), .Y(n299) );
  nr2d1_hd U2947 ( .A(n714), .B(n725), .Y(n301) );
  ivd1_hd U2948 ( .A(n301), .Y(n431) );
  clknd2d1_hd U2949 ( .A(n714), .B(n725), .Y(n302) );
  ivd1_hd U2950 ( .A(n308), .Y(n307) );
  clknd2d1_hd U2951 ( .A(n726), .B(n737), .Y(n314) );
  nr2d1_hd U2952 ( .A(n318), .B(n323), .Y(n316) );
  oa21d1_hd U2953 ( .A(n318), .B(n324), .C(n319), .Y(n317) );
  nr2d1_hd U2954 ( .A(n738), .B(n749), .Y(n318) );
  ivd1_hd U2955 ( .A(n324), .Y(n322) );
  clknd2d1_hd U2956 ( .A(n738), .B(n749), .Y(n319) );
  clknd2d1_hd U2957 ( .A(n750), .B(n759), .Y(n324) );
  ivd1_hd U2958 ( .A(n326), .Y(n325) );
  ivd1_hd U2959 ( .A(n323), .Y(n434) );
  nr2d1_hd U2960 ( .A(n760), .B(n769), .Y(n329) );
  clknd2d1_hd U2961 ( .A(n760), .B(n769), .Y(n330) );
  nr2d1_hd U2962 ( .A(n770), .B(n779), .Y(n332) );
  ivd1_hd U2963 ( .A(n335), .Y(n334) );
  clknd2d1_hd U2964 ( .A(n770), .B(n779), .Y(n333) );
  clknd2d1_hd U2965 ( .A(n780), .B(n787), .Y(n341) );
  nr2d1_hd U2966 ( .A(n345), .B(n350), .Y(n343) );
  oa21d1_hd U2967 ( .A(n345), .B(n351), .C(n346), .Y(n344) );
  nr2d1_hd U2968 ( .A(n788), .B(n795), .Y(n345) );
  ivd1_hd U2969 ( .A(n351), .Y(n349) );
  clknd2d1_hd U2970 ( .A(n788), .B(n795), .Y(n346) );
  clknd2d1_hd U2971 ( .A(n796), .B(n803), .Y(n351) );
  ivd1_hd U2972 ( .A(n353), .Y(n352) );
  ivd1_hd U2973 ( .A(n350), .Y(n439) );
  nr2d1_hd U2974 ( .A(n804), .B(n809), .Y(n356) );
  clknd2d1_hd U2975 ( .A(n804), .B(n809), .Y(n357) );
  nr2d1_hd U2976 ( .A(n810), .B(n815), .Y(n359) );
  ivd1_hd U2977 ( .A(n362), .Y(n361) );
  clknd2d1_hd U2978 ( .A(n810), .B(n815), .Y(n360) );
  clknd2d1_hd U2979 ( .A(n816), .B(n821), .Y(n368) );
  ivd1_hd U2980 ( .A(n373), .Y(n371) );
  clknd2d1_hd U2981 ( .A(n822), .B(n825), .Y(n373) );
  ivd1_hd U2982 ( .A(n375), .Y(n374) );
  clknd2d1_hd U2983 ( .A(n826), .B(n829), .Y(n379) );
  oa21d1_hd U2984 ( .A(n383), .B(n381), .C(n382), .Y(n380) );
  ao21d1_hd U2985 ( .A(n388), .B(n1982), .C(n385), .Y(n383) );
  ivd1_hd U2986 ( .A(n387), .Y(n385) );
  nr2d1_hd U2987 ( .A(n830), .B(n1314), .Y(n381) );
  clknd2d1_hd U2988 ( .A(n830), .B(n1314), .Y(n382) );
  clknd2d1_hd U2989 ( .A(n834), .B(n1315), .Y(n387) );
  oa21d1_hd U2990 ( .A(n391), .B(n389), .C(n390), .Y(n388) );
  ao21d1_hd U2991 ( .A(n396), .B(n1981), .C(n393), .Y(n391) );
  ivd1_hd U2992 ( .A(n395), .Y(n393) );
  nr2d1_hd U2993 ( .A(n1316), .B(n836), .Y(n389) );
  clknd2d1_hd U2994 ( .A(n1316), .B(n836), .Y(n390) );
  clknd2d1_hd U2995 ( .A(n1317), .B(n838), .Y(n395) );
  oa21d1_hd U2996 ( .A(n1999), .B(n9), .C(n1734), .Y(n1708) );
  ao222d1_hd U2997 ( .A(n3), .B(a[2]), .C(n5), .D(a[1]), .E(n11), .F(a[0]), 
        .Y(n1734) );
  ivd1_hd U2998 ( .A(n403), .Y(n401) );
  xo2d1_hd U2999 ( .A(b[2]), .B(n1709), .Y(n399) );
  oa21d1_hd U3000 ( .A(n9), .B(n1761), .C(n1984), .Y(n1709) );
  xo2d1_hd U3001 ( .A(b[2]), .B(n1710), .Y(n1320) );
  oa21d1_hd U3002 ( .A(n9), .B(n1762), .C(n1991), .Y(n1710) );
  clknd2d1_hd U3003 ( .A(n1320), .B(b[2]), .Y(n403) );
  clknd2d1_hd U3005 ( .A(n2029), .B(n179), .Y(n132) );
  clknd2d1_hd U3007 ( .A(n451), .B(n450), .Y(n179) );
  xo2d1_hd U3008 ( .A(n133), .B(n183), .Y(product[46]) );
  clknd2d1_hd U3009 ( .A(n405), .B(n182), .Y(n133) );
  ivd1_hd U3010 ( .A(n181), .Y(n405) );
  xn2d1_hd U3011 ( .A(n188), .B(n134), .Y(product[45]) );
  clknd2d1_hd U3012 ( .A(n2028), .B(n187), .Y(n134) );
  xo2d1_hd U3013 ( .A(n135), .B(n191), .Y(product[44]) );
  clknd2d1_hd U3014 ( .A(n407), .B(n190), .Y(n135) );
  ivd1_hd U3015 ( .A(n189), .Y(n407) );
  xn2d1_hd U3016 ( .A(n196), .B(n136), .Y(product[43]) );
  clknd2d1_hd U3017 ( .A(n2027), .B(n195), .Y(n136) );
  xo2d1_hd U3018 ( .A(n137), .B(n199), .Y(product[42]) );
  clknd2d1_hd U3019 ( .A(n409), .B(n198), .Y(n137) );
  ivd1_hd U3020 ( .A(n197), .Y(n409) );
  xn2d1_hd U3021 ( .A(n204), .B(n138), .Y(product[41]) );
  clknd2d1_hd U3022 ( .A(n2026), .B(n203), .Y(n138) );
  xo2d1_hd U3023 ( .A(n139), .B(n207), .Y(product[40]) );
  clknd2d1_hd U3024 ( .A(n411), .B(n206), .Y(n139) );
  ivd1_hd U3025 ( .A(n205), .Y(n411) );
  xn2d1_hd U3026 ( .A(n212), .B(n140), .Y(product[39]) );
  clknd2d1_hd U3027 ( .A(n2025), .B(n211), .Y(n140) );
  xo2d1_hd U3028 ( .A(n141), .B(n215), .Y(product[38]) );
  clknd2d1_hd U3029 ( .A(n413), .B(n214), .Y(n141) );
  ivd1_hd U3030 ( .A(n213), .Y(n413) );
  xn2d1_hd U3031 ( .A(n220), .B(n142), .Y(product[37]) );
  clknd2d1_hd U3032 ( .A(n2022), .B(n219), .Y(n142) );
  xo2d1_hd U3033 ( .A(n143), .B(n223), .Y(product[36]) );
  clknd2d1_hd U3034 ( .A(n415), .B(n222), .Y(n143) );
  ivd1_hd U3035 ( .A(n221), .Y(n415) );
  xn2d1_hd U3036 ( .A(n228), .B(n144), .Y(product[35]) );
  clknd2d1_hd U3037 ( .A(n2021), .B(n227), .Y(n144) );
  xo2d1_hd U3038 ( .A(n145), .B(n231), .Y(product[34]) );
  clknd2d1_hd U3039 ( .A(n417), .B(n230), .Y(n145) );
  ivd1_hd U3040 ( .A(n229), .Y(n417) );
  xn2d1_hd U3041 ( .A(n236), .B(n146), .Y(product[33]) );
  clknd2d1_hd U3042 ( .A(n1980), .B(n235), .Y(n146) );
  xo2d1_hd U3043 ( .A(n147), .B(n239), .Y(product[32]) );
  clknd2d1_hd U3044 ( .A(n419), .B(n238), .Y(n147) );
  ivd1_hd U3045 ( .A(n237), .Y(n419) );
  xn2d1_hd U3046 ( .A(n244), .B(n148), .Y(product[31]) );
  clknd2d1_hd U3047 ( .A(n420), .B(n243), .Y(n148) );
  oa21d1_hd U3048 ( .A(n266), .B(n245), .C(n246), .Y(n244) );
  ivd1_hd U3049 ( .A(n242), .Y(n420) );
  xo2d1_hd U3050 ( .A(n149), .B(n251), .Y(product[30]) );
  clknd2d1_hd U3051 ( .A(n421), .B(n250), .Y(n149) );
  ao21d1_hd U3052 ( .A(n256), .B(n422), .C(n253), .Y(n251) );
  ivd1_hd U3053 ( .A(n249), .Y(n421) );
  xn2d1_hd U3054 ( .A(n256), .B(n150), .Y(product[29]) );
  clknd2d1_hd U3055 ( .A(n422), .B(n255), .Y(n150) );
  xn2d1_hd U3056 ( .A(n263), .B(n151), .Y(product[28]) );
  clknd2d1_hd U3057 ( .A(n423), .B(n262), .Y(n151) );
  oa21d1_hd U3058 ( .A(n266), .B(n264), .C(n265), .Y(n263) );
  ivd1_hd U3059 ( .A(n261), .Y(n423) );
  xo2d1_hd U3060 ( .A(n152), .B(n266), .Y(product[27]) );
  clknd2d1_hd U3061 ( .A(n424), .B(n265), .Y(n152) );
  ivd1_hd U3062 ( .A(n264), .Y(n424) );
  xn2d1_hd U3063 ( .A(n274), .B(n153), .Y(product[26]) );
  clknd2d1_hd U3064 ( .A(n425), .B(n273), .Y(n153) );
  oa21d1_hd U3065 ( .A(n277), .B(n275), .C(n276), .Y(n274) );
  ivd1_hd U3066 ( .A(n272), .Y(n425) );
  xo2d1_hd U3067 ( .A(n154), .B(n277), .Y(product[25]) );
  clknd2d1_hd U3068 ( .A(n426), .B(n276), .Y(n154) );
  ivd1_hd U3069 ( .A(n275), .Y(n426) );
  xo2d1_hd U3070 ( .A(n155), .B(n282), .Y(product[24]) );
  clknd2d1_hd U3071 ( .A(n427), .B(n281), .Y(n155) );
  ao21d1_hd U3072 ( .A(n287), .B(n428), .C(n284), .Y(n282) );
  ivd1_hd U3073 ( .A(n280), .Y(n427) );
  xn2d1_hd U3074 ( .A(n287), .B(n156), .Y(product[23]) );
  clknd2d1_hd U3075 ( .A(n428), .B(n286), .Y(n156) );
  xn2d1_hd U3076 ( .A(n293), .B(n157), .Y(product[22]) );
  clknd2d1_hd U3077 ( .A(n429), .B(n292), .Y(n157) );
  oa21d1_hd U3078 ( .A(n307), .B(n294), .C(n295), .Y(n293) );
  ivd1_hd U3079 ( .A(n291), .Y(n429) );
  xn2d1_hd U3080 ( .A(n300), .B(n158), .Y(product[21]) );
  clknd2d1_hd U3081 ( .A(n1973), .B(n299), .Y(n158) );
  oa21d1_hd U3082 ( .A(n307), .B(n301), .C(n302), .Y(n300) );
  xo2d1_hd U3083 ( .A(n159), .B(n307), .Y(product[20]) );
  clknd2d1_hd U3084 ( .A(n431), .B(n302), .Y(n159) );
  xo2d1_hd U3085 ( .A(n160), .B(n315), .Y(product[19]) );
  clknd2d1_hd U3086 ( .A(n1977), .B(n314), .Y(n160) );
  ao21d1_hd U3087 ( .A(n325), .B(n316), .C(n317), .Y(n315) );
  xo2d1_hd U3088 ( .A(n161), .B(n320), .Y(product[18]) );
  clknd2d1_hd U3089 ( .A(n433), .B(n319), .Y(n161) );
  ao21d1_hd U3090 ( .A(n325), .B(n434), .C(n322), .Y(n320) );
  ivd1_hd U3091 ( .A(n318), .Y(n433) );
  xn2d1_hd U3092 ( .A(n325), .B(n162), .Y(product[17]) );
  clknd2d1_hd U3093 ( .A(n434), .B(n324), .Y(n162) );
  xn2d1_hd U3094 ( .A(n331), .B(n163), .Y(product[16]) );
  clknd2d1_hd U3095 ( .A(n435), .B(n330), .Y(n163) );
  oa21d1_hd U3096 ( .A(n334), .B(n332), .C(n333), .Y(n331) );
  ivd1_hd U3097 ( .A(n329), .Y(n435) );
  xo2d1_hd U3098 ( .A(n164), .B(n334), .Y(product[15]) );
  clknd2d1_hd U3099 ( .A(n436), .B(n333), .Y(n164) );
  ivd1_hd U3100 ( .A(n332), .Y(n436) );
  xo2d1_hd U3101 ( .A(n165), .B(n342), .Y(product[14]) );
  clknd2d1_hd U3102 ( .A(n1976), .B(n341), .Y(n165) );
  ao21d1_hd U3103 ( .A(n352), .B(n343), .C(n344), .Y(n342) );
  xo2d1_hd U3104 ( .A(n166), .B(n347), .Y(product[13]) );
  clknd2d1_hd U3105 ( .A(n438), .B(n346), .Y(n166) );
  ao21d1_hd U3106 ( .A(n352), .B(n439), .C(n349), .Y(n347) );
  ivd1_hd U3107 ( .A(n345), .Y(n438) );
  xn2d1_hd U3108 ( .A(n352), .B(n167), .Y(product[12]) );
  clknd2d1_hd U3109 ( .A(n439), .B(n351), .Y(n167) );
  xn2d1_hd U3110 ( .A(n358), .B(n168), .Y(product[11]) );
  clknd2d1_hd U3111 ( .A(n440), .B(n357), .Y(n168) );
  oa21d1_hd U3112 ( .A(n361), .B(n359), .C(n360), .Y(n358) );
  ivd1_hd U3113 ( .A(n356), .Y(n440) );
  xo2d1_hd U3114 ( .A(n169), .B(n361), .Y(product[10]) );
  clknd2d1_hd U3115 ( .A(n441), .B(n360), .Y(n169) );
  ivd1_hd U3116 ( .A(n359), .Y(n441) );
  xo2d1_hd U3117 ( .A(n170), .B(n369), .Y(product[9]) );
  ao21d1_hd U3118 ( .A(n374), .B(n1971), .C(n371), .Y(n369) );
  clknd2d1_hd U3119 ( .A(n1978), .B(n368), .Y(n170) );
  xn2d1_hd U3120 ( .A(n171), .B(n374), .Y(product[8]) );
  clknd2d1_hd U3121 ( .A(n1971), .B(n373), .Y(n171) );
  xn2d1_hd U3122 ( .A(n172), .B(n380), .Y(product[7]) );
  clknd2d1_hd U3123 ( .A(n1979), .B(n379), .Y(n172) );
  xo2d1_hd U3124 ( .A(n383), .B(n173), .Y(product[6]) );
  clknd2d1_hd U3125 ( .A(n445), .B(n382), .Y(n173) );
  ivd1_hd U3126 ( .A(n381), .Y(n445) );
  xn2d1_hd U3127 ( .A(n388), .B(n174), .Y(product[5]) );
  clknd2d1_hd U3128 ( .A(n1982), .B(n387), .Y(n174) );
  xo2d1_hd U3129 ( .A(n391), .B(n175), .Y(product[4]) );
  clknd2d1_hd U3130 ( .A(n447), .B(n390), .Y(n175) );
  ivd1_hd U3131 ( .A(n389), .Y(n447) );
  xn2d1_hd U3132 ( .A(n176), .B(n396), .Y(product[3]) );
  clknd2d1_hd U3133 ( .A(n1981), .B(n395), .Y(n176) );
  xo2d1_hd U3134 ( .A(n398), .B(n1983), .Y(product[2]) );
  xn2d1_hd U3135 ( .A(n400), .B(n401), .Y(product[1]) );
  ivd1_hd U3136 ( .A(n399), .Y(n400) );
  or2d1_hd U3137 ( .A(n822), .B(n825), .Y(n1971) );
  or2d1_hd U3138 ( .A(n914), .B(n945), .Y(n1972) );
  or2d1_hd U3139 ( .A(n700), .B(n713), .Y(n1973) );
  ao22d1_hd U3140 ( .A(n75), .B(a[0]), .C(n73), .D(a[1]), .Y(n1974) );
  clknd2d1_hd U3141 ( .A(n73), .B(a[0]), .Y(n1975) );
  or2d1_hd U3142 ( .A(n780), .B(n787), .Y(n1976) );
  or2d1_hd U3143 ( .A(n726), .B(n737), .Y(n1977) );
  or2d1_hd U3144 ( .A(n816), .B(n821), .Y(n1978) );
  or2d1_hd U3145 ( .A(n826), .B(n829), .Y(n1979) );
  or2d1_hd U3146 ( .A(n549), .B(n539), .Y(n1980) );
  or2d1_hd U3147 ( .A(n1317), .B(n838), .Y(n1981) );
  or2d1_hd U3148 ( .A(n834), .B(n1315), .Y(n1982) );
  xn2d1_hd U3149 ( .A(b[2]), .B(n1708), .Y(n1983) );
  ao22d1_hd U3150 ( .A(n5), .B(a[0]), .C(n3), .D(a[1]), .Y(n1984) );
  ao22d1_hd U3151 ( .A(n15), .B(a[0]), .C(n13), .D(a[1]), .Y(n1985) );
  ao22d1_hd U3152 ( .A(n25), .B(a[0]), .C(n23), .D(a[1]), .Y(n1986) );
  ao22d1_hd U3153 ( .A(n35), .B(a[0]), .C(n33), .D(a[1]), .Y(n1987) );
  ao22d1_hd U3154 ( .A(n45), .B(a[0]), .C(n43), .D(a[1]), .Y(n1988) );
  ao22d1_hd U3155 ( .A(n55), .B(a[0]), .C(n53), .D(a[1]), .Y(n1989) );
  ao22d1_hd U3156 ( .A(n65), .B(a[0]), .C(n63), .D(a[1]), .Y(n1990) );
  clknd2d1_hd U3157 ( .A(n3), .B(a[0]), .Y(n1991) );
  clknd2d1_hd U3158 ( .A(n13), .B(a[0]), .Y(n1992) );
  clknd2d1_hd U3159 ( .A(n23), .B(a[0]), .Y(n1993) );
  clknd2d1_hd U3160 ( .A(n33), .B(a[0]), .Y(n1994) );
  clknd2d1_hd U3161 ( .A(n43), .B(a[0]), .Y(n1995) );
  clknd2d1_hd U3162 ( .A(n53), .B(a[0]), .Y(n1996) );
  clknd2d1_hd U3163 ( .A(n63), .B(a[0]), .Y(n1997) );
  or2d1_hd U3164 ( .A(n527), .B(n518), .Y(n2021) );
  or2d1_hd U3165 ( .A(n508), .B(n500), .Y(n2022) );
  or2d1_hd U3166 ( .A(a[0]), .B(a[1]), .Y(n2023) );
  scg9d1_hd U3167 ( .A(n914), .B(n946), .C(n915), .Y(n2024) );
  or2d1_hd U3168 ( .A(n491), .B(n485), .Y(n2025) );
  or2d1_hd U3169 ( .A(n477), .B(n472), .Y(n2026) );
  or2d1_hd U3170 ( .A(n466), .B(n462), .Y(n2027) );
  or2d1_hd U3171 ( .A(n457), .B(n455), .Y(n2028) );
  or2d1_hd U3172 ( .A(n451), .B(n450), .Y(n2029) );
  or2d1_hd U3173 ( .A(n1320), .B(b[2]), .Y(n2030) );
  ad2d1_hd U3174 ( .A(n2030), .B(n403), .Y(product[0]) );
  clknd2d1_hd U1 ( .A(a[0]), .B(a[1]), .Y(n1078) );
  xo2d1_hd U2 ( .A(b[11]), .B(b[10]), .Y(n1833) );
  xo2d1_hd U3 ( .A(b[14]), .B(b[13]), .Y(n1832) );
  nr2d2_hd U4 ( .A(n1831), .B(n1815), .Y(n53) );
  xn2d1_hd U5 ( .A(b[15]), .B(b[14]), .Y(n1815) );
  ao21d2_hd U6 ( .A(n212), .B(n2025), .C(n209), .Y(n207) );
  or2bd2_hd U7 ( .B(n1813), .AN(n1829), .Y(n79) );
  nr2d1_hd U9 ( .A(n1003), .B(n1010), .Y(n997) );
  or2bd2_hd U10 ( .B(n1816), .AN(n1832), .Y(n49) );
  xo2d1_hd U11 ( .A(n955), .B(n890), .Y(n2016) );
  xo2d1_hd U12 ( .A(n926), .B(n887), .Y(n2019) );
  oa21d1_hd U13 ( .A(n309), .B(n326), .C(n310), .Y(n308) );
  ao21d4_hd U20 ( .A(n236), .B(n1980), .C(n233), .Y(n231) );
  oa21d4_hd U21 ( .A(n239), .B(n237), .C(n238), .Y(n236) );
  oa21d2_hd U23 ( .A(n223), .B(n221), .C(n222), .Y(n220) );
  had1_hd U24 ( .A(n1210), .B(n793), .CO(n785), .S(n786) );
  xo2d1_hd U25 ( .A(b[8]), .B(b[7]), .Y(n1834) );
  xn2d1_hd U26 ( .A(b[6]), .B(b[5]), .Y(n1818) );
  xo2d1_hd U27 ( .A(n1030), .B(n899), .Y(n2008) );
  xn2d1_hd U28 ( .A(b[9]), .B(b[8]), .Y(n1817) );
  nr2d1_hd U29 ( .A(a[9]), .B(a[10]), .Y(n1039) );
  nr2bd2_hd U30 ( .AN(n1818), .B(n1826), .Y(n25) );
  nr2d2_hd U31 ( .A(n1834), .B(n1818), .Y(n23) );
  xo2d1_hd U32 ( .A(n1012), .B(n897), .Y(n2010) );
  xn2d1_hd U33 ( .A(b[12]), .B(b[13]), .Y(n1824) );
  xo2d1_hd U34 ( .A(n994), .B(n895), .Y(n2012) );
  xo2d1_hd U35 ( .A(b[16]), .B(b[17]), .Y(n1831) );
  xn2d1_hd U36 ( .A(b[18]), .B(b[17]), .Y(n1814) );
  ivd1_hd U37 ( .A(a[0]), .Y(n1762) );
  xo2d1_hd U38 ( .A(b[2]), .B(b[1]), .Y(n1836) );
  or2bd2_hd U39 ( .B(n1819), .AN(n1835), .Y(n19) );
  fad1_hd U40 ( .A(n1250), .B(n709), .CI(n1202), .CO(n693), .S(n694) );
  nr2d2_hd U41 ( .A(n1832), .B(n1816), .Y(n43) );
  nr2bd2_hd U42 ( .AN(n1816), .B(n1824), .Y(n45) );
  nr2bd2_hd U43 ( .AN(n1815), .B(n1823), .Y(n55) );
  or2bd2_hd U44 ( .B(n1815), .AN(n1831), .Y(n59) );
  nr2d2_hd U45 ( .A(n1830), .B(n1814), .Y(n63) );
  nr2d1_hd U46 ( .A(n953), .B(n960), .Y(n951) );
  xn2d1_hd U47 ( .A(b[21]), .B(b[20]), .Y(n1813) );
  clknd2d1_hd U48 ( .A(n997), .B(n981), .Y(n979) );
  ao21d2_hd U8 ( .A(n204), .B(n2026), .C(n201), .Y(n199) );
  oa21d1_hd U14 ( .A(n1066), .B(n1046), .C(n1047), .Y(n1045) );
  oa21d2_hd U15 ( .A(n207), .B(n205), .C(n206), .Y(n204) );
  xn2d2_hd U16 ( .A(n180), .B(n132), .Y(product[47]) );
  oa21d2_hd U17 ( .A(n246), .B(n242), .C(n243), .Y(n241) );
  ao21d4_hd U18 ( .A(n228), .B(n2021), .C(n225), .Y(n223) );
  oa21d8_hd U19 ( .A(n231), .B(n229), .C(n230), .Y(n228) );
  oa21d4_hd U22 ( .A(n199), .B(n197), .C(n198), .Y(n196) );
  ao21d2_hd U49 ( .A(n240), .B(n267), .C(n241), .Y(n239) );
  oa21d2_hd U50 ( .A(n268), .B(n288), .C(n269), .Y(n267) );
  ivd6_hd U51 ( .A(n1045), .Y(n1044) );
  ao21d1_hd U52 ( .A(n188), .B(n2028), .C(n185), .Y(n183) );
  oa21d2_hd U53 ( .A(n191), .B(n189), .C(n190), .Y(n188) );
  oa21d2_hd U54 ( .A(n215), .B(n213), .C(n214), .Y(n212) );
  nr2d2_hd U55 ( .A(n1829), .B(n1813), .Y(n73) );
  ao21d2_hd U56 ( .A(n220), .B(n2022), .C(n217), .Y(n215) );
  oa21d1_hd U57 ( .A(n183), .B(n181), .C(n182), .Y(n180) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_float_multiplier_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module float_multiplier ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n469,
         n502, N33, guard, round_bit, sticky, N41, N45, N85, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N286,
         N287, N288, N289, N290, N291, N292, N350, N380, N382, N406, N408,
         N419, N430, N463, N498, N501, N502, C76_DATA2_0, C76_DATA2_1,
         C76_DATA2_2, C76_DATA2_3, C76_DATA2_4, C76_DATA2_5, C76_DATA2_6,
         C76_DATA2_7, C76_DATA2_8, C76_DATA2_9, C72_DATA2_0, C72_DATA2_1,
         C72_DATA2_2, C72_DATA2_3, C72_DATA2_4, C72_DATA2_5, C72_DATA2_6,
         C72_DATA2_7, C72_DATA2_8, C72_DATA2_9, n4, n5, n6, n7, n8, n9, C1_Z_9,
         C1_Z_8, C1_Z_7, C1_Z_6, C1_Z_5, C1_Z_4, C1_Z_3, C1_Z_2, C1_Z_1,
         C1_Z_0, C2_Z_0, n1, DP_OP_105_124_8121_n9, DP_OP_105_124_8121_n8,
         DP_OP_105_124_8121_n7, DP_OP_105_124_8121_n6, DP_OP_105_124_8121_n5,
         DP_OP_105_124_8121_n4, DP_OP_105_124_8121_n3, DP_OP_102_127_8889_n9,
         DP_OP_102_127_8889_n8, DP_OP_102_127_8889_n7, DP_OP_102_127_8889_n6,
         DP_OP_102_127_8889_n5, DP_OP_102_127_8889_n4, DP_OP_102_127_8889_n3,
         n37, n39, n40, n41, n45, n46, n47, n49, n50, n51, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n2, n3, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n48, n72, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267,
         n269, n271, n273, n275, n277, n279, n281, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n301, n303, n305, n307, n309, n311, n313, n315, n317,
         n319, n321, n323, n325, n327, n329, n331, n333, n335, n337, n339,
         n341, n343, n344, n346, n347, n349, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n552;
  wire   [3:1] state;
  wire   [9:0] a_e;
  wire   [23:0] a_m;
  wire   [9:0] b_e;
  wire   [23:0] b_m;
  wire   [49:2] product;
  wire   [9:0] z_e;
  wire   [23:0] z_m;

  ivd1_hd U11 ( .A(i_RST), .Y(n4) );
  ivd1_hd U14 ( .A(i_RST), .Y(n5) );
  ivd1_hd U15 ( .A(i_RST), .Y(n6) );
  ivd1_hd U16 ( .A(i_RST), .Y(n7) );
  ivd1_hd U17 ( .A(i_RST), .Y(n8) );
  ivd1_hd U18 ( .A(i_RST), .Y(n9) );
  fad1_hd DP_OP_105_124_8121_U11 ( .A(n157), .B(n208), .CI(
        DP_OP_105_124_8121_n9), .CO(DP_OP_105_124_8121_n8), .S(C76_DATA2_1) );
  fad1_hd DP_OP_105_124_8121_U10 ( .A(n157), .B(n209), .CI(
        DP_OP_105_124_8121_n8), .CO(DP_OP_105_124_8121_n7), .S(C76_DATA2_2) );
  fad1_hd DP_OP_105_124_8121_U9 ( .A(n157), .B(n210), .CI(
        DP_OP_105_124_8121_n7), .CO(DP_OP_105_124_8121_n6), .S(C76_DATA2_3) );
  fad1_hd DP_OP_105_124_8121_U8 ( .A(n157), .B(n211), .CI(
        DP_OP_105_124_8121_n6), .CO(DP_OP_105_124_8121_n5), .S(C76_DATA2_4) );
  fad1_hd DP_OP_105_124_8121_U7 ( .A(n157), .B(n212), .CI(
        DP_OP_105_124_8121_n5), .CO(DP_OP_105_124_8121_n4), .S(C76_DATA2_5) );
  fad1_hd DP_OP_105_124_8121_U6 ( .A(n157), .B(n213), .CI(
        DP_OP_105_124_8121_n4), .CO(DP_OP_105_124_8121_n3), .S(C76_DATA2_6) );
  fad1_hd DP_OP_102_127_8889_U11 ( .A(n157), .B(C1_Z_1), .CI(
        DP_OP_102_127_8889_n9), .CO(DP_OP_102_127_8889_n8), .S(C72_DATA2_1) );
  fad1_hd DP_OP_102_127_8889_U10 ( .A(n157), .B(C1_Z_2), .CI(
        DP_OP_102_127_8889_n8), .CO(DP_OP_102_127_8889_n7), .S(C72_DATA2_2) );
  fad1_hd DP_OP_102_127_8889_U9 ( .A(n157), .B(C1_Z_3), .CI(
        DP_OP_102_127_8889_n7), .CO(DP_OP_102_127_8889_n6), .S(C72_DATA2_3) );
  fad1_hd DP_OP_102_127_8889_U8 ( .A(n157), .B(C1_Z_4), .CI(
        DP_OP_102_127_8889_n6), .CO(DP_OP_102_127_8889_n5), .S(C72_DATA2_4) );
  fad1_hd DP_OP_102_127_8889_U7 ( .A(n157), .B(C1_Z_5), .CI(
        DP_OP_102_127_8889_n5), .CO(DP_OP_102_127_8889_n4), .S(C72_DATA2_5) );
  fad1_hd DP_OP_102_127_8889_U6 ( .A(n157), .B(C1_Z_6), .CI(
        DP_OP_102_127_8889_n4), .CO(DP_OP_102_127_8889_n3), .S(C72_DATA2_6) );
  nr2d1_hd U186 ( .A(n139), .B(n135), .Y(n132) );
  or2d2_hd U188 ( .A(n201), .B(n191), .Y(n157) );
  or2d1_hd U189 ( .A(n217), .B(n72), .Y(n191) );
  clknd2d2_hd U193 ( .A(n129), .B(n136), .Y(n144) );
  scg2d1_hd U198 ( .A(N45), .B(n417), .C(n99), .D(n298), .Y(n212) );
  scg2d1_hd U199 ( .A(N45), .B(n448), .C(n162), .D(n292), .Y(C1_Z_5) );
  scg2d1_hd U200 ( .A(N45), .B(n416), .C(n99), .D(n297), .Y(n211) );
  scg2d1_hd U201 ( .A(N45), .B(n447), .C(n162), .D(n291), .Y(C1_Z_4) );
  scg2d1_hd U202 ( .A(N45), .B(n445), .C(n162), .D(n289), .Y(C1_Z_2) );
  scg2d1_hd U203 ( .A(N45), .B(n414), .C(n99), .D(n295), .Y(n209) );
  scg2d1_hd U204 ( .A(N45), .B(n446), .C(n162), .D(n290), .Y(C1_Z_3) );
  scg2d1_hd U205 ( .A(N45), .B(n418), .C(n99), .D(n299), .Y(n213) );
  scg2d1_hd U206 ( .A(N45), .B(n444), .C(n162), .D(n258), .Y(C1_Z_1) );
  scg2d1_hd U207 ( .A(N45), .B(n449), .C(n162), .D(n293), .Y(C1_Z_6) );
  scg2d1_hd U208 ( .A(N45), .B(n415), .C(n99), .D(n296), .Y(n210) );
  scg2d1_hd U209 ( .A(N45), .B(n413), .C(n99), .D(n262), .Y(n208) );
  scg2d1_hd U210 ( .A(N45), .B(n412), .C(n99), .D(n294), .Y(n207) );
  clknd2d1_hd U211 ( .A(n198), .B(n199), .Y(n100) );
  clknd2d1_hd U212 ( .A(n257), .B(n190), .Y(n201) );
  clknd2d1_hd U213 ( .A(n154), .B(n155), .Y(n153) );
  ivd1_hd U214 ( .A(n217), .Y(n205) );
  clknd2d1_hd U215 ( .A(n72), .B(n217), .Y(n193) );
  clknd2d1_hd U216 ( .A(n167), .B(n148), .Y(n163) );
  ivd1_hd U217 ( .A(n285), .Y(n190) );
  nr2bd1_hd U218 ( .AN(n217), .B(n72), .Y(n199) );
  scg2d1_hd U219 ( .A(N45), .B(n419), .C(n99), .D(n263), .Y(n214) );
  clknd2d1_hd U220 ( .A(n388), .B(n203), .Y(n119) );
  clknd2d1_hd U221 ( .A(n142), .B(n141), .Y(n204) );
  clknd2d1_hd U222 ( .A(n150), .B(n152), .Y(n149) );
  clknd2d1_hd U223 ( .A(n85), .B(n84), .Y(n88) );
  clknd2d1_hd U224 ( .A(n91), .B(n90), .Y(n94) );
  clknd2d1_hd U225 ( .A(n257), .B(n285), .Y(n196) );
  clknd2d1_hd U226 ( .A(n51), .B(n118), .Y(n111) );
  scg2d1_hd U227 ( .A(N45), .B(n443), .C(n162), .D(n288), .Y(C1_Z_0) );
  scg2d1_hd U228 ( .A(N45), .B(n451), .C(n162), .D(n259), .Y(C1_Z_7) );
  ivd2_hd U230 ( .A(n100), .Y(n99) );
  ivd1_hd U231 ( .A(n199), .Y(n192) );
  scg2d1_hd U232 ( .A(N45), .B(n406), .C(n99), .D(n231), .Y(b_m[17]) );
  scg2d1_hd U233 ( .A(N45), .B(n394), .C(n99), .D(n223), .Y(b_m[5]) );
  scg2d1_hd U235 ( .A(N45), .B(n397), .C(n99), .D(n225), .Y(b_m[8]) );
  scg2d1_hd U236 ( .A(N45), .B(n409), .C(n99), .D(n254), .Y(b_m[20]) );
  scg2d1_hd U237 ( .A(N45), .B(n400), .C(n99), .D(n227), .Y(b_m[11]) );
  scg2d1_hd U238 ( .A(N45), .B(n391), .C(n99), .D(n221), .Y(b_m[2]) );
  xo2d1_hd U239 ( .A(C1_Z_8), .B(n76), .Y(C72_DATA2_8) );
  scg2d1_hd U240 ( .A(N45), .B(n411), .C(n99), .D(n255), .Y(b_m[22]) );
  scg2d1_hd U241 ( .A(N45), .B(n410), .C(n99), .D(n455), .Y(b_m[21]) );
  scg2d1_hd U242 ( .A(N45), .B(n408), .C(n99), .D(n253), .Y(b_m[19]) );
  scg2d1_hd U243 ( .A(N45), .B(n407), .C(n99), .D(n462), .Y(b_m[18]) );
  xo2d1_hd U244 ( .A(n215), .B(n80), .Y(C76_DATA2_8) );
  xo2d1_hd U245 ( .A(n216), .B(n81), .Y(C76_DATA2_9) );
  scg2d1_hd U246 ( .A(n99), .B(n452), .C(n162), .D(n461), .Y(n197) );
  clknd2d1_hd U247 ( .A(i_Z_ACK), .B(o_Z_STB), .Y(n502) );
  clknd2d1_hd U248 ( .A(i_AB_STB), .B(o_AB_ACK), .Y(n469) );
  clknd2d1_hd U249 ( .A(n127), .B(n128), .Y(n470) );
  xo2d1_hd U250 ( .A(n386), .B(n98), .Y(N292) );
  clknd2d1_hd U251 ( .A(n97), .B(n96), .Y(n98) );
  clknd2d1_hd U252 ( .A(n41), .B(n112), .Y(N502) );
  scg2d1_hd U253 ( .A(N45), .B(n441), .C(n162), .D(n251), .Y(a_m[21]) );
  scg2d1_hd U254 ( .A(N45), .B(n440), .C(n162), .D(n250), .Y(a_m[20]) );
  scg2d1_hd U255 ( .A(N45), .B(n439), .C(n162), .D(n249), .Y(a_m[19]) );
  scg2d1_hd U256 ( .A(N45), .B(n438), .C(n162), .D(n248), .Y(a_m[18]) );
  scg2d1_hd U257 ( .A(N45), .B(n437), .C(n162), .D(n247), .Y(a_m[17]) );
  scg2d1_hd U258 ( .A(N45), .B(n436), .C(n162), .D(n246), .Y(a_m[16]) );
  scg2d1_hd U259 ( .A(N45), .B(n435), .C(n162), .D(n245), .Y(a_m[15]) );
  scg2d1_hd U260 ( .A(N45), .B(n434), .C(n162), .D(n244), .Y(a_m[14]) );
  scg2d1_hd U261 ( .A(N45), .B(n433), .C(n162), .D(n243), .Y(a_m[13]) );
  scg2d1_hd U262 ( .A(N45), .B(n432), .C(n162), .D(n242), .Y(a_m[12]) );
  scg2d1_hd U263 ( .A(N45), .B(n431), .C(n162), .D(n241), .Y(a_m[11]) );
  scg2d1_hd U264 ( .A(N45), .B(n430), .C(n162), .D(n240), .Y(a_m[10]) );
  scg2d1_hd U265 ( .A(N45), .B(n429), .C(n162), .D(n239), .Y(a_m[9]) );
  scg2d1_hd U266 ( .A(N45), .B(n428), .C(n162), .D(n238), .Y(a_m[8]) );
  scg2d1_hd U267 ( .A(N45), .B(n427), .C(n162), .D(n237), .Y(a_m[7]) );
  scg2d1_hd U268 ( .A(N45), .B(n426), .C(n162), .D(n236), .Y(a_m[6]) );
  scg2d1_hd U269 ( .A(N45), .B(n425), .C(n162), .D(n235), .Y(a_m[5]) );
  scg2d1_hd U270 ( .A(N45), .B(n424), .C(n162), .D(n234), .Y(a_m[4]) );
  scg2d1_hd U271 ( .A(N45), .B(n423), .C(n162), .D(n233), .Y(a_m[3]) );
  scg2d1_hd U272 ( .A(N45), .B(n422), .C(n162), .D(n232), .Y(a_m[2]) );
  scg2d1_hd U273 ( .A(N45), .B(n421), .C(n162), .D(n286), .Y(a_m[1]) );
  xo2d1_hd U274 ( .A(C1_Z_9), .B(n77), .Y(C72_DATA2_9) );
  xo2d1_hd U275 ( .A(n207), .B(n206), .Y(C76_DATA2_0) );
  scg2d1_hd U276 ( .A(N45), .B(n405), .C(n99), .D(n230), .Y(b_m[16]) );
  scg2d1_hd U277 ( .A(N45), .B(n404), .C(n99), .D(n460), .Y(b_m[15]) );
  scg2d1_hd U278 ( .A(N45), .B(n402), .C(n99), .D(n228), .Y(b_m[13]) );
  scg2d1_hd U279 ( .A(N45), .B(n401), .C(n99), .D(n454), .Y(b_m[12]) );
  scg2d1_hd U280 ( .A(N45), .B(n399), .C(n99), .D(n226), .Y(b_m[10]) );
  scg2d1_hd U281 ( .A(N45), .B(n398), .C(n99), .D(n456), .Y(b_m[9]) );
  scg2d1_hd U282 ( .A(N45), .B(n396), .C(n99), .D(n224), .Y(b_m[7]) );
  scg2d1_hd U283 ( .A(N45), .B(n395), .C(n99), .D(n457), .Y(b_m[6]) );
  scg2d1_hd U284 ( .A(N45), .B(n393), .C(n99), .D(n222), .Y(b_m[4]) );
  scg2d1_hd U285 ( .A(N45), .B(n392), .C(n99), .D(n453), .Y(b_m[3]) );
  scg2d1_hd U286 ( .A(N45), .B(n390), .C(n99), .D(n287), .Y(b_m[1]) );
  xo2d1_hd U287 ( .A(i_B[31]), .B(i_A[31]), .Y(N33) );
  ivd1_hd U288 ( .A(N41), .Y(n73) );
  or2d1_hd U289 ( .A(n201), .B(n193), .Y(n37) );
  scg9d1_hd U291 ( .A(n461), .B(n164), .C(n157), .Y(n39) );
  or2d1_hd U292 ( .A(n469), .B(n73), .Y(n40) );
  ivd4_hd U293 ( .A(n157), .Y(N45) );
  or2d1_hd U294 ( .A(n193), .B(n165), .Y(n41) );
  xo2d1_hd U297 ( .A(C1_Z_0), .B(C2_Z_0), .Y(C72_DATA2_0) );
  nr2ad1_hd U298 ( .A(n217), .B(n201), .Y(C2_Z_0) );
  oa21d2_hd U299 ( .A(n190), .B(n191), .C(n37), .Y(n1) );
  nr2ad1_hd U300 ( .A(n165), .B(n166), .Y(n147) );
  oa21d2_hd U302 ( .A(n158), .B(n159), .C(n160), .Y(N419) );
  nr2d4_hd U303 ( .A(n191), .B(n196), .Y(n115) );
  ivd1_hd U304 ( .A(n41), .Y(n46) );
  ivd1_hd U305 ( .A(n41), .Y(n47) );
  ivd1_hd U307 ( .A(n37), .Y(n49) );
  ivd1_hd U308 ( .A(n37), .Y(n50) );
  ivd1_hd U309 ( .A(n37), .Y(n51) );
  oa21d2_hd U325 ( .A(n161), .B(n159), .C(n39), .Y(N408) );
  scg2d1_hd U327 ( .A(n47), .B(n352), .C(n102), .D(n48), .Y(round_bit) );
  nr2d4_hd U328 ( .A(n191), .B(n202), .Y(n102) );
  nr2d4_hd U331 ( .A(n201), .B(n166), .Y(n162) );
  clknd2d1_hd U332 ( .A(n72), .B(n205), .Y(n166) );
  ivd1_hd U334 ( .A(DP_OP_102_127_8889_n3), .Y(n75) );
  ivd1_hd U335 ( .A(C1_Z_7), .Y(n74) );
  ao22d1_hd U336 ( .A(C1_Z_7), .B(n75), .C(DP_OP_102_127_8889_n3), .D(n74), 
        .Y(C72_DATA2_7) );
  nr2d1_hd U337 ( .A(C1_Z_7), .B(DP_OP_102_127_8889_n3), .Y(n76) );
  nr3d1_hd U338 ( .A(DP_OP_102_127_8889_n3), .B(C1_Z_7), .C(C1_Z_8), .Y(n77)
         );
  nd2bd1_hd U339 ( .AN(C1_Z_0), .B(C2_Z_0), .Y(DP_OP_102_127_8889_n9) );
  ivd1_hd U340 ( .A(DP_OP_105_124_8121_n3), .Y(n79) );
  ivd1_hd U341 ( .A(n214), .Y(n78) );
  ao22d1_hd U342 ( .A(n214), .B(n79), .C(DP_OP_105_124_8121_n3), .D(n78), .Y(
        C76_DATA2_7) );
  nr2d1_hd U343 ( .A(n214), .B(DP_OP_105_124_8121_n3), .Y(n80) );
  nr3d1_hd U344 ( .A(DP_OP_105_124_8121_n3), .B(n214), .C(n215), .Y(n81) );
  nd2bd1_hd U345 ( .AN(n207), .B(n206), .Y(DP_OP_105_124_8121_n9) );
  ivd1_hd U346 ( .A(n380), .Y(n82) );
  ao22d1_hd U347 ( .A(n380), .B(n143), .C(n379), .D(n82), .Y(N286) );
  nr2d1_hd U348 ( .A(n380), .B(n379), .Y(n85) );
  ivd1_hd U349 ( .A(n85), .Y(n83) );
  ivd1_hd U350 ( .A(n381), .Y(n84) );
  ao22d1_hd U351 ( .A(n381), .B(n85), .C(n83), .D(n84), .Y(N287) );
  ivd1_hd U352 ( .A(n88), .Y(n87) );
  ivd1_hd U353 ( .A(n382), .Y(n86) );
  ao22d1_hd U354 ( .A(n382), .B(n87), .C(n88), .D(n86), .Y(N288) );
  nr2d1_hd U355 ( .A(n382), .B(n88), .Y(n91) );
  ivd1_hd U356 ( .A(n91), .Y(n89) );
  ivd1_hd U357 ( .A(n383), .Y(n90) );
  ao22d1_hd U358 ( .A(n383), .B(n91), .C(n89), .D(n90), .Y(N289) );
  ivd1_hd U359 ( .A(n94), .Y(n93) );
  ivd1_hd U360 ( .A(n384), .Y(n92) );
  ao22d1_hd U361 ( .A(n384), .B(n93), .C(n94), .D(n92), .Y(N290) );
  nr2d1_hd U362 ( .A(n384), .B(n94), .Y(n96) );
  ivd1_hd U363 ( .A(n96), .Y(n95) );
  ivd1_hd U364 ( .A(n385), .Y(n97) );
  ao22d1_hd U365 ( .A(n385), .B(n96), .C(n95), .D(n97), .Y(N291) );
  nr2bd1_hd U366 ( .AN(n265), .B(n100), .Y(n216) );
  nr2bd1_hd U367 ( .AN(n264), .B(n100), .Y(n215) );
  oa22ad1_hd U368 ( .A(n218), .B(n41), .C(n102), .D(n103), .Y(sticky) );
  nr4d1_hd U369 ( .A(product[11]), .B(product[10]), .C(n104), .D(n105), .Y(
        n101) );
  nd4d1_hd U370 ( .A(n106), .B(n107), .C(n108), .D(n109), .Y(n105) );
  nr4d1_hd U371 ( .A(product[4]), .B(product[6]), .C(product[5]), .D(
        product[3]), .Y(n109) );
  nr4d1_hd U372 ( .A(product[2]), .B(product[22]), .C(product[21]), .D(
        product[18]), .Y(n108) );
  nr4d1_hd U373 ( .A(product[16]), .B(product[12]), .C(product[14]), .D(
        product[13]), .Y(n107) );
  nr4d1_hd U374 ( .A(product[20]), .B(product[19]), .C(product[15]), .D(
        product[17]), .Y(n106) );
  or4d1_hd U375 ( .A(product[23]), .B(product[7]), .C(product[8]), .D(
        product[9]), .Y(n104) );
  scg5d1_hd U376 ( .A(n46), .B(n353), .C(n51), .D(n220), .E(n14), .F(n102), 
        .Y(guard) );
  nd2bd1_hd U377 ( .AN(N502), .B(n111), .Y(N501) );
  oa21d1_hd U378 ( .A(n37), .B(n113), .C(n114), .Y(z_m[23]) );
  ao22d1_hd U379 ( .A(n115), .B(N273), .C(n47), .D(n378), .Y(n114) );
  scg4d1_hd U380 ( .A(n115), .B(N272), .C(n47), .D(n376), .E(n284), .F(n102), 
        .G(n35), .H(n51), .Y(z_m[22]) );
  scg4d1_hd U381 ( .A(n115), .B(N271), .C(n36), .D(n102), .E(n46), .F(n375), 
        .G(n34), .H(n50), .Y(z_m[21]) );
  scg4d1_hd U382 ( .A(n115), .B(N270), .C(n46), .D(n374), .E(n35), .F(n102), 
        .G(n33), .H(n51), .Y(z_m[20]) );
  scg4d1_hd U383 ( .A(n115), .B(N269), .C(n47), .D(n373), .E(n34), .F(n102), 
        .G(n32), .H(n50), .Y(z_m[19]) );
  scg4d1_hd U384 ( .A(n115), .B(N268), .C(n46), .D(n372), .E(n33), .F(n102), 
        .G(n31), .H(n51), .Y(z_m[18]) );
  scg4d1_hd U385 ( .A(n115), .B(N267), .C(n47), .D(n371), .E(n32), .F(n102), 
        .G(n30), .H(n50), .Y(z_m[17]) );
  scg4d1_hd U386 ( .A(n115), .B(N266), .C(n46), .D(n370), .E(n31), .F(n102), 
        .G(n29), .H(n51), .Y(z_m[16]) );
  scg4d1_hd U387 ( .A(n115), .B(N265), .C(n47), .D(n369), .E(n30), .F(n102), 
        .G(n28), .H(n50), .Y(z_m[15]) );
  scg4d1_hd U388 ( .A(n115), .B(N264), .C(n46), .D(n368), .E(n29), .F(n102), 
        .G(n27), .H(n50), .Y(z_m[14]) );
  scg4d1_hd U389 ( .A(n115), .B(N263), .C(n47), .D(n367), .E(n28), .F(n102), 
        .G(n26), .H(n51), .Y(z_m[13]) );
  scg4d1_hd U390 ( .A(n115), .B(N262), .C(n46), .D(n366), .E(n27), .F(n102), 
        .G(n25), .H(n50), .Y(z_m[12]) );
  scg4d1_hd U391 ( .A(n115), .B(N261), .C(n47), .D(n365), .E(n26), .F(n102), 
        .G(n24), .H(n51), .Y(z_m[11]) );
  scg4d1_hd U392 ( .A(n115), .B(N260), .C(n46), .D(n364), .E(n25), .F(n102), 
        .G(n23), .H(n50), .Y(z_m[10]) );
  scg4d1_hd U393 ( .A(n115), .B(N259), .C(n47), .D(n363), .E(n24), .F(n102), 
        .G(n22), .H(n51), .Y(z_m[9]) );
  scg4d1_hd U394 ( .A(n115), .B(N258), .C(n46), .D(n362), .E(n23), .F(n102), 
        .G(n21), .H(n50), .Y(z_m[8]) );
  scg4d1_hd U395 ( .A(n115), .B(N257), .C(n47), .D(n361), .E(n22), .F(n102), 
        .G(n20), .H(n51), .Y(z_m[7]) );
  scg4d1_hd U396 ( .A(n115), .B(N256), .C(n46), .D(n360), .E(n21), .F(n102), 
        .G(n19), .H(n51), .Y(z_m[6]) );
  scg4d1_hd U397 ( .A(n115), .B(N255), .C(n47), .D(n359), .E(n20), .F(n102), 
        .G(n18), .H(n51), .Y(z_m[5]) );
  scg4d1_hd U398 ( .A(n115), .B(N254), .C(n46), .D(n358), .E(n19), .F(n102), 
        .G(n17), .H(n50), .Y(z_m[4]) );
  scg4d1_hd U399 ( .A(n115), .B(N253), .C(n47), .D(n357), .E(n18), .F(n102), 
        .G(n51), .H(n16), .Y(z_m[3]) );
  scg4d1_hd U400 ( .A(n115), .B(N252), .C(n46), .D(n356), .E(n17), .F(n102), 
        .G(n50), .H(n15), .Y(z_m[2]) );
  scg4d1_hd U401 ( .A(n115), .B(N251), .C(n47), .D(n355), .E(n14), .F(n50), 
        .G(n16), .H(n102), .Y(z_m[1]) );
  scg4d1_hd U402 ( .A(n115), .B(N250), .C(n46), .D(n354), .E(n48), .F(n50), 
        .G(n15), .H(n102), .Y(z_m[0]) );
  scg18d1_hd U403 ( .A(n116), .B(n117), .C(n506), .D(n112), .E(n111), .Y(N463)
         );
  nd2bd1_hd U404 ( .AN(n119), .B(n102), .Y(n112) );
  nr2d1_hd U405 ( .A(n120), .B(n121), .Y(n117) );
  nd4d1_hd U406 ( .A(n35), .B(n34), .C(n33), .D(n32), .Y(n121) );
  or4d1_hd U407 ( .A(n122), .B(n123), .C(n124), .D(n125), .Y(n120) );
  nd4d1_hd U408 ( .A(n36), .B(n284), .C(n14), .D(n15), .Y(n125) );
  nd4d1_hd U409 ( .A(n19), .B(n18), .C(n17), .D(n16), .Y(n124) );
  nd4d1_hd U410 ( .A(n23), .B(n22), .C(n21), .D(n20), .Y(n123) );
  nd4d1_hd U411 ( .A(n27), .B(n26), .C(n25), .D(n24), .Y(n122) );
  nr2d1_hd U412 ( .A(n126), .B(n110), .Y(n116) );
  oa211d1_hd U413 ( .A(n14), .B(n103), .C(n48), .D(n115), .Y(n110) );
  or2d1_hd U414 ( .A(n220), .B(n219), .Y(n103) );
  nd4d1_hd U415 ( .A(n31), .B(n30), .C(n29), .D(n28), .Y(n126) );
  ao22d1_hd U416 ( .A(n129), .B(n344), .C(n346), .D(n130), .Y(n127) );
  ivd1_hd U417 ( .A(n131), .Y(n130) );
  scg6d1_hd U418 ( .A(N292), .B(n132), .C(n503), .Y(n471) );
  scg6d1_hd U419 ( .A(n132), .B(N291), .C(n503), .Y(n472) );
  scg6d1_hd U420 ( .A(n132), .B(N290), .C(n503), .Y(n473) );
  scg6d1_hd U421 ( .A(n132), .B(N289), .C(n503), .Y(n474) );
  scg6d1_hd U422 ( .A(n132), .B(N288), .C(n503), .Y(n475) );
  scg6d1_hd U423 ( .A(n132), .B(N287), .C(n503), .Y(n476) );
  scg6d1_hd U424 ( .A(n132), .B(N286), .C(n503), .Y(n477) );
  scg6d1_hd U425 ( .A(n132), .B(n143), .C(n503), .Y(n478) );
  nr2d1_hd U426 ( .A(n137), .B(n138), .Y(n133) );
  ad4d1_hd U427 ( .A(n140), .B(n141), .C(n142), .D(n143), .Y(n139) );
  ivd1_hd U428 ( .A(n379), .Y(n143) );
  ad4d1_hd U429 ( .A(n380), .B(n387), .C(n386), .D(n118), .Y(n140) );
  ivd1_hd U430 ( .A(n284), .Y(n118) );
  oa21d1_hd U431 ( .A(n113), .B(n144), .C(n128), .Y(n479) );
  oa21d1_hd U432 ( .A(n145), .B(n146), .C(n147), .Y(n128) );
  oa22d1_hd U433 ( .A(n148), .B(n149), .C(n150), .D(n151), .Y(n146) );
  oa22d1_hd U434 ( .A(n151), .B(n153), .C(n154), .D(n148), .Y(n145) );
  ivd1_hd U435 ( .A(n36), .Y(n113) );
  nr2bd1_hd U436 ( .AN(n35), .B(n144), .Y(n480) );
  nr2bd1_hd U437 ( .AN(n34), .B(n144), .Y(n481) );
  nr2bd1_hd U438 ( .AN(n33), .B(n144), .Y(n482) );
  nr2bd1_hd U439 ( .AN(n32), .B(n144), .Y(n483) );
  nr2bd1_hd U440 ( .AN(n31), .B(n144), .Y(n484) );
  nr2bd1_hd U441 ( .AN(n30), .B(n144), .Y(n485) );
  nr2bd1_hd U442 ( .AN(n29), .B(n144), .Y(n486) );
  nr2bd1_hd U443 ( .AN(n28), .B(n144), .Y(n487) );
  nr2bd1_hd U444 ( .AN(n27), .B(n144), .Y(n488) );
  nr2bd1_hd U445 ( .AN(n26), .B(n144), .Y(n489) );
  nr2bd1_hd U446 ( .AN(n25), .B(n144), .Y(n490) );
  nr2bd1_hd U447 ( .AN(n24), .B(n144), .Y(n491) );
  nr2bd1_hd U448 ( .AN(n23), .B(n144), .Y(n492) );
  nr2bd1_hd U449 ( .AN(n22), .B(n144), .Y(n493) );
  nr2bd1_hd U450 ( .AN(n21), .B(n144), .Y(n494) );
  nr2bd1_hd U451 ( .AN(n20), .B(n144), .Y(n495) );
  nr2bd1_hd U452 ( .AN(n19), .B(n144), .Y(n496) );
  nr2bd1_hd U453 ( .AN(n18), .B(n144), .Y(n497) );
  nr2bd1_hd U454 ( .AN(n17), .B(n144), .Y(n498) );
  nr2bd1_hd U455 ( .AN(n16), .B(n144), .Y(n499) );
  nr2bd1_hd U456 ( .AN(n15), .B(n144), .Y(n500) );
  nr2bd1_hd U457 ( .AN(n14), .B(n144), .Y(n501) );
  oa21d1_hd U458 ( .A(n387), .B(n386), .C(n156), .Y(n136) );
  ivd1_hd U459 ( .A(n388), .Y(n156) );
  scg6d1_hd U460 ( .A(C76_DATA2_9), .B(n206), .C(n147), .Y(b_e[9]) );
  scg6d1_hd U461 ( .A(C76_DATA2_8), .B(n206), .C(n147), .Y(b_e[8]) );
  scg6d1_hd U462 ( .A(C76_DATA2_7), .B(n206), .C(n147), .Y(b_e[7]) );
  ad2d1_hd U463 ( .A(C76_DATA2_6), .B(n206), .Y(b_e[6]) );
  ad2d1_hd U464 ( .A(C76_DATA2_5), .B(n206), .Y(b_e[5]) );
  ad2d1_hd U465 ( .A(C76_DATA2_4), .B(n206), .Y(b_e[4]) );
  ad2d1_hd U466 ( .A(C76_DATA2_3), .B(n206), .Y(b_e[3]) );
  ad2d1_hd U467 ( .A(C76_DATA2_2), .B(n206), .Y(b_e[2]) );
  scg6d1_hd U468 ( .A(C76_DATA2_1), .B(n206), .C(n147), .Y(b_e[1]) );
  ad2d1_hd U469 ( .A(C76_DATA2_0), .B(n206), .Y(b_e[0]) );
  scg6d1_hd U470 ( .A(C72_DATA2_9), .B(C2_Z_0), .C(n147), .Y(a_e[9]) );
  scg6d1_hd U471 ( .A(C72_DATA2_8), .B(C2_Z_0), .C(n147), .Y(a_e[8]) );
  scg6d1_hd U472 ( .A(C72_DATA2_7), .B(C2_Z_0), .C(n147), .Y(a_e[7]) );
  ad2d1_hd U473 ( .A(C72_DATA2_6), .B(C2_Z_0), .Y(a_e[6]) );
  ad2d1_hd U474 ( .A(C72_DATA2_5), .B(C2_Z_0), .Y(a_e[5]) );
  ad2d1_hd U475 ( .A(C72_DATA2_4), .B(C2_Z_0), .Y(a_e[4]) );
  ad2d1_hd U476 ( .A(C72_DATA2_3), .B(C2_Z_0), .Y(a_e[3]) );
  ad2d1_hd U477 ( .A(C72_DATA2_2), .B(C2_Z_0), .Y(a_e[2]) );
  scg6d1_hd U478 ( .A(C72_DATA2_1), .B(C2_Z_0), .C(n147), .Y(a_e[1]) );
  ad2d1_hd U479 ( .A(C72_DATA2_0), .B(C2_Z_0), .Y(a_e[0]) );
  scg14d1_hd U480 ( .A(n99), .B(n256), .C(n134), .Y(b_m[23]) );
  oa21d1_hd U481 ( .A(n155), .B(n159), .C(n160), .Y(N406) );
  ivd1_hd U482 ( .A(N382), .Y(n160) );
  nr2bd1_hd U483 ( .AN(n389), .B(n157), .Y(b_m[0]) );
  scg14d1_hd U484 ( .A(n162), .B(n459), .C(n134), .Y(a_m[23]) );
  ivd1_hd U485 ( .A(n147), .Y(n134) );
  oa21d1_hd U486 ( .A(n152), .B(n159), .C(n39), .Y(N380) );
  nd3bd1_hd U487 ( .AN(n163), .B(n147), .C(n151), .Y(n159) );
  ivd1_hd U488 ( .A(n137), .Y(n151) );
  nr2bd1_hd U489 ( .AN(n420), .B(n157), .Y(a_m[0]) );
  or2d1_hd U490 ( .A(n1), .B(N430), .Y(state[3]) );
  oa21d1_hd U491 ( .A(n137), .B(n163), .C(n147), .Y(n131) );
  ivd1_hd U492 ( .A(n138), .Y(n148) );
  nr4d1_hd U493 ( .A(n265), .B(n294), .C(n264), .D(n168), .Y(n138) );
  ao22d1_hd U494 ( .A(n150), .B(n152), .C(n154), .D(n155), .Y(n167) );
  ivd1_hd U495 ( .A(n158), .Y(n155) );
  nd4d1_hd U496 ( .A(n265), .B(n294), .C(n264), .D(n169), .Y(n158) );
  ivd1_hd U497 ( .A(n168), .Y(n169) );
  nd3d1_hd U498 ( .A(n263), .B(n170), .C(n171), .Y(n168) );
  nr2d1_hd U499 ( .A(n299), .B(n296), .Y(n171) );
  nr4d1_hd U500 ( .A(n262), .B(n298), .C(n295), .D(n297), .Y(n170) );
  scg12d1_hd U501 ( .A(n172), .B(n173), .C(n174), .Y(n154) );
  nd4d1_hd U502 ( .A(n175), .B(n176), .C(n177), .D(n178), .Y(n174) );
  nr4d1_hd U503 ( .A(n228), .B(n229), .C(n456), .D(n223), .Y(n178) );
  nr4d1_hd U504 ( .A(n457), .B(n222), .C(n453), .D(n455), .Y(n177) );
  nr4d1_hd U505 ( .A(n225), .B(n255), .C(n226), .D(n224), .Y(n176) );
  nr4d1_hd U506 ( .A(n253), .B(n221), .C(n254), .D(n230), .Y(n175) );
  nr4d1_hd U507 ( .A(n452), .B(n256), .C(n287), .D(n227), .Y(n173) );
  nr4d1_hd U508 ( .A(n462), .B(n231), .C(n460), .D(n454), .Y(n172) );
  ivd1_hd U509 ( .A(n161), .Y(n152) );
  nd4d1_hd U510 ( .A(n179), .B(n288), .C(n261), .D(n260), .Y(n161) );
  ivd1_hd U511 ( .A(n180), .Y(n179) );
  scg12d1_hd U512 ( .A(n181), .B(n182), .C(n183), .Y(n150) );
  nd4d1_hd U513 ( .A(n184), .B(n185), .C(n186), .D(n187), .Y(n183) );
  nr4d1_hd U514 ( .A(n237), .B(n234), .C(n252), .D(n249), .Y(n187) );
  nr4d1_hd U515 ( .A(n232), .B(n246), .C(n238), .D(n243), .Y(n186) );
  nr4d1_hd U516 ( .A(n239), .B(n233), .C(n236), .D(n251), .Y(n185) );
  nr4d1_hd U517 ( .A(n248), .B(n245), .C(n240), .D(n242), .Y(n184) );
  nr4d1_hd U518 ( .A(n461), .B(n459), .C(n286), .D(n241), .Y(n182) );
  nr4d1_hd U519 ( .A(n235), .B(n250), .C(n247), .D(n244), .Y(n181) );
  nr4d1_hd U520 ( .A(n261), .B(n288), .C(n260), .D(n180), .Y(n137) );
  nd3d1_hd U521 ( .A(n259), .B(n188), .C(n189), .Y(n180) );
  nr2d1_hd U522 ( .A(n292), .B(n293), .Y(n189) );
  nr4d1_hd U523 ( .A(n291), .B(n290), .C(n289), .D(n258), .Y(n188) );
  ivd1_hd U524 ( .A(n129), .Y(n135) );
  oa211d1_hd U525 ( .A(n285), .B(n192), .C(n164), .D(n41), .Y(state[2]) );
  scg18d1_hd U527 ( .A(n102), .B(n119), .C(n45), .D(n194), .E(n195), .Y(N350)
         );
  nd2bd1_hd U528 ( .AN(n502), .B(N85), .Y(n195) );
  ao211d1_hd U529 ( .A(n50), .B(n284), .C(state[1]), .D(n197), .Y(n194) );
  scg17d1_hd U530 ( .A(n198), .B(n72), .C(n129), .D(n200), .Y(state[1]) );
  scg20d1_hd U531 ( .A(n72), .B(n201), .C(n115), .Y(n200) );
  nr2d1_hd U532 ( .A(n202), .B(n166), .Y(n129) );
  nr2d1_hd U533 ( .A(n191), .B(n165), .Y(N41) );
  ivd1_hd U534 ( .A(n198), .Y(n165) );
  nr2d1_hd U535 ( .A(n257), .B(n285), .Y(n198) );
  oa211d1_hd U536 ( .A(n380), .B(n204), .C(n387), .D(n386), .Y(n203) );
  nr3d1_hd U537 ( .A(n381), .B(n383), .C(n382), .Y(n141) );
  nr2d1_hd U538 ( .A(n385), .B(n384), .Y(n142) );
  or2d1_hd U539 ( .A(n190), .B(n257), .Y(n202) );
  ad2d1_hd U540 ( .A(n162), .B(n261), .Y(C1_Z_9) );
  nr2bd1_hd U541 ( .AN(n260), .B(n164), .Y(C1_Z_8) );
  ivd1_hd U542 ( .A(n162), .Y(n164) );
  fd1eqd4_hd clk_r_REG105_S5 ( .D(b_m[23]), .E(N406), .CK(n515), .Q(n452) );
  ivd1_hd U1 ( .A(i_RST), .Y(n2) );
  ivd1_hd U2 ( .A(i_RST), .Y(n3) );
  ivd1_hd U3 ( .A(i_RST), .Y(n10) );
  ivd1_hd U4 ( .A(i_RST), .Y(n11) );
  ivd1_hd U5 ( .A(i_RST), .Y(n12) );
  ivd1_hd U6 ( .A(i_RST), .Y(n13) );
  ivd6_hd U12 ( .A(n4) );
  ivd6_hd U13 ( .A(n9) );
  ivd6_hd U19 ( .A(n8) );
  ivd6_hd U20 ( .A(n6) );
  ivd6_hd U21 ( .A(n7) );
  ivd6_hd U22 ( .A(n5) );
  fds2eqd1_hd clk_r_REG201_S4 ( .CRN(n3), .D(state[2]), .E(N350), .CK(i_CLK), 
        .Q(n217) );
  fds2eqd1_hd clk_r_REG9_S3 ( .CRN(n11), .D(state[3]), .E(N350), .CK(i_CLK), 
        .Q(n285) );
  fd1eqd2_hd clk_r_REG177_S5 ( .D(a_m[23]), .E(N380), .CK(n515), .Q(n461) );
  fd1eqd1_hd clk_r_REG79_S5 ( .D(z_e[9]), .E(N463), .CK(n515), .Q(n388) );
  fd1eqd1_hd clk_r_REG78_S5 ( .D(z_e[8]), .E(N463), .CK(n515), .Q(n387) );
  fd1eqd1_hd clk_r_REG33_S5 ( .D(z_e[7]), .E(N463), .CK(n515), .Q(n386) );
  fd1eqd1_hd clk_r_REG27_S5 ( .D(z_e[1]), .E(N463), .CK(n515), .Q(n380) );
  fd1eqd1_hd clk_r_REG1_S2 ( .D(n347), .E(N45), .CK(n511), .Q(n346) );
  fd1eqd1_hd clk_r_REG84_S4 ( .D(b_e[6]), .E(N419), .CK(n512), .Q(n299) );
  fd1eqd1_hd clk_r_REG83_S4 ( .D(b_e[5]), .E(N419), .CK(n512), .Q(n298) );
  fd1eqd1_hd clk_r_REG82_S4 ( .D(b_e[4]), .E(N419), .CK(n512), .Q(n297) );
  fd1eqd1_hd clk_r_REG81_S4 ( .D(b_e[3]), .E(N419), .CK(n512), .Q(n296) );
  fd1eqd1_hd clk_r_REG80_S4 ( .D(b_e[2]), .E(N419), .CK(n512), .Q(n295) );
  fd1eqd1_hd clk_r_REG96_S4 ( .D(b_e[0]), .E(N419), .CK(n515), .Q(n294) );
  fd1eqd1_hd clk_r_REG93_S4 ( .D(a_e[6]), .E(N408), .CK(n511), .Q(n293) );
  fd1eqd1_hd clk_r_REG92_S4 ( .D(a_e[5]), .E(N408), .CK(n511), .Q(n292) );
  fd1eqd1_hd clk_r_REG91_S4 ( .D(a_e[4]), .E(N408), .CK(n511), .Q(n291) );
  fd1eqd1_hd clk_r_REG90_S4 ( .D(a_e[3]), .E(N408), .CK(n511), .Q(n290) );
  fd1eqd1_hd clk_r_REG89_S4 ( .D(a_e[2]), .E(N408), .CK(n511), .Q(n289) );
  fd1eqd1_hd clk_r_REG98_S4 ( .D(a_e[0]), .E(N408), .CK(n515), .Q(n288) );
  fd1eqd1_hd clk_r_REG107_S7 ( .D(z_m[23]), .E(N498), .CK(n515), .Q(n284) );
  fd1eqd1_hd clk_r_REG87_S4 ( .D(b_e[9]), .E(N419), .CK(n512), .Q(n265) );
  fd1eqd1_hd clk_r_REG86_S4 ( .D(b_e[8]), .E(N419), .CK(n512), .Q(n264) );
  fd1eqd1_hd clk_r_REG85_S4 ( .D(b_e[7]), .E(N419), .CK(n512), .Q(n263) );
  fd1eqd1_hd clk_r_REG10_S4 ( .D(b_e[1]), .E(N419), .CK(n515), .Q(n262) );
  fd1eqd1_hd clk_r_REG95_S2 ( .D(a_e[9]), .E(N408), .CK(n511), .Q(n261) );
  fd1eqd1_hd clk_r_REG94_S2 ( .D(a_e[8]), .E(N408), .CK(n511), .Q(n260) );
  fd1eqd1_hd clk_r_REG6_S2 ( .D(a_e[7]), .E(N408), .CK(n511), .Q(n259) );
  fd1eqd1_hd clk_r_REG88_S4 ( .D(a_e[1]), .E(N408), .CK(n515), .Q(n258) );
  fd1eqd1_hd clk_r_REG133_S33 ( .D(sticky), .E(N502), .CK(n513), .Q(n219) );
  fd1eqd1_hd clk_r_REG130_S30 ( .D(z_m[0]), .E(N498), .CK(n515), .Q(n14) );
  oa22d1_hd U8 ( .A(n133), .B(n134), .C(n135), .D(n136), .Y(n503) );
  scg2d1_hd U9 ( .A(N45), .B(n442), .C(n162), .D(n252), .Y(n504) );
  scg2d1_hd U10 ( .A(N45), .B(n403), .C(n99), .D(n229), .Y(n505) );
  fd1qd1_hd clk_r_REG0_S1 ( .D(N33), .CK(n507), .Q(n347) );
  fd1qd1_hd clk_r_REG264_S1 ( .D(i_B[0]), .CK(n507), .Q(n389) );
  fd1qd1_hd clk_r_REG263_S1 ( .D(i_B[1]), .CK(n507), .Q(n390) );
  fd1qd1_hd clk_r_REG262_S1 ( .D(i_B[2]), .CK(n507), .Q(n391) );
  fd1qd1_hd clk_r_REG261_S1 ( .D(i_B[3]), .CK(n507), .Q(n392) );
  fd1qd1_hd clk_r_REG260_S1 ( .D(i_B[4]), .CK(n507), .Q(n393) );
  fd1qd1_hd clk_r_REG259_S1 ( .D(i_B[5]), .CK(n507), .Q(n394) );
  fd1qd1_hd clk_r_REG258_S1 ( .D(i_B[6]), .CK(n507), .Q(n395) );
  fd1qd1_hd clk_r_REG257_S1 ( .D(i_B[7]), .CK(n507), .Q(n396) );
  fd1qd1_hd clk_r_REG256_S1 ( .D(i_B[8]), .CK(n507), .Q(n397) );
  fd1qd1_hd clk_r_REG255_S1 ( .D(i_B[9]), .CK(n507), .Q(n398) );
  fd1qd1_hd clk_r_REG254_S1 ( .D(i_B[10]), .CK(n507), .Q(n399) );
  fd1qd1_hd clk_r_REG253_S1 ( .D(i_B[11]), .CK(n507), .Q(n400) );
  fd1qd1_hd clk_r_REG252_S1 ( .D(i_B[12]), .CK(n507), .Q(n401) );
  fd1qd1_hd clk_r_REG251_S1 ( .D(i_B[13]), .CK(n507), .Q(n402) );
  fd1qd1_hd clk_r_REG250_S1 ( .D(i_B[14]), .CK(n507), .Q(n403) );
  fd1qd1_hd clk_r_REG249_S1 ( .D(i_B[15]), .CK(n507), .Q(n404) );
  fd1qd1_hd clk_r_REG248_S1 ( .D(i_B[16]), .CK(n507), .Q(n405) );
  fd1qd1_hd clk_r_REG247_S1 ( .D(i_B[17]), .CK(n507), .Q(n406) );
  fd1qd1_hd clk_r_REG246_S1 ( .D(i_B[18]), .CK(n507), .Q(n407) );
  fd1qd1_hd clk_r_REG245_S1 ( .D(i_B[19]), .CK(n507), .Q(n408) );
  fd1qd1_hd clk_r_REG244_S1 ( .D(i_B[20]), .CK(n507), .Q(n409) );
  fd1qd1_hd clk_r_REG243_S1 ( .D(i_B[21]), .CK(n507), .Q(n410) );
  fd1qd1_hd clk_r_REG242_S1 ( .D(i_B[22]), .CK(n507), .Q(n411) );
  fd1qd1_hd clk_r_REG241_S1 ( .D(i_B[23]), .CK(n507), .Q(n412) );
  fd1qd1_hd clk_r_REG240_S1 ( .D(i_B[24]), .CK(n507), .Q(n413) );
  fd1qd1_hd clk_r_REG239_S1 ( .D(i_B[25]), .CK(n507), .Q(n414) );
  fd1qd1_hd clk_r_REG238_S1 ( .D(i_B[26]), .CK(n507), .Q(n415) );
  fd1qd1_hd clk_r_REG237_S1 ( .D(i_B[27]), .CK(n507), .Q(n416) );
  fd1qd1_hd clk_r_REG236_S1 ( .D(i_B[28]), .CK(n507), .Q(n417) );
  fd1qd1_hd clk_r_REG235_S1 ( .D(i_B[29]), .CK(n507), .Q(n418) );
  fd1qd1_hd clk_r_REG234_S1 ( .D(i_B[30]), .CK(n507), .Q(n419) );
  fd1qd1_hd clk_r_REG233_S1 ( .D(i_A[0]), .CK(n507), .Q(n420) );
  fd1qd1_hd clk_r_REG232_S1 ( .D(i_A[1]), .CK(n507), .Q(n421) );
  fd1qd1_hd clk_r_REG231_S1 ( .D(i_A[2]), .CK(n507), .Q(n422) );
  fd1qd1_hd clk_r_REG230_S1 ( .D(i_A[3]), .CK(n507), .Q(n423) );
  fd1qd1_hd clk_r_REG229_S1 ( .D(i_A[4]), .CK(n507), .Q(n424) );
  fd1qd1_hd clk_r_REG228_S1 ( .D(i_A[5]), .CK(n507), .Q(n425) );
  fd1qd1_hd clk_r_REG227_S1 ( .D(i_A[6]), .CK(n507), .Q(n426) );
  fd1qd1_hd clk_r_REG226_S1 ( .D(i_A[7]), .CK(n507), .Q(n427) );
  fd1qd1_hd clk_r_REG225_S1 ( .D(i_A[8]), .CK(n507), .Q(n428) );
  fd1qd1_hd clk_r_REG224_S1 ( .D(i_A[9]), .CK(n507), .Q(n429) );
  fd1qd1_hd clk_r_REG223_S1 ( .D(i_A[10]), .CK(n507), .Q(n430) );
  fd1qd1_hd clk_r_REG222_S1 ( .D(i_A[11]), .CK(n507), .Q(n431) );
  fd1qd1_hd clk_r_REG221_S1 ( .D(i_A[12]), .CK(n507), .Q(n432) );
  fd1qd1_hd clk_r_REG220_S1 ( .D(i_A[13]), .CK(n507), .Q(n433) );
  fd1qd1_hd clk_r_REG219_S1 ( .D(i_A[14]), .CK(n507), .Q(n434) );
  fd1qd1_hd clk_r_REG218_S1 ( .D(i_A[15]), .CK(n507), .Q(n435) );
  fd1qd1_hd clk_r_REG217_S1 ( .D(i_A[16]), .CK(n507), .Q(n436) );
  fd1qd1_hd clk_r_REG216_S1 ( .D(i_A[17]), .CK(n507), .Q(n437) );
  fd1qd1_hd clk_r_REG215_S1 ( .D(i_A[18]), .CK(n507), .Q(n438) );
  fd1qd1_hd clk_r_REG214_S1 ( .D(i_A[19]), .CK(n507), .Q(n439) );
  fd1qd1_hd clk_r_REG213_S1 ( .D(i_A[20]), .CK(n507), .Q(n440) );
  fd1qd1_hd clk_r_REG212_S1 ( .D(i_A[21]), .CK(n507), .Q(n441) );
  fd1qd1_hd clk_r_REG211_S1 ( .D(i_A[22]), .CK(n507), .Q(n442) );
  fd1qd1_hd clk_r_REG210_S1 ( .D(i_A[23]), .CK(n507), .Q(n443) );
  fd1qd1_hd clk_r_REG209_S1 ( .D(i_A[24]), .CK(n507), .Q(n444) );
  fd1qd1_hd clk_r_REG208_S1 ( .D(i_A[25]), .CK(n507), .Q(n445) );
  fd1qd1_hd clk_r_REG207_S1 ( .D(i_A[26]), .CK(n507), .Q(n446) );
  fd1qd1_hd clk_r_REG206_S1 ( .D(i_A[27]), .CK(n507), .Q(n447) );
  fd1qd1_hd clk_r_REG205_S1 ( .D(i_A[28]), .CK(n507), .Q(n448) );
  fd1qd1_hd clk_r_REG204_S1 ( .D(i_A[29]), .CK(n507), .Q(n449) );
  fd1qd1_hd clk_r_REG5_S1 ( .D(i_A[30]), .CK(n507), .Q(n451) );
  fd1qd1_hd clk_r_REG8_S4 ( .D(n267), .CK(n508), .Q(o_Z[22]) );
  fd1qd1_hd clk_r_REG26_S6 ( .D(n269), .CK(n508), .Q(o_Z[23]) );
  fd1qd1_hd clk_r_REG24_S6 ( .D(n271), .CK(n508), .Q(o_Z[24]) );
  fd1qd1_hd clk_r_REG22_S6 ( .D(n273), .CK(n508), .Q(o_Z[25]) );
  fd1qd1_hd clk_r_REG20_S6 ( .D(n275), .CK(n508), .Q(o_Z[26]) );
  fd1qd1_hd clk_r_REG18_S6 ( .D(n277), .CK(n508), .Q(o_Z[27]) );
  fd1qd1_hd clk_r_REG16_S6 ( .D(n279), .CK(n508), .Q(o_Z[28]) );
  fd1qd1_hd clk_r_REG14_S6 ( .D(n281), .CK(n508), .Q(o_Z[29]) );
  fd1qd1_hd clk_r_REG12_S6 ( .D(n283), .CK(n508), .Q(o_Z[30]) );
  fd1qd1_hd clk_r_REG75_S7 ( .D(n303), .CK(n508), .Q(o_Z[1]) );
  fd1qd1_hd clk_r_REG73_S7 ( .D(n305), .CK(n508), .Q(o_Z[2]) );
  fd1qd1_hd clk_r_REG71_S7 ( .D(n307), .CK(n508), .Q(o_Z[3]) );
  fd1qd1_hd clk_r_REG69_S7 ( .D(n309), .CK(n508), .Q(o_Z[4]) );
  fd1qd1_hd clk_r_REG67_S7 ( .D(n311), .CK(n508), .Q(o_Z[5]) );
  fd1qd1_hd clk_r_REG65_S7 ( .D(n313), .CK(n508), .Q(o_Z[6]) );
  fd1qd1_hd clk_r_REG63_S7 ( .D(n315), .CK(n508), .Q(o_Z[7]) );
  fd1qd1_hd clk_r_REG61_S7 ( .D(n317), .CK(n508), .Q(o_Z[8]) );
  fd1qd1_hd clk_r_REG59_S7 ( .D(n319), .CK(n508), .Q(o_Z[9]) );
  fd1qd1_hd clk_r_REG57_S7 ( .D(n321), .CK(n508), .Q(o_Z[10]) );
  fd1qd1_hd clk_r_REG55_S7 ( .D(n323), .CK(n508), .Q(o_Z[11]) );
  fd1qd1_hd clk_r_REG53_S7 ( .D(n325), .CK(n508), .Q(o_Z[12]) );
  fd1qd1_hd clk_r_REG51_S7 ( .D(n327), .CK(n508), .Q(o_Z[13]) );
  fd1qd1_hd clk_r_REG49_S7 ( .D(n329), .CK(n508), .Q(o_Z[14]) );
  fd1qd1_hd clk_r_REG47_S7 ( .D(n331), .CK(n508), .Q(o_Z[15]) );
  fd1qd1_hd clk_r_REG45_S7 ( .D(n333), .CK(n508), .Q(o_Z[16]) );
  fd1qd1_hd clk_r_REG43_S7 ( .D(n335), .CK(n508), .Q(o_Z[17]) );
  fd1qd1_hd clk_r_REG41_S7 ( .D(n337), .CK(n508), .Q(o_Z[18]) );
  fd1qd1_hd clk_r_REG39_S7 ( .D(n339), .CK(n508), .Q(o_Z[19]) );
  fd1qd1_hd clk_r_REG37_S7 ( .D(n341), .CK(n508), .Q(o_Z[20]) );
  fd1qd1_hd clk_r_REG35_S7 ( .D(n343), .CK(n508), .Q(o_Z[21]) );
  fd1qd1_hd clk_r_REG4_S4 ( .D(n349), .CK(n508), .Q(o_Z[31]) );
  fd1qd1_hd clk_r_REG77_S7 ( .D(n301), .CK(n508), .Q(o_Z[0]) );
  fd1qd1_hd clk_r_REG7_S3 ( .D(n479), .CK(n509), .Q(n267) );
  fd1qd1_hd clk_r_REG25_S5 ( .D(n478), .CK(n509), .Q(n269) );
  fd1qd1_hd clk_r_REG23_S5 ( .D(n477), .CK(n509), .Q(n271) );
  fd1qd1_hd clk_r_REG21_S5 ( .D(n476), .CK(n509), .Q(n273) );
  fd1qd1_hd clk_r_REG19_S5 ( .D(n475), .CK(n509), .Q(n275) );
  fd1qd1_hd clk_r_REG17_S5 ( .D(n474), .CK(n509), .Q(n277) );
  fd1qd1_hd clk_r_REG15_S5 ( .D(n473), .CK(n509), .Q(n279) );
  fd1qd1_hd clk_r_REG13_S5 ( .D(n472), .CK(n509), .Q(n281) );
  fd1qd1_hd clk_r_REG11_S5 ( .D(n471), .CK(n509), .Q(n283) );
  fd1qd1_hd clk_r_REG76_S6 ( .D(n501), .CK(n509), .Q(n301) );
  fd1qd1_hd clk_r_REG74_S6 ( .D(n500), .CK(n509), .Q(n303) );
  fd1qd1_hd clk_r_REG72_S6 ( .D(n499), .CK(n509), .Q(n305) );
  fd1qd1_hd clk_r_REG70_S6 ( .D(n498), .CK(n509), .Q(n307) );
  fd1qd1_hd clk_r_REG68_S6 ( .D(n497), .CK(n509), .Q(n309) );
  fd1qd1_hd clk_r_REG66_S6 ( .D(n496), .CK(n509), .Q(n311) );
  fd1qd1_hd clk_r_REG64_S6 ( .D(n495), .CK(n509), .Q(n313) );
  fd1qd1_hd clk_r_REG62_S6 ( .D(n494), .CK(n509), .Q(n315) );
  fd1qd1_hd clk_r_REG60_S6 ( .D(n493), .CK(n509), .Q(n317) );
  fd1qd1_hd clk_r_REG58_S6 ( .D(n492), .CK(n509), .Q(n319) );
  fd1qd1_hd clk_r_REG56_S6 ( .D(n491), .CK(n509), .Q(n321) );
  fd1qd1_hd clk_r_REG54_S6 ( .D(n490), .CK(n509), .Q(n323) );
  fd1qd1_hd clk_r_REG52_S6 ( .D(n489), .CK(n509), .Q(n325) );
  fd1qd1_hd clk_r_REG50_S6 ( .D(n488), .CK(n509), .Q(n327) );
  fd1qd1_hd clk_r_REG48_S6 ( .D(n487), .CK(n509), .Q(n329) );
  fd1qd1_hd clk_r_REG46_S6 ( .D(n486), .CK(n509), .Q(n331) );
  fd1qd1_hd clk_r_REG44_S6 ( .D(n485), .CK(n509), .Q(n333) );
  fd1qd1_hd clk_r_REG42_S6 ( .D(n484), .CK(n509), .Q(n335) );
  fd1qd1_hd clk_r_REG40_S6 ( .D(n483), .CK(n509), .Q(n337) );
  fd1qd1_hd clk_r_REG38_S6 ( .D(n482), .CK(n509), .Q(n339) );
  fd1qd1_hd clk_r_REG36_S6 ( .D(n481), .CK(n509), .Q(n341) );
  fd1qd1_hd clk_r_REG34_S6 ( .D(n480), .CK(n509), .Q(n343) );
  fd1qd1_hd clk_r_REG3_S3 ( .D(n470), .CK(n509), .Q(n349) );
  fd1qd1_hd clk_r_REG159_S6 ( .D(n101), .CK(n510), .Q(n218) );
  fd1qd1_hd clk_r_REG2_S3 ( .D(n346), .CK(n510), .Q(n344) );
  fd1qd1_hd clk_r_REG158_S6 ( .D(product[24]), .CK(n510), .Q(n352) );
  fd1qd1_hd clk_r_REG157_S6 ( .D(product[25]), .CK(n510), .Q(n353) );
  fd1qd1_hd clk_r_REG156_S6 ( .D(product[26]), .CK(n510), .Q(n354) );
  fd1qd1_hd clk_r_REG155_S6 ( .D(product[27]), .CK(n510), .Q(n355) );
  fd1qd1_hd clk_r_REG154_S6 ( .D(product[28]), .CK(n510), .Q(n356) );
  fd1qd1_hd clk_r_REG153_S6 ( .D(product[29]), .CK(n510), .Q(n357) );
  fd1qd1_hd clk_r_REG152_S6 ( .D(product[30]), .CK(n510), .Q(n358) );
  fd1qd1_hd clk_r_REG150_S6 ( .D(product[31]), .CK(n510), .Q(n359) );
  fd1qd1_hd clk_r_REG149_S6 ( .D(product[32]), .CK(n510), .Q(n360) );
  fd1qd1_hd clk_r_REG151_S6 ( .D(product[33]), .CK(n510), .Q(n361) );
  fd1qd1_hd clk_r_REG148_S6 ( .D(product[34]), .CK(n510), .Q(n362) );
  fd1qd1_hd clk_r_REG147_S6 ( .D(product[35]), .CK(n510), .Q(n363) );
  fd1qd1_hd clk_r_REG146_S6 ( .D(product[36]), .CK(n510), .Q(n364) );
  fd1qd1_hd clk_r_REG145_S6 ( .D(product[37]), .CK(n510), .Q(n365) );
  fd1qd1_hd clk_r_REG144_S6 ( .D(product[38]), .CK(n510), .Q(n366) );
  fd1qd1_hd clk_r_REG143_S6 ( .D(product[39]), .CK(n510), .Q(n367) );
  fd1qd1_hd clk_r_REG142_S6 ( .D(product[40]), .CK(n510), .Q(n368) );
  fd1qd1_hd clk_r_REG141_S6 ( .D(product[41]), .CK(n510), .Q(n369) );
  fd1qd1_hd clk_r_REG140_S6 ( .D(product[42]), .CK(n510), .Q(n370) );
  fd1qd1_hd clk_r_REG139_S6 ( .D(product[43]), .CK(n510), .Q(n371) );
  fd1qd1_hd clk_r_REG138_S6 ( .D(product[44]), .CK(n510), .Q(n372) );
  fd1qd1_hd clk_r_REG137_S6 ( .D(product[45]), .CK(n510), .Q(n373) );
  fd1qd1_hd clk_r_REG136_S6 ( .D(product[46]), .CK(n510), .Q(n374) );
  fd1qd1_hd clk_r_REG135_S6 ( .D(product[47]), .CK(n510), .Q(n375) );
  fd1qd1_hd clk_r_REG134_S6 ( .D(product[48]), .CK(n510), .Q(n376) );
  fd1qd2_hd clk_r_REG188_S4 ( .D(a_m[10]), .CK(n511), .Q(n241) );
  fd1qd2_hd clk_r_REG187_S4 ( .D(a_m[11]), .CK(n511), .Q(n242) );
  fd1qd2_hd clk_r_REG186_S4 ( .D(a_m[12]), .CK(n511), .Q(n243) );
  fd1qd2_hd clk_r_REG185_S4 ( .D(a_m[13]), .CK(n511), .Q(n244) );
  fd1qd2_hd clk_r_REG184_S4 ( .D(a_m[14]), .CK(n511), .Q(n245) );
  fd1qd2_hd clk_r_REG183_S4 ( .D(a_m[15]), .CK(n511), .Q(n246) );
  fd1qd2_hd clk_r_REG182_S4 ( .D(a_m[16]), .CK(n511), .Q(n247) );
  fd1qd2_hd clk_r_REG181_S4 ( .D(a_m[17]), .CK(n511), .Q(n248) );
  fd1qd2_hd clk_r_REG180_S4 ( .D(a_m[18]), .CK(n511), .Q(n249) );
  fd1qd2_hd clk_r_REG179_S4 ( .D(a_m[19]), .CK(n511), .Q(n250) );
  fd1qd2_hd clk_r_REG178_S4 ( .D(a_m[20]), .CK(n511), .Q(n251) );
  fd1qd2_hd clk_r_REG175_S4 ( .D(a_m[21]), .CK(n511), .Q(n252) );
  fd1qd2_hd clk_r_REG176_S4 ( .D(n504), .CK(n511), .Q(n459) );
  fd1qd4_hd clk_r_REG197_S4 ( .D(a_m[1]), .CK(n511), .Q(n232) );
  fd1qd4_hd clk_r_REG200_S4 ( .D(a_m[0]), .CK(n511), .Q(n286) );
  fd1qd4_hd clk_r_REG169_S4 ( .D(n505), .CK(n512), .Q(n460) );
  fd1qd1_hd clk_r_REG198_S4 ( .D(b_m[1]), .CK(n512), .Q(n221) );
  fd1qd1_hd clk_r_REG173_S4 ( .D(b_m[3]), .CK(n512), .Q(n222) );
  fd1qd1_hd clk_r_REG174_S4 ( .D(b_m[4]), .CK(n512), .Q(n223) );
  fd1qd1_hd clk_r_REG161_S4 ( .D(b_m[6]), .CK(n512), .Q(n224) );
  fd1qd1_hd clk_r_REG162_S4 ( .D(b_m[7]), .CK(n512), .Q(n225) );
  fd1qd1_hd clk_r_REG164_S4 ( .D(b_m[9]), .CK(n512), .Q(n226) );
  fd1qd1_hd clk_r_REG165_S4 ( .D(b_m[10]), .CK(n512), .Q(n227) );
  fd1qd1_hd clk_r_REG167_S4 ( .D(b_m[12]), .CK(n512), .Q(n228) );
  fd1qd1_hd clk_r_REG168_S4 ( .D(b_m[13]), .CK(n512), .Q(n229) );
  fd1qd1_hd clk_r_REG170_S4 ( .D(b_m[15]), .CK(n512), .Q(n230) );
  fd1qd1_hd clk_r_REG171_S4 ( .D(b_m[16]), .CK(n512), .Q(n231) );
  fd1qd1_hd clk_r_REG100_S4 ( .D(b_m[18]), .CK(n512), .Q(n253) );
  fd1qd1_hd clk_r_REG101_S4 ( .D(b_m[19]), .CK(n512), .Q(n254) );
  fd1qd1_hd clk_r_REG103_S4 ( .D(b_m[21]), .CK(n512), .Q(n255) );
  fd1qd1_hd clk_r_REG104_S4 ( .D(b_m[22]), .CK(n512), .Q(n256) );
  fd1qd1_hd clk_r_REG199_S4 ( .D(b_m[0]), .CK(n512), .Q(n287) );
  fd1qd4_hd clk_r_REG172_S4 ( .D(b_m[2]), .CK(n512), .Q(n453) );
  fd1qd4_hd clk_r_REG166_S4 ( .D(b_m[11]), .CK(n512), .Q(n454) );
  fd1qd4_hd clk_r_REG102_S4 ( .D(b_m[20]), .CK(n512), .Q(n455) );
  fd1qd4_hd clk_r_REG163_S4 ( .D(b_m[8]), .CK(n512), .Q(n456) );
  fd1qd4_hd clk_r_REG99_S4 ( .D(b_m[17]), .CK(n512), .Q(n462) );
  fd1qd1_hd clk_r_REG129_S29 ( .D(z_m[1]), .CK(n513), .Q(n15) );
  fd1qd1_hd clk_r_REG128_S28 ( .D(z_m[2]), .CK(n513), .Q(n16) );
  fd1qd1_hd clk_r_REG127_S27 ( .D(z_m[3]), .CK(n513), .Q(n17) );
  fd1qd1_hd clk_r_REG126_S26 ( .D(z_m[4]), .CK(n513), .Q(n18) );
  fd1qd1_hd clk_r_REG125_S25 ( .D(z_m[5]), .CK(n513), .Q(n19) );
  fd1qd1_hd clk_r_REG124_S24 ( .D(z_m[6]), .CK(n513), .Q(n20) );
  fd1qd1_hd clk_r_REG123_S23 ( .D(z_m[7]), .CK(n513), .Q(n21) );
  fd1qd1_hd clk_r_REG122_S22 ( .D(z_m[8]), .CK(n513), .Q(n22) );
  fd1qd1_hd clk_r_REG121_S21 ( .D(z_m[9]), .CK(n513), .Q(n23) );
  fd1qd1_hd clk_r_REG120_S20 ( .D(z_m[10]), .CK(n513), .Q(n24) );
  fd1qd1_hd clk_r_REG119_S19 ( .D(z_m[11]), .CK(n513), .Q(n25) );
  fd1qd1_hd clk_r_REG118_S18 ( .D(z_m[12]), .CK(n513), .Q(n26) );
  fd1qd1_hd clk_r_REG117_S17 ( .D(z_m[13]), .CK(n513), .Q(n27) );
  fd1qd1_hd clk_r_REG116_S16 ( .D(z_m[14]), .CK(n513), .Q(n28) );
  fd1qd1_hd clk_r_REG115_S15 ( .D(z_m[15]), .CK(n513), .Q(n29) );
  fd1qd1_hd clk_r_REG114_S14 ( .D(z_m[16]), .CK(n513), .Q(n30) );
  fd1qd1_hd clk_r_REG113_S13 ( .D(z_m[17]), .CK(n513), .Q(n31) );
  fd1qd1_hd clk_r_REG112_S12 ( .D(z_m[18]), .CK(n513), .Q(n32) );
  fd1qd1_hd clk_r_REG111_S11 ( .D(z_m[19]), .CK(n513), .Q(n33) );
  fd1qd1_hd clk_r_REG110_S10 ( .D(z_m[20]), .CK(n513), .Q(n34) );
  fd1qd1_hd clk_r_REG109_S9 ( .D(z_m[21]), .CK(n513), .Q(n35) );
  fd1qd1_hd clk_r_REG108_S8 ( .D(z_m[22]), .CK(n513), .Q(n36) );
  fd1qd1_hd clk_r_REG97_S5 ( .D(z_e[0]), .CK(n514), .Q(n379) );
  fd1qd1_hd clk_r_REG28_S5 ( .D(z_e[2]), .CK(n514), .Q(n381) );
  fd1qd1_hd clk_r_REG29_S5 ( .D(z_e[3]), .CK(n514), .Q(n382) );
  fd1qd1_hd clk_r_REG30_S5 ( .D(z_e[4]), .CK(n514), .Q(n383) );
  fd1qd1_hd clk_r_REG31_S5 ( .D(z_e[5]), .CK(n514), .Q(n384) );
  fd1qd1_hd clk_r_REG32_S5 ( .D(z_e[6]), .CK(n514), .Q(n385) );
  fd1eqd1_hd clk_r_REG202_S4 ( .D(n522), .E(n544), .CK(i_CLK), .Q(n72) );
  fd1eqd1_hd clk_r_REG203_S4 ( .D(n520), .E(n546), .CK(i_CLK), .Q(n257) );
  fd1eqd1_hd clk_r_REG265_S1 ( .D(n518), .E(n548), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1eqd1_hd clk_r_REG266_S1 ( .D(n516), .E(n550), .CK(i_CLK), .Q(o_Z_STB) );
  fd1eqd1_hd clk_r_REG132_S32 ( .D(round_bit), .E(N501), .CK(n513), .Q(n220)
         );
  fd1eqd1_hd clk_r_REG131_S31 ( .D(guard), .E(N501), .CK(n513), .Q(n48) );
  float_multiplier_DW01_inc_0 add_x_3 ( .A({n284, n36, n35, n34, n33, n32, n31, 
        n30, n29, n28, n27, n26, n25, n24, n23, n22, n21, n20, n19, n18, n17, 
        n16, n15, n14}), .SUM({N273, N272, N271, N270, N269, N268, N267, N266, 
        N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, 
        N253, N252, N251, N250}) );
  float_multiplier_DP_OP_114_130_61_0 DP_OP_114_130_61 ( .I1({n261, n260, n259, 
        n293, n292, n291, n290, n289, n258, n288}), .I2({n265, n264, n263, 
        n299, n298, n297, n296, n295, n262, n294}), .I3(n506), .I4({n388, n387, 
        n386, n385, n384, n383, n382, n381, n380, n379}), .I5(n1), .I6(n49), 
        .O1(z_e) );
  float_multiplier_DW_mult_uns_2 mult_x_1 ( .a({n461, n459, n252, n251, n250, 
        n249, n248, n247, n246, n245, n244, n243, n242, n241, n240, n239, n238, 
        n237, n236, n235, n234, n233, n232, n286}), .b({n452, n256, n255, n455, 
        n254, n253, n462, n231, n230, n460, n229, n228, n454, n227, n226, n456, 
        n225, n224, n457, n223, n222, n453, n221, n287}), .product(product) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_14 clk_gate_clk_r_REG98_S4_0 ( .CLK(
        i_CLK), .EN(n552), .ENCLK(n515), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_15 clk_gate_clk_r_REG97_S5_0 ( .CLK(
        i_CLK), .EN(N463), .ENCLK(n514), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_16 clk_gate_clk_r_REG131_S31_0 ( .CLK(
        i_CLK), .EN(N498), .ENCLK(n513), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_17 clk_gate_clk_r_REG169_S4_0 ( .CLK(
        i_CLK), .EN(N382), .ENCLK(n512), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_18 clk_gate_clk_r_REG188_S4_0 ( .CLK(
        i_CLK), .EN(n458), .ENCLK(n511), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_19 clk_gate_clk_r_REG159_S6_0 ( .CLK(
        i_CLK), .EN(n506), .ENCLK(n510), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_20 clk_gate_clk_r_REG7_S3_0 ( .CLK(
        i_CLK), .EN(N430), .ENCLK(n509), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_21 clk_gate_clk_r_REG8_S4_0 ( .CLK(
        i_CLK), .EN(N85), .ENCLK(n508), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_float_multiplier_22 clk_gate_clk_r_REG0_S1_0 ( .CLK(
        i_CLK), .EN(n45), .ENCLK(n507), .TE(1'b0) );
  fd1qd1_hd clk_r_REG106_S6 ( .D(product[49]), .CK(n510), .Q(n378) );
  fd1qd2_hd clk_r_REG196_S4 ( .D(a_m[2]), .CK(n511), .Q(n233) );
  fd1qd2_hd clk_r_REG195_S4 ( .D(a_m[3]), .CK(n511), .Q(n234) );
  fd1qd2_hd clk_r_REG194_S4 ( .D(a_m[4]), .CK(n511), .Q(n235) );
  fd1qd2_hd clk_r_REG193_S4 ( .D(a_m[5]), .CK(n511), .Q(n236) );
  fd1qd2_hd clk_r_REG192_S4 ( .D(a_m[6]), .CK(n511), .Q(n237) );
  fd1qd2_hd clk_r_REG191_S4 ( .D(a_m[7]), .CK(n511), .Q(n238) );
  fd1qd2_hd clk_r_REG190_S4 ( .D(a_m[8]), .CK(n511), .Q(n239) );
  fd1qd2_hd clk_r_REG189_S4 ( .D(a_m[9]), .CK(n511), .Q(n240) );
  fd1qd2_hd clk_r_REG160_S4 ( .D(b_m[5]), .CK(n512), .Q(n457) );
  clknd2d1_hd U7 ( .A(n217), .B(n257), .Y(n541) );
  clknd2d1_hd U23 ( .A(n285), .B(n502), .Y(n529) );
  clknd2d1_hd U24 ( .A(n100), .B(n157), .Y(n206) );
  nr2d1_hd U25 ( .A(n196), .B(n166), .Y(N85) );
  clknd2d1_hd U26 ( .A(n135), .B(n131), .Y(N430) );
  ivd1_hd U27 ( .A(n39), .Y(n458) );
  oa21d1_hd U28 ( .A(n452), .B(n100), .C(n157), .Y(N382) );
  mx2d1_hd U29 ( .D0(n190), .D1(n165), .S(n542), .Y(n552) );
  ivd1_hd U30 ( .A(n517), .Y(n516) );
  clknd2d1_hd U31 ( .A(n13), .B(n549), .Y(n517) );
  ivd1_hd U32 ( .A(n519), .Y(n518) );
  clknd2d1_hd U33 ( .A(n12), .B(n547), .Y(n519) );
  ivd1_hd U34 ( .A(n521), .Y(n520) );
  clknd2d1_hd U35 ( .A(n10), .B(n545), .Y(n521) );
  clknd2d1_hd U36 ( .A(n530), .B(n2), .Y(n544) );
  ivd1_hd U37 ( .A(n523), .Y(n522) );
  clknd2d1_hd U38 ( .A(n2), .B(n543), .Y(n523) );
  nd2bd1_hd U39 ( .AN(N501), .B(n110), .Y(N498) );
  nr2ad1_hd U40 ( .A(n201), .B(n192), .Y(n506) );
  ivd1_hd U41 ( .A(n40), .Y(n45) );
  ao21d1_hd U42 ( .A(n524), .B(n525), .C(n526), .Y(n543) );
  ivd1_hd U43 ( .A(n2), .Y(n526) );
  nd3d1_hd U44 ( .A(n72), .B(n217), .C(n527), .Y(n525) );
  nr2d1_hd U45 ( .A(n284), .B(n285), .Y(n527) );
  ao22d1_hd U46 ( .A(n190), .B(n536), .C(n205), .D(n528), .Y(n524) );
  oa211d1_hd U47 ( .A(n285), .B(n461), .C(n72), .D(n529), .Y(n528) );
  scg14d1_hd U48 ( .A(n285), .B(n217), .C(n257), .Y(n530) );
  ad2d1_hd U49 ( .A(n10), .B(n531), .Y(n545) );
  oa22d1_hd U50 ( .A(n45), .B(n532), .C(n257), .D(n533), .Y(n531) );
  ao211d1_hd U51 ( .A(n72), .B(n190), .C(n534), .D(n535), .Y(n533) );
  ao21d1_hd U52 ( .A(n536), .B(n537), .C(n217), .Y(n535) );
  oa21d1_hd U53 ( .A(n45), .B(n119), .C(n285), .Y(n537) );
  ivd1_hd U54 ( .A(n72), .Y(n536) );
  nr3d1_hd U55 ( .A(n538), .B(n285), .C(n72), .Y(n534) );
  ao21d1_hd U56 ( .A(n199), .B(n452), .C(n45), .Y(n538) );
  oa211d1_hd U57 ( .A(n285), .B(n539), .C(n540), .D(n72), .Y(n532) );
  scg16d1_hd U58 ( .A(n502), .B(n217), .C(n285), .Y(n540) );
  oa22d1_hd U59 ( .A(n284), .B(n541), .C(n461), .D(n217), .Y(n539) );
  nd4d1_hd U60 ( .A(n285), .B(n217), .C(n10), .D(n40), .Y(n546) );
  ad2d1_hd U61 ( .A(n469), .B(n12), .Y(n547) );
  nd2bd1_hd U62 ( .AN(N41), .B(n12), .Y(n548) );
  ad2d1_hd U63 ( .A(n502), .B(n13), .Y(n549) );
  nd2bd1_hd U64 ( .AN(N85), .B(n13), .Y(n550) );
  nr2d1_hd U65 ( .A(n217), .B(n72), .Y(n542) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_lpf_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_lpf_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_lpf_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_lpf_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module iir_lpf ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   w_rstn, w_rst, r_add_AB_STB, w_add_AB_ACK, w_add_Z_STB, r_add_Z_ACK,
         w_mult_1_AB_ACK, w_mult_2_AB_ACK, w_mult_AB_ACK, w_mult_1_Z_STB,
         w_mult_2_Z_STB, w_mult_Z_STB, r_mult_AB_STB, r_mult_Z_ACK, N27, N28,
         N29, N35, N39, N40, N41, N46, N111, N435, N440, N561, N564, N766,
         N768, N769, N770, N771, N772, N773, N774, N775, N776, N777, N778,
         N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789,
         N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, N802,
         N804, N806, N812, N813, N814, N817, N818, alt20_n15, alt20_n16, n163,
         n164, n165, n167, n170, n171, n173, n175, n176, n177, n178, n179,
         n180, n183, n184, n185, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n254, n255, n287, n289, n292, n355, n577, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n978, n979, n980, n981, n982, n1000, n172, n186, n579, n596,
         n598, n599, n602, n603, n616, n631, n632, n633, n634, n636, n665,
         n666, n668, n732, n733, n792, n857, n858, n859, n864, n915, n1002,
         n1116, n1338, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1607;
  wire   [31:0] r_add_A;
  wire   [31:0] r_add_B;
  wire   [31:0] w_add_Z;
  wire   [29:0] r_mult_1_A;
  wire   [31:0] r_mult_1_B;
  wire   [31:0] w_mult_1_Z;
  wire   [29:0] r_mult_2_A;
  wire   [31:0] r_mult_2_B;
  wire   [31:0] w_mult_2_Z;
  wire   [95:0] r_x_data;
  wire   [63:0] r_y_data;
  wire   [1:0] r_pstate;
  wire   [1:0] r_counter;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  float_adder add ( .i_A(r_add_A), .i_B(r_add_B), .i_AB_STB(r_add_AB_STB), 
        .o_AB_ACK(w_add_AB_ACK), .o_Z(w_add_Z), .o_Z_STB(w_add_Z_STB), 
        .i_Z_ACK(r_add_Z_ACK), .i_CLK(i_CLK), .i_RST(n577) );
  float_multiplier mult_1 ( .i_A({1'b0, 1'b0, r_mult_1_A[29:26], n1376, n1376, 
        r_mult_1_A[23:22], 1'b0, r_mult_1_A[20:19], 1'b0, r_mult_1_A[17:16], 
        n1376, n1376, 1'b0, n1376, r_mult_1_A[11:10], n1375, n1376, 
        r_mult_1_A[7:5], n1375, r_mult_1_A[3:0]}), .i_B(r_mult_1_B), 
        .i_AB_STB(r_mult_AB_STB), .o_AB_ACK(w_mult_1_AB_ACK), .o_Z(w_mult_1_Z), 
        .o_Z_STB(w_mult_1_Z_STB), .i_Z_ACK(r_mult_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(n577) );
  float_multiplier mult_2 ( .i_A({n1375, 1'b0, r_mult_2_A[29:26], n1375, n1375, 
        1'b0, r_mult_2_A[22], n1376, r_mult_2_A[20:19], 1'b0, 
        r_mult_2_A[17:16], 1'b0, n1376, n1376, 1'b0, r_mult_2_A[11:10], 1'b0, 
        n1376, r_mult_2_A[7:5], n1376, r_mult_2_A[3:0]}), .i_B(r_mult_2_B), 
        .i_AB_STB(r_mult_AB_STB), .o_AB_ACK(w_mult_2_AB_ACK), .o_Z(w_mult_2_Z), 
        .o_Z_STB(w_mult_2_Z_STB), .i_Z_ACK(r_mult_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(w_rst) );
  ao211d1_hd U188 ( .A(n173), .B(n165), .C(n179), .D(N561), .Y(n177) );
  oa21d1_hd U193 ( .A(N435), .B(n962), .C(n171), .Y(n184) );
  ivd1_hd U194 ( .A(n966), .Y(n171) );
  oa21d1_hd U195 ( .A(n965), .B(N440), .C(w_add_Z_STB), .Y(n183) );
  ivd1_hd U200 ( .A(n967), .Y(n164) );
  oa22d1_hd U205 ( .A(n966), .B(n167), .C(n173), .D(n178), .Y(n188) );
  ivd1_hd U206 ( .A(w_add_Z_STB), .Y(n173) );
  oa22d1_hd U207 ( .A(n167), .B(n189), .C(n178), .D(n190), .Y(N799) );
  oa22d1_hd U208 ( .A(n167), .B(n191), .C(n178), .D(n192), .Y(N798) );
  oa22d1_hd U209 ( .A(n167), .B(n193), .C(n178), .D(n194), .Y(N797) );
  oa22d1_hd U210 ( .A(n167), .B(n195), .C(n178), .D(n196), .Y(N796) );
  oa22d1_hd U211 ( .A(n167), .B(n197), .C(n178), .D(n198), .Y(N795) );
  oa22d1_hd U212 ( .A(n167), .B(n199), .C(n178), .D(n200), .Y(N794) );
  oa22d1_hd U213 ( .A(n167), .B(n201), .C(n178), .D(n202), .Y(N793) );
  oa22d1_hd U214 ( .A(n167), .B(n203), .C(n178), .D(n204), .Y(N792) );
  oa22d1_hd U215 ( .A(n167), .B(n205), .C(n178), .D(n206), .Y(N791) );
  oa22d1_hd U216 ( .A(n167), .B(n207), .C(n178), .D(n208), .Y(N790) );
  oa22d1_hd U217 ( .A(n167), .B(n209), .C(n178), .D(n210), .Y(N789) );
  oa22d1_hd U218 ( .A(n167), .B(n211), .C(n178), .D(n212), .Y(N788) );
  oa22d1_hd U219 ( .A(n167), .B(n213), .C(n178), .D(n214), .Y(N787) );
  oa22d1_hd U220 ( .A(n167), .B(n215), .C(n178), .D(n216), .Y(N786) );
  oa22d1_hd U221 ( .A(n167), .B(n217), .C(n178), .D(n218), .Y(N785) );
  oa22d1_hd U222 ( .A(n167), .B(n219), .C(n178), .D(n220), .Y(N784) );
  oa22d1_hd U223 ( .A(n167), .B(n221), .C(n178), .D(n222), .Y(N783) );
  oa22d1_hd U224 ( .A(n167), .B(n223), .C(n178), .D(n224), .Y(N782) );
  oa22d1_hd U225 ( .A(n167), .B(n225), .C(n178), .D(n226), .Y(N781) );
  oa22d1_hd U226 ( .A(n167), .B(n227), .C(n178), .D(n228), .Y(N780) );
  oa22d1_hd U227 ( .A(n167), .B(n229), .C(n178), .D(n230), .Y(N779) );
  oa22d1_hd U228 ( .A(n167), .B(n231), .C(n178), .D(n232), .Y(N778) );
  oa22d1_hd U229 ( .A(n167), .B(n233), .C(n178), .D(n234), .Y(N777) );
  oa22d1_hd U230 ( .A(n167), .B(n235), .C(n178), .D(n236), .Y(N776) );
  oa22d1_hd U231 ( .A(n167), .B(n237), .C(n178), .D(n238), .Y(N775) );
  oa22d1_hd U232 ( .A(n167), .B(n239), .C(n178), .D(n240), .Y(N774) );
  oa22d1_hd U233 ( .A(n167), .B(n241), .C(n178), .D(n242), .Y(N773) );
  oa22d1_hd U234 ( .A(n167), .B(n243), .C(n178), .D(n244), .Y(N772) );
  oa22d1_hd U235 ( .A(n167), .B(n245), .C(n178), .D(n246), .Y(N771) );
  oa22d1_hd U236 ( .A(n167), .B(n247), .C(n178), .D(n248), .Y(N770) );
  oa22d1_hd U237 ( .A(n167), .B(n249), .C(n178), .D(n250), .Y(N769) );
  oa22d1_hd U238 ( .A(n167), .B(n251), .C(n178), .D(n252), .Y(N768) );
  nr2bd1_hd U240 ( .AN(N111), .B(n164), .Y(N766) );
  ivd1_hd U243 ( .A(w_add_Z[31]), .Y(n190) );
  ivd1_hd U246 ( .A(w_add_Z[30]), .Y(n192) );
  ivd1_hd U249 ( .A(w_add_Z[29]), .Y(n194) );
  ivd1_hd U252 ( .A(w_add_Z[28]), .Y(n196) );
  ivd1_hd U255 ( .A(w_add_Z[27]), .Y(n198) );
  ivd1_hd U258 ( .A(w_add_Z[26]), .Y(n200) );
  ivd1_hd U261 ( .A(w_add_Z[25]), .Y(n202) );
  ivd1_hd U264 ( .A(w_add_Z[24]), .Y(n204) );
  ivd1_hd U267 ( .A(w_add_Z[23]), .Y(n206) );
  ivd1_hd U270 ( .A(w_add_Z[22]), .Y(n208) );
  ivd1_hd U273 ( .A(w_add_Z[21]), .Y(n210) );
  ivd1_hd U276 ( .A(w_add_Z[20]), .Y(n212) );
  ivd1_hd U279 ( .A(w_add_Z[19]), .Y(n214) );
  ivd1_hd U282 ( .A(w_add_Z[18]), .Y(n216) );
  ivd1_hd U285 ( .A(w_add_Z[17]), .Y(n218) );
  ivd1_hd U288 ( .A(w_add_Z[16]), .Y(n220) );
  ivd1_hd U291 ( .A(w_add_Z[15]), .Y(n222) );
  ivd1_hd U294 ( .A(w_add_Z[14]), .Y(n224) );
  ivd1_hd U297 ( .A(w_add_Z[13]), .Y(n226) );
  ivd1_hd U300 ( .A(w_add_Z[12]), .Y(n228) );
  ivd1_hd U303 ( .A(w_add_Z[11]), .Y(n230) );
  ivd1_hd U306 ( .A(w_add_Z[10]), .Y(n232) );
  ivd1_hd U309 ( .A(w_add_Z[9]), .Y(n234) );
  ivd1_hd U312 ( .A(w_add_Z[8]), .Y(n236) );
  ivd1_hd U315 ( .A(w_add_Z[7]), .Y(n238) );
  ivd1_hd U318 ( .A(w_add_Z[6]), .Y(n240) );
  ivd1_hd U321 ( .A(w_add_Z[5]), .Y(n242) );
  ivd1_hd U324 ( .A(w_add_Z[4]), .Y(n244) );
  ivd1_hd U327 ( .A(w_add_Z[3]), .Y(n246) );
  ivd1_hd U330 ( .A(w_add_Z[2]), .Y(n248) );
  ivd1_hd U333 ( .A(w_add_Z[1]), .Y(n250) );
  ivd1_hd U336 ( .A(w_add_Z[0]), .Y(n252) );
  ivd1_hd U460 ( .A(w_mult_1_Z[31]), .Y(n189) );
  ivd1_hd U464 ( .A(w_mult_1_Z[30]), .Y(n191) );
  ivd1_hd U468 ( .A(w_mult_1_Z[29]), .Y(n193) );
  ivd1_hd U472 ( .A(w_mult_1_Z[28]), .Y(n195) );
  ivd1_hd U476 ( .A(w_mult_1_Z[27]), .Y(n197) );
  ivd1_hd U480 ( .A(w_mult_1_Z[26]), .Y(n199) );
  ivd1_hd U484 ( .A(w_mult_1_Z[25]), .Y(n201) );
  ivd1_hd U488 ( .A(w_mult_1_Z[24]), .Y(n203) );
  ivd1_hd U492 ( .A(w_mult_1_Z[23]), .Y(n205) );
  ivd1_hd U496 ( .A(w_mult_1_Z[22]), .Y(n207) );
  ivd1_hd U500 ( .A(w_mult_1_Z[21]), .Y(n209) );
  ivd1_hd U504 ( .A(w_mult_1_Z[20]), .Y(n211) );
  ivd1_hd U508 ( .A(w_mult_1_Z[19]), .Y(n213) );
  ivd1_hd U512 ( .A(w_mult_1_Z[18]), .Y(n215) );
  ivd1_hd U516 ( .A(w_mult_1_Z[17]), .Y(n217) );
  ivd1_hd U520 ( .A(w_mult_1_Z[16]), .Y(n219) );
  ivd1_hd U524 ( .A(w_mult_1_Z[15]), .Y(n221) );
  ivd1_hd U528 ( .A(w_mult_1_Z[14]), .Y(n223) );
  ivd1_hd U532 ( .A(w_mult_1_Z[13]), .Y(n225) );
  ivd1_hd U536 ( .A(w_mult_1_Z[12]), .Y(n227) );
  ivd1_hd U540 ( .A(w_mult_1_Z[11]), .Y(n229) );
  ivd1_hd U544 ( .A(w_mult_1_Z[10]), .Y(n231) );
  ivd1_hd U548 ( .A(w_mult_1_Z[9]), .Y(n233) );
  ivd1_hd U552 ( .A(w_mult_1_Z[8]), .Y(n235) );
  ivd1_hd U556 ( .A(w_mult_1_Z[7]), .Y(n237) );
  ivd1_hd U560 ( .A(w_mult_1_Z[6]), .Y(n239) );
  ivd1_hd U564 ( .A(w_mult_1_Z[5]), .Y(n241) );
  ivd1_hd U568 ( .A(w_mult_1_Z[4]), .Y(n243) );
  ivd1_hd U572 ( .A(w_mult_1_Z[3]), .Y(n245) );
  ivd1_hd U576 ( .A(w_mult_1_Z[2]), .Y(n247) );
  ivd1_hd U580 ( .A(w_mult_1_Z[1]), .Y(n249) );
  scg20d1_hd U583 ( .A(n969), .B(N818), .C(n164), .Y(n255) );
  ad2d1_hd U584 ( .A(n179), .B(N41), .Y(n254) );
  nr2d1_hd U585 ( .A(n969), .B(n164), .Y(n179) );
  ivd1_hd U589 ( .A(w_mult_1_Z[0]), .Y(n251) );
  nr2d1_hd U591 ( .A(n355), .B(r_counter[0]), .Y(N564) );
  nr2d1_hd U592 ( .A(n165), .B(n175), .Y(n355) );
  ad2d1_hd U598 ( .A(alt20_n16), .B(n968), .Y(N561) );
  clknd2d3_hd U820 ( .A(n964), .B(N440), .Y(n178) );
  ad2d1_hd U821 ( .A(N39), .B(N40), .Y(N435) );
  or3d1_hd U822 ( .A(n963), .B(n971), .C(N46), .Y(N818) );
  nr2d1_hd U824 ( .A(n966), .B(n167), .Y(n973) );
  ad2d1_hd U825 ( .A(r_pstate[1]), .B(r_pstate[0]), .Y(alt20_n16) );
  ivd1_hd U827 ( .A(alt20_n16), .Y(alt20_n15) );
  ad2d1_hd U828 ( .A(N39), .B(N40), .Y(N41) );
  oa21d1_hd U829 ( .A(n969), .B(n164), .C(n185), .Y(N802) );
  clknd2d1_hd U830 ( .A(w_mult_AB_ACK), .B(w_add_AB_ACK), .Y(n969) );
  ad2d1_hd U831 ( .A(w_mult_1_AB_ACK), .B(w_mult_2_AB_ACK), .Y(w_mult_AB_ACK)
         );
  clknd2d1_hd U832 ( .A(n964), .B(n1000), .Y(n163) );
  clknd2d1_hd U833 ( .A(n183), .B(n184), .Y(n1000) );
  ad2d1_hd U834 ( .A(N27), .B(N28), .Y(N29) );
  ad2d1_hd U835 ( .A(w_mult_1_Z_STB), .B(w_mult_2_Z_STB), .Y(w_mult_Z_STB) );
  clknd2d1_hd U836 ( .A(n170), .B(n167), .Y(n175) );
  clknd2d1_hd U837 ( .A(n163), .B(n180), .Y(N806) );
  ivd1_hd U1180 ( .A(n972), .Y(N812) );
  or2d1_hd U1182 ( .A(N29), .B(alt20_n16), .Y(N804) );
  or2d1_hd U1217 ( .A(N41), .B(n963), .Y(N111) );
  clknd2d1_hd U1219 ( .A(n163), .B(n164), .Y(N813) );
  ad2d1_hd U1222 ( .A(N29), .B(n616), .Y(N814) );
  clknd2d1_hd U1223 ( .A(n177), .B(n178), .Y(n176) );
  ad2d1_hd U1231 ( .A(r_counter[1]), .B(r_counter[0]), .Y(N46) );
  ivd1_hd U1232 ( .A(r_counter[0]), .Y(N40) );
  nr2d1_hd U1234 ( .A(n1374), .B(n973), .Y(n972) );
  clknd2d4_hd U1239 ( .A(n964), .B(n962), .Y(n167) );
  ivd1_hd U1622 ( .A(r_pstate[0]), .Y(N28) );
  nid3_hd U1625 ( .A(n254), .Y(n978) );
  scg6d1_hd U1628 ( .A(n175), .B(n966), .C(n176), .Y(n961) );
  ad2d1_hd U1630 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(N35) );
  nid2_hd U1635 ( .A(n980), .Y(n979) );
  nr2d1_hd U1636 ( .A(r_counter[1]), .B(N40), .Y(n963) );
  nr2d4_hd U1644 ( .A(N27), .B(r_pstate[0]), .Y(n964) );
  clknd2d1_hd U1646 ( .A(w_add_Z_STB), .B(w_mult_Z_STB), .Y(n966) );
  nr2d1_hd U1647 ( .A(r_pstate[1]), .B(N28), .Y(n967) );
  clknd2d1_hd U1648 ( .A(o_Y_DATA_VALID), .B(i_Y_ACK), .Y(n968) );
  scg8d1_hd U1649 ( .A(n179), .B(n963), .C(alt20_n16), .D(n188), .Y(n970) );
  ad2d1_hd U1655 ( .A(r_counter[1]), .B(r_counter[0]), .Y(N440) );
  nid1_hd U1656 ( .A(n254), .Y(n981) );
  nid2_hd U1657 ( .A(n981), .Y(n980) );
  nr2d1_hd U1658 ( .A(N39), .B(r_counter[0]), .Y(n971) );
  ivd1_hd U1659 ( .A(N29), .Y(n180) );
  ivd1_hd U6 ( .A(n1002), .Y(n172) );
  ivd1_hd U9 ( .A(n1002), .Y(n186) );
  ivd1_hd U11 ( .A(n1002), .Y(n579) );
  ivd1_hd U28 ( .A(n1116), .Y(n596) );
  ivd1_hd U30 ( .A(n1116), .Y(n598) );
  ivd1_hd U31 ( .A(n1338), .Y(n599) );
  ivd1_hd U34 ( .A(n1338), .Y(n602) );
  ivd1_hd U35 ( .A(n1116), .Y(n603) );
  ivd1_hd U48 ( .A(n1338), .Y(n616) );
  ivd1_hd U63 ( .A(n1002), .Y(n631) );
  ivd1_hd U64 ( .A(n1002), .Y(n632) );
  ivd1_hd U65 ( .A(n1338), .Y(n633) );
  ivd1_hd U66 ( .A(n1116), .Y(n634) );
  ivd1_hd U68 ( .A(n1116), .Y(n636) );
  ivd1_hd U97 ( .A(n1002), .Y(n665) );
  ivd1_hd U98 ( .A(n1002), .Y(n666) );
  ivd1_hd U100 ( .A(n1338), .Y(n668) );
  ivd1_hd U164 ( .A(n1116), .Y(n732) );
  ivd1_hd U165 ( .A(n1116), .Y(n733) );
  ivd1_hd U613 ( .A(n1338), .Y(n792) );
  ivd1_hd U678 ( .A(n1002), .Y(n857) );
  ivd1_hd U679 ( .A(n1116), .Y(n858) );
  ivd1_hd U680 ( .A(n1116), .Y(n859) );
  ivd1_hd U685 ( .A(n1002), .Y(n864) );
  ivd1_hd U736 ( .A(n1338), .Y(n915) );
  ivd1_hd U784 ( .A(w_rstn), .Y(n1002) );
  ivd1_hd U1322 ( .A(w_rstn), .Y(n1116) );
  ivd1_hd U1544 ( .A(w_rstn), .Y(n1338) );
  SNPS_CLOCK_GATE_HIGH_iir_lpf_12 clk_gate_o_Y_DATA_reg_31__0 ( .CLK(i_CLK), 
        .EN(N817), .ENCLK(n1380), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_lpf_13 clk_gate_r_add_B_reg_31__0 ( .CLK(i_CLK), 
        .EN(n1536), .ENCLK(n1379), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_lpf_14 clk_gate_r_mult_2_B_reg_31__0 ( .CLK(i_CLK), 
        .EN(n1607), .ENCLK(n1378), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_lpf_15 clk_gate_r_y_data_reg_63__0 ( .CLK(i_CLK), 
        .EN(N35), .ENCLK(n1377), .TE(1'b0) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n982), .E(N814), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_pstate_reg_1_ ( .D(n961), .CK(i_CLK), .RN(n599), .Q(r_pstate[1])
         );
  fd2qd1_hd r_counter_reg_1_ ( .D(n1385), .CK(i_CLK), .RN(n915), .Q(
        r_counter[1]) );
  fd2qd1_hd r_x_data_reg_65_ ( .D(r_x_data[33]), .CK(n1377), .RN(n579), .Q(
        r_x_data[65]) );
  fd2qd1_hd r_y_data_reg_0_ ( .D(o_Y_DATA[0]), .CK(n1377), .RN(n668), .Q(
        r_y_data[0]) );
  fd2qd1_hd r_y_data_reg_60_ ( .D(r_y_data[28]), .CK(n1377), .RN(n636), .Q(
        r_y_data[60]) );
  fd2qd1_hd r_y_data_reg_34_ ( .D(r_y_data[2]), .CK(n1377), .RN(n633), .Q(
        r_y_data[34]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(o_Y_DATA[27]), .CK(n1377), .RN(n668), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_x_data_reg_73_ ( .D(r_x_data[41]), .CK(n1377), .RN(n636), .Q(
        r_x_data[73]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(o_Y_DATA[29]), .CK(n1377), .RN(n596), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(o_Y_DATA[20]), .CK(n1377), .RN(n631), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_61_ ( .D(r_y_data[29]), .CK(n1377), .RN(n636), .Q(
        r_y_data[61]) );
  fd2qd1_hd r_y_data_reg_57_ ( .D(r_y_data[25]), .CK(n1377), .RN(n636), .Q(
        r_y_data[57]) );
  fd2qd1_hd r_y_data_reg_59_ ( .D(r_y_data[27]), .CK(n1377), .RN(n732), .Q(
        r_y_data[59]) );
  fd2qd1_hd r_y_data_reg_41_ ( .D(r_y_data[9]), .CK(n1377), .RN(n631), .Q(
        r_y_data[41]) );
  fd2qd1_hd r_y_data_reg_40_ ( .D(r_y_data[8]), .CK(n1377), .RN(n792), .Q(
        r_y_data[40]) );
  fd2qd1_hd r_y_data_reg_39_ ( .D(r_y_data[7]), .CK(n1377), .RN(n857), .Q(
        r_y_data[39]) );
  fd2qd1_hd r_y_data_reg_38_ ( .D(r_y_data[6]), .CK(n1377), .RN(n859), .Q(
        r_y_data[38]) );
  fd2qd1_hd r_y_data_reg_37_ ( .D(r_y_data[5]), .CK(n1377), .RN(n858), .Q(
        r_y_data[37]) );
  fd2qd1_hd r_y_data_reg_35_ ( .D(r_y_data[3]), .CK(n1377), .RN(n666), .Q(
        r_y_data[35]) );
  fd2qd1_hd r_y_data_reg_32_ ( .D(r_y_data[0]), .CK(n1377), .RN(n857), .Q(
        r_y_data[32]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(o_Y_DATA[26]), .CK(n1377), .RN(n599), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(o_Y_DATA[9]), .CK(n1377), .RN(n864), .Q(
        r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(o_Y_DATA[8]), .CK(n1377), .RN(n733), .Q(
        r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(o_Y_DATA[7]), .CK(n1377), .RN(n598), .Q(
        r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(o_Y_DATA[6]), .CK(n1377), .RN(n858), .Q(
        r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(o_Y_DATA[5]), .CK(n1377), .RN(n864), .Q(
        r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(o_Y_DATA[4]), .CK(n1377), .RN(n859), .Q(
        r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_1_ ( .D(o_Y_DATA[1]), .CK(n1377), .RN(n665), .Q(
        r_y_data[1]) );
  fd2qd1_hd r_x_data_reg_71_ ( .D(r_x_data[39]), .CK(n1377), .RN(n596), .Q(
        r_x_data[71]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(r_x_data[10]), .CK(n1377), .RN(n792), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(o_Y_DATA[30]), .CK(n1377), .RN(n792), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_x_data_reg_95_ ( .D(r_x_data[63]), .CK(n1377), .RN(n864), .Q(
        r_x_data[95]) );
  fd2qd1_hd r_x_data_reg_94_ ( .D(r_x_data[62]), .CK(n1377), .RN(n733), .Q(
        r_x_data[94]) );
  fd2qd1_hd r_x_data_reg_69_ ( .D(r_x_data[37]), .CK(n1377), .RN(n859), .Q(
        r_x_data[69]) );
  fd2qd1_hd r_x_data_reg_64_ ( .D(r_x_data[32]), .CK(n1377), .RN(n858), .Q(
        r_x_data[64]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(r_x_data[31]), .CK(n1377), .RN(n792), .Q(
        r_x_data[63]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(r_x_data[30]), .CK(n1377), .RN(n792), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(r_x_data[29]), .CK(n1377), .RN(n634), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(r_x_data[7]), .CK(n1377), .RN(n603), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(r_x_data[4]), .CK(n1377), .RN(n668), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_y_data_reg_56_ ( .D(r_y_data[24]), .CK(n1377), .RN(n616), .Q(
        r_y_data[56]) );
  fd2qd1_hd r_y_data_reg_55_ ( .D(r_y_data[23]), .CK(n1377), .RN(n732), .Q(
        r_y_data[55]) );
  fd2qd1_hd r_y_data_reg_54_ ( .D(r_y_data[22]), .CK(n1377), .RN(n733), .Q(
        r_y_data[54]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(o_Y_DATA[3]), .CK(n1377), .RN(n665), .Q(
        r_y_data[3]) );
  fd2qd1_hd r_x_data_reg_72_ ( .D(r_x_data[40]), .CK(n1377), .RN(n732), .Q(
        r_x_data[72]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(r_x_data[8]), .CK(n1377), .RN(n733), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(r_x_data[5]), .CK(n1377), .RN(n857), .Q(
        r_x_data[37]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(r_x_data[1]), .CK(n1377), .RN(n172), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_y_data_reg_63_ ( .D(r_y_data[31]), .CK(n1377), .RN(n864), .Q(
        r_y_data[63]) );
  fd2qd1_hd r_y_data_reg_62_ ( .D(r_y_data[30]), .CK(n1377), .RN(n632), .Q(
        r_y_data[62]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(o_Y_DATA[24]), .CK(n1377), .RN(n602), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(o_Y_DATA[23]), .CK(n1377), .RN(n632), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(o_Y_DATA[22]), .CK(n1377), .RN(n859), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(o_Y_DATA[21]), .CK(n1377), .RN(n596), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_52_ ( .D(r_y_data[20]), .CK(n1377), .RN(n732), .Q(
        r_y_data[52]) );
  fd2qd1_hd r_x_data_reg_79_ ( .D(r_x_data[47]), .CK(n1377), .RN(n668), .Q(
        r_x_data[79]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(o_Y_DATA[28]), .CK(n1377), .RN(n792), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_x_data_reg_93_ ( .D(r_x_data[61]), .CK(n1377), .RN(n634), .Q(
        r_x_data[93]) );
  fd2qd1_hd r_x_data_reg_92_ ( .D(r_x_data[60]), .CK(n1377), .RN(n631), .Q(
        r_x_data[92]) );
  fd2qd1_hd r_x_data_reg_91_ ( .D(r_x_data[59]), .CK(n1377), .RN(n599), .Q(
        r_x_data[91]) );
  fd2qd1_hd r_x_data_reg_90_ ( .D(r_x_data[58]), .CK(n1377), .RN(n632), .Q(
        r_x_data[90]) );
  fd2qd1_hd r_x_data_reg_89_ ( .D(r_x_data[57]), .CK(n1377), .RN(n864), .Q(
        r_x_data[89]) );
  fd2qd1_hd r_x_data_reg_88_ ( .D(r_x_data[56]), .CK(n1377), .RN(n732), .Q(
        r_x_data[88]) );
  fd2qd1_hd r_x_data_reg_86_ ( .D(r_x_data[54]), .CK(n1377), .RN(n732), .Q(
        r_x_data[86]) );
  fd2qd1_hd r_x_data_reg_85_ ( .D(r_x_data[53]), .CK(n1377), .RN(n915), .Q(
        r_x_data[85]) );
  fd2qd1_hd r_x_data_reg_84_ ( .D(r_x_data[52]), .CK(n1377), .RN(n634), .Q(
        r_x_data[84]) );
  fd2qd1_hd r_x_data_reg_83_ ( .D(r_x_data[51]), .CK(n1377), .RN(n859), .Q(
        r_x_data[83]) );
  fd2qd1_hd r_x_data_reg_82_ ( .D(r_x_data[50]), .CK(n1377), .RN(n603), .Q(
        r_x_data[82]) );
  fd2qd1_hd r_x_data_reg_81_ ( .D(r_x_data[49]), .CK(n1377), .RN(n634), .Q(
        r_x_data[81]) );
  fd2qd1_hd r_x_data_reg_78_ ( .D(r_x_data[46]), .CK(n1377), .RN(n915), .Q(
        r_x_data[78]) );
  fd2qd1_hd r_x_data_reg_77_ ( .D(r_x_data[45]), .CK(n1377), .RN(n857), .Q(
        r_x_data[77]) );
  fd2qd1_hd r_x_data_reg_76_ ( .D(r_x_data[44]), .CK(n1377), .RN(n732), .Q(
        r_x_data[76]) );
  fd2qd1_hd r_x_data_reg_75_ ( .D(r_x_data[43]), .CK(n1377), .RN(n666), .Q(
        r_x_data[75]) );
  fd2qd1_hd r_x_data_reg_74_ ( .D(r_x_data[42]), .CK(n1377), .RN(n858), .Q(
        r_x_data[74]) );
  fd2qd1_hd r_x_data_reg_68_ ( .D(r_x_data[36]), .CK(n1377), .RN(n616), .Q(
        r_x_data[68]) );
  fd2qd1_hd r_x_data_reg_67_ ( .D(r_x_data[35]), .CK(n1377), .RN(n631), .Q(
        r_x_data[67]) );
  fd2qd1_hd r_x_data_reg_66_ ( .D(r_x_data[34]), .CK(n1377), .RN(n858), .Q(
        r_x_data[66]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(r_x_data[28]), .CK(n1377), .RN(n858), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(r_x_data[27]), .CK(n1377), .RN(n631), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(r_x_data[26]), .CK(n1377), .RN(n733), .Q(
        r_x_data[58]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(r_x_data[25]), .CK(n1377), .RN(n598), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(r_x_data[24]), .CK(n1377), .RN(n599), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(r_x_data[23]), .CK(n1377), .RN(n859), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(r_x_data[22]), .CK(n1377), .RN(n616), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(r_x_data[21]), .CK(n1377), .RN(n603), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(r_x_data[20]), .CK(n1377), .RN(n666), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(r_x_data[19]), .CK(n1377), .RN(n602), .Q(
        r_x_data[51]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(r_x_data[18]), .CK(n1377), .RN(n857), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(r_x_data[17]), .CK(n1377), .RN(n915), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(r_x_data[16]), .CK(n1377), .RN(n631), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(r_x_data[15]), .CK(n1377), .RN(n632), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(r_x_data[14]), .CK(n1377), .RN(n633), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(r_x_data[13]), .CK(n1377), .RN(n602), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(r_x_data[12]), .CK(n1377), .RN(n733), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(r_x_data[11]), .CK(n1377), .RN(n915), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(r_x_data[3]), .CK(n1377), .RN(n603), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(r_x_data[2]), .CK(n1377), .RN(n668), .Q(
        r_x_data[34]) );
  fd2qd1_hd r_x_data_reg_32_ ( .D(r_x_data[0]), .CK(n1377), .RN(n172), .Q(
        r_x_data[32]) );
  fd2qd1_hd r_y_data_reg_51_ ( .D(r_y_data[19]), .CK(n1377), .RN(n857), .Q(
        r_y_data[51]) );
  fd2qd1_hd r_y_data_reg_50_ ( .D(r_y_data[18]), .CK(n1377), .RN(n579), .Q(
        r_y_data[50]) );
  fd2qd1_hd r_y_data_reg_49_ ( .D(r_y_data[17]), .CK(n1377), .RN(n186), .Q(
        r_y_data[49]) );
  fd2qd1_hd r_y_data_reg_43_ ( .D(r_y_data[11]), .CK(n1377), .RN(n633), .Q(
        r_y_data[43]) );
  fd2qd1_hd r_y_data_reg_42_ ( .D(r_y_data[10]), .CK(n1377), .RN(n579), .Q(
        r_y_data[42]) );
  fd2qd1_hd r_y_data_reg_36_ ( .D(r_y_data[4]), .CK(n1377), .RN(n186), .Q(
        r_y_data[36]) );
  fd2qd1_hd r_y_data_reg_33_ ( .D(r_y_data[1]), .CK(n1377), .RN(n579), .Q(
        r_y_data[33]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(o_Y_DATA[31]), .CK(n1377), .RN(n186), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(o_Y_DATA[25]), .CK(n1377), .RN(n632), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(o_Y_DATA[17]), .CK(n1377), .RN(n631), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(o_Y_DATA[16]), .CK(n1377), .RN(n915), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(o_Y_DATA[15]), .CK(n1377), .RN(n599), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(o_Y_DATA[14]), .CK(n1377), .RN(n579), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(o_Y_DATA[13]), .CK(n1377), .RN(n633), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(o_Y_DATA[12]), .CK(n1377), .RN(n186), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(o_Y_DATA[11]), .CK(n1377), .RN(n579), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_x_data_reg_87_ ( .D(r_x_data[55]), .CK(n1377), .RN(n172), .Q(
        r_x_data[87]) );
  fd2qd1_hd r_x_data_reg_80_ ( .D(r_x_data[48]), .CK(n1377), .RN(n186), .Q(
        r_x_data[80]) );
  fd2qd1_hd r_x_data_reg_70_ ( .D(r_x_data[38]), .CK(n1377), .RN(n665), .Q(
        r_x_data[70]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(r_x_data[9]), .CK(n1377), .RN(n596), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_y_data_reg_58_ ( .D(r_y_data[26]), .CK(n1377), .RN(n732), .Q(
        r_y_data[58]) );
  fd2qd1_hd r_y_data_reg_53_ ( .D(r_y_data[21]), .CK(n1377), .RN(n857), .Q(
        r_y_data[53]) );
  fd2qd1_hd r_y_data_reg_48_ ( .D(r_y_data[16]), .CK(n1377), .RN(n857), .Q(
        r_y_data[48]) );
  fd2qd1_hd r_y_data_reg_47_ ( .D(r_y_data[15]), .CK(n1377), .RN(n665), .Q(
        r_y_data[47]) );
  fd2qd1_hd r_y_data_reg_46_ ( .D(r_y_data[14]), .CK(n1377), .RN(n915), .Q(
        r_y_data[46]) );
  fd2qd1_hd r_y_data_reg_45_ ( .D(r_y_data[13]), .CK(n1377), .RN(n596), .Q(
        r_y_data[45]) );
  fd2qd1_hd r_y_data_reg_44_ ( .D(r_y_data[12]), .CK(n1377), .RN(n596), .Q(
        r_y_data[44]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(o_Y_DATA[19]), .CK(n1377), .RN(n668), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(o_Y_DATA[18]), .CK(n1377), .RN(n598), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(o_Y_DATA[10]), .CK(n1377), .RN(n632), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_2_ ( .D(o_Y_DATA[2]), .CK(n1377), .RN(n668), .Q(
        r_y_data[2]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(r_x_data[6]), .CK(n1377), .RN(n859), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_mult_2_A_reg_22_ ( .D(n1537), .CK(n1378), .RN(n186), .Q(
        r_mult_2_A[22]) );
  fd2qd1_hd r_mult_2_A_reg_19_ ( .D(n1538), .CK(n1378), .RN(n186), .Q(
        r_mult_2_A[19]) );
  fd2qd1_hd r_mult_2_A_reg_2_ ( .D(n1539), .CK(n1378), .RN(n186), .Q(
        r_mult_2_A[2]) );
  fd2qd1_hd r_mult_2_A_reg_1_ ( .D(n1539), .CK(n1378), .RN(n732), .Q(
        r_mult_2_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_19_ ( .D(n1538), .CK(n1378), .RN(n733), .Q(
        r_mult_1_A[19]) );
  fd2qd1_hd r_mult_1_A_reg_16_ ( .D(n1537), .CK(n1378), .RN(n858), .Q(
        r_mult_1_A[16]) );
  fd2qd1_hd r_mult_1_A_reg_2_ ( .D(n1539), .CK(n1378), .RN(n666), .Q(
        r_mult_1_A[2]) );
  fd2qd1_hd r_mult_1_A_reg_1_ ( .D(n1538), .CK(n1378), .RN(n666), .Q(
        r_mult_1_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_0_ ( .D(n1537), .CK(n1378), .RN(w_rstn), .Q(
        r_mult_1_A[0]) );
  fd2qd1_hd r_mult_1_B_reg_30_ ( .D(n1572), .CK(n1378), .RN(n666), .Q(
        r_mult_1_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_28_ ( .D(n1570), .CK(n1378), .RN(n668), .Q(
        r_mult_1_B[28]) );
  fd2qd1_hd r_mult_1_B_reg_25_ ( .D(n1567), .CK(n1378), .RN(n602), .Q(
        r_mult_1_B[25]) );
  fd2qd1_hd r_mult_1_B_reg_24_ ( .D(n1566), .CK(n1378), .RN(n598), .Q(
        r_mult_1_B[24]) );
  fd2qd1_hd r_mult_1_B_reg_22_ ( .D(n1564), .CK(n1378), .RN(n634), .Q(
        r_mult_1_B[22]) );
  fd2qd1_hd r_mult_1_B_reg_21_ ( .D(n1563), .CK(n1378), .RN(n616), .Q(
        r_mult_1_B[21]) );
  fd2qd1_hd r_mult_1_B_reg_20_ ( .D(n1562), .CK(n1378), .RN(n579), .Q(
        r_mult_1_B[20]) );
  fd2qd1_hd r_mult_1_B_reg_19_ ( .D(n1561), .CK(n1378), .RN(n186), .Q(
        r_mult_1_B[19]) );
  fd2qd1_hd r_mult_1_B_reg_18_ ( .D(n1560), .CK(n1378), .RN(n665), .Q(
        r_mult_1_B[18]) );
  fd2qd1_hd r_mult_1_B_reg_15_ ( .D(n1557), .CK(n1378), .RN(n602), .Q(
        r_mult_1_B[15]) );
  fd2qd1_hd r_mult_1_B_reg_13_ ( .D(n1555), .CK(n1378), .RN(n666), .Q(
        r_mult_1_B[13]) );
  fd2qd1_hd r_mult_1_B_reg_9_ ( .D(n1551), .CK(n1378), .RN(n172), .Q(
        r_mult_1_B[9]) );
  fd2qd1_hd r_mult_1_B_reg_7_ ( .D(n1549), .CK(n1378), .RN(n616), .Q(
        r_mult_1_B[7]) );
  fd2qd1_hd r_mult_1_B_reg_3_ ( .D(n1545), .CK(n1378), .RN(n602), .Q(
        r_mult_1_B[3]) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(i_X_DATA[31]), .CK(n1377), .RN(n668), .Q(
        r_x_data[31]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(i_X_DATA[30]), .CK(n1377), .RN(n632), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(i_X_DATA[29]), .CK(n1377), .RN(n616), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(i_X_DATA[28]), .CK(n1377), .RN(n631), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(i_X_DATA[27]), .CK(n1377), .RN(n859), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(i_X_DATA[26]), .CK(n1377), .RN(n665), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(i_X_DATA[25]), .CK(n1377), .RN(n732), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(i_X_DATA[24]), .CK(n1377), .RN(n631), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(i_X_DATA[23]), .CK(n1377), .RN(n632), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(i_X_DATA[22]), .CK(n1377), .RN(n665), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(i_X_DATA[21]), .CK(n1377), .RN(n666), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(i_X_DATA[20]), .CK(n1377), .RN(n859), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(i_X_DATA[19]), .CK(n1377), .RN(n599), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(i_X_DATA[18]), .CK(n1377), .RN(n668), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(i_X_DATA[17]), .CK(n1377), .RN(n732), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(i_X_DATA[16]), .CK(n1377), .RN(n172), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(i_X_DATA[15]), .CK(n1377), .RN(n665), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(i_X_DATA[14]), .CK(n1377), .RN(n634), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(i_X_DATA[13]), .CK(n1377), .RN(n864), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(i_X_DATA[12]), .CK(n1377), .RN(n603), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(i_X_DATA[11]), .CK(n1377), .RN(n599), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(i_X_DATA[10]), .CK(n1377), .RN(n602), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(i_X_DATA[9]), .CK(n1377), .RN(n859), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(i_X_DATA[8]), .CK(n1377), .RN(n633), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(i_X_DATA[7]), .CK(n1377), .RN(n603), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(i_X_DATA[6]), .CK(n1377), .RN(n172), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(i_X_DATA[5]), .CK(n1377), .RN(n634), .Q(
        r_x_data[5]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(i_X_DATA[4]), .CK(n1377), .RN(n579), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(i_X_DATA[3]), .CK(n1377), .RN(n636), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(i_X_DATA[2]), .CK(n1377), .RN(w_rstn), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(i_X_DATA[1]), .CK(n1377), .RN(n666), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(i_X_DATA[0]), .CK(n1377), .RN(n859), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_add_B_reg_1_ ( .D(n1504), .CK(n1379), .RN(n915), .Q(r_add_B[1])
         );
  fd2qd1_hd r_mult_AB_STB_reg ( .D(n1381), .CK(i_CLK), .RN(n858), .Q(
        r_mult_AB_STB) );
  fd2qd1_hd r_add_AB_STB_reg ( .D(n1382), .CK(i_CLK), .RN(n596), .Q(
        r_add_AB_STB) );
  fd2qd1_hd r_mult_2_B_reg_31_ ( .D(n1605), .CK(n1378), .RN(n633), .Q(
        r_mult_2_B[31]) );
  fd2qd1_hd R_1 ( .D(n980), .CK(n1378), .RN(n598), .Q(n1376) );
  fd2qd1_hd r_mult_1_B_reg_31_ ( .D(n1573), .CK(n1378), .RN(n665), .Q(
        r_mult_1_B[31]) );
  fd2qd1_hd r_mult_1_B_reg_29_ ( .D(n1571), .CK(n1378), .RN(n602), .Q(
        r_mult_1_B[29]) );
  fd2qd1_hd r_mult_1_B_reg_27_ ( .D(n1569), .CK(n1378), .RN(n864), .Q(
        r_mult_1_B[27]) );
  fd2qd1_hd r_mult_1_B_reg_26_ ( .D(n1568), .CK(n1378), .RN(n596), .Q(
        r_mult_1_B[26]) );
  fd2qd1_hd r_mult_1_B_reg_23_ ( .D(n1565), .CK(n1378), .RN(n598), .Q(
        r_mult_1_B[23]) );
  fd2qd1_hd r_mult_1_B_reg_17_ ( .D(n1559), .CK(n1378), .RN(n579), .Q(
        r_mult_1_B[17]) );
  fd2qd1_hd r_mult_1_B_reg_11_ ( .D(n1553), .CK(n1378), .RN(n792), .Q(
        r_mult_1_B[11]) );
  fd2qd1_hd r_mult_1_B_reg_5_ ( .D(n1547), .CK(n1378), .RN(n633), .Q(
        r_mult_1_B[5]) );
  fd2qd1_hd r_mult_1_B_reg_1_ ( .D(n1543), .CK(n1378), .RN(n666), .Q(
        r_mult_1_B[1]) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n1388), .CK(i_CLK), .RN(n633), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_add_B_reg_31_ ( .D(n1534), .CK(n1379), .RN(n636), .Q(r_add_B[31]) );
  fd2qd1_hd r_add_B_reg_28_ ( .D(n1531), .CK(n1379), .RN(n616), .Q(r_add_B[28]) );
  fd2qd1_hd r_add_B_reg_24_ ( .D(n1527), .CK(n1379), .RN(n634), .Q(r_add_B[24]) );
  fd2qd1_hd r_add_B_reg_23_ ( .D(n1526), .CK(n1379), .RN(n633), .Q(r_add_B[23]) );
  fd2qd1_hd r_add_B_reg_21_ ( .D(n1524), .CK(n1379), .RN(n858), .Q(r_add_B[21]) );
  fd2qd1_hd r_add_B_reg_20_ ( .D(n1523), .CK(n1379), .RN(n632), .Q(r_add_B[20]) );
  fd2qd1_hd r_add_B_reg_19_ ( .D(n1522), .CK(n1379), .RN(n733), .Q(r_add_B[19]) );
  fd2qd1_hd r_add_B_reg_18_ ( .D(n1521), .CK(n1379), .RN(n732), .Q(r_add_B[18]) );
  fd2qd1_hd r_add_B_reg_17_ ( .D(n1520), .CK(n1379), .RN(n634), .Q(r_add_B[17]) );
  fd2qd1_hd r_add_B_reg_15_ ( .D(n1518), .CK(n1379), .RN(n596), .Q(r_add_B[15]) );
  fd2qd1_hd r_add_B_reg_13_ ( .D(n1516), .CK(n1379), .RN(n596), .Q(r_add_B[13]) );
  fd2qd1_hd r_add_B_reg_11_ ( .D(n1514), .CK(n1379), .RN(n598), .Q(r_add_B[11]) );
  fd2qd1_hd r_add_B_reg_9_ ( .D(n1512), .CK(n1379), .RN(n579), .Q(r_add_B[9])
         );
  fd2qd1_hd r_add_B_reg_8_ ( .D(n1511), .CK(n1379), .RN(n636), .Q(r_add_B[8])
         );
  fd2qd1_hd r_add_B_reg_7_ ( .D(n1510), .CK(n1379), .RN(n666), .Q(r_add_B[7])
         );
  fd2qd1_hd r_add_B_reg_5_ ( .D(n1508), .CK(n1379), .RN(n858), .Q(r_add_B[5])
         );
  fd2qd1_hd r_add_B_reg_3_ ( .D(n1506), .CK(n1379), .RN(n857), .Q(r_add_B[3])
         );
  fd2qd1_hd r_add_Z_ACK_reg ( .D(n1387), .CK(i_CLK), .RN(n864), .Q(r_add_Z_ACK) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(N799), .CK(n1380), .RN(n598), .Q(
        o_Y_DATA[31]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(N798), .CK(n1380), .RN(n172), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(N797), .CK(n1380), .RN(n596), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(N796), .CK(n1380), .RN(n186), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(N795), .CK(n1380), .RN(n186), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(N794), .CK(n1380), .RN(n579), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(N793), .CK(n1380), .RN(n579), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(N792), .CK(n1380), .RN(n599), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(N791), .CK(n1380), .RN(n859), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(N790), .CK(n1380), .RN(n666), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(N789), .CK(n1380), .RN(n603), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(N788), .CK(n1380), .RN(n633), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(N787), .CK(n1380), .RN(n634), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(N786), .CK(n1380), .RN(n915), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(N785), .CK(n1380), .RN(n666), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(N784), .CK(n1380), .RN(n186), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(N783), .CK(n1380), .RN(n864), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(N782), .CK(n1380), .RN(n186), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(N781), .CK(n1380), .RN(n792), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(N780), .CK(n1380), .RN(n636), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(N779), .CK(n1380), .RN(n631), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(N778), .CK(n1380), .RN(n172), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(N777), .CK(n1380), .RN(n602), .Q(o_Y_DATA[9])
         );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(N776), .CK(n1380), .RN(n596), .Q(o_Y_DATA[8])
         );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(N775), .CK(n1380), .RN(n636), .Q(o_Y_DATA[7])
         );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(N774), .CK(n1380), .RN(n598), .Q(o_Y_DATA[6])
         );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(N773), .CK(n1380), .RN(n599), .Q(o_Y_DATA[5])
         );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(N772), .CK(n1380), .RN(n733), .Q(o_Y_DATA[4])
         );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(N771), .CK(n1380), .RN(n579), .Q(o_Y_DATA[3])
         );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(N770), .CK(n1380), .RN(n602), .Q(o_Y_DATA[2])
         );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(N769), .CK(n1380), .RN(n603), .Q(o_Y_DATA[1])
         );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(N768), .CK(n1380), .RN(n598), .Q(o_Y_DATA[0])
         );
  fd2qd1_hd R_2 ( .D(n979), .CK(n1378), .RN(n596), .Q(n1375) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(n1383), .CK(i_CLK), .RN(n858), .Q(r_pstate[0]) );
  fd2qd1_hd r_mult_1_B_reg_16_ ( .D(n1558), .CK(n1378), .RN(n186), .Q(
        r_mult_1_B[16]) );
  fd2qd1_hd r_mult_1_B_reg_14_ ( .D(n1556), .CK(n1378), .RN(n632), .Q(
        r_mult_1_B[14]) );
  fd2qd1_hd r_mult_1_B_reg_12_ ( .D(n1554), .CK(n1378), .RN(n599), .Q(
        r_mult_1_B[12]) );
  fd2qd1_hd r_mult_1_B_reg_10_ ( .D(n1552), .CK(n1378), .RN(n172), .Q(
        r_mult_1_B[10]) );
  fd2qd1_hd r_mult_1_B_reg_8_ ( .D(n1550), .CK(n1378), .RN(n732), .Q(
        r_mult_1_B[8]) );
  fd2qd1_hd r_mult_1_B_reg_6_ ( .D(n1548), .CK(n1378), .RN(n857), .Q(
        r_mult_1_B[6]) );
  fd2qd1_hd r_mult_1_B_reg_4_ ( .D(n1546), .CK(n1378), .RN(n859), .Q(
        r_mult_1_B[4]) );
  fd2qd1_hd r_mult_1_B_reg_2_ ( .D(n1544), .CK(n1378), .RN(n631), .Q(
        r_mult_1_B[2]) );
  fd2qd1_hd r_mult_1_B_reg_0_ ( .D(n1542), .CK(n1378), .RN(n599), .Q(
        r_mult_1_B[0]) );
  fd2qd1_hd r_mult_2_B_reg_30_ ( .D(n1604), .CK(n1378), .RN(n633), .Q(
        r_mult_2_B[30]) );
  fd2qd1_hd r_mult_2_B_reg_29_ ( .D(n1603), .CK(n1378), .RN(n859), .Q(
        r_mult_2_B[29]) );
  fd2qd1_hd r_mult_2_B_reg_28_ ( .D(n1602), .CK(n1378), .RN(n915), .Q(
        r_mult_2_B[28]) );
  fd2qd1_hd r_mult_2_B_reg_27_ ( .D(n1601), .CK(n1378), .RN(n733), .Q(
        r_mult_2_B[27]) );
  fd2qd1_hd r_mult_2_B_reg_26_ ( .D(n1600), .CK(n1378), .RN(n186), .Q(
        r_mult_2_B[26]) );
  fd2qd1_hd r_mult_2_B_reg_25_ ( .D(n1599), .CK(n1378), .RN(n668), .Q(
        r_mult_2_B[25]) );
  fd2qd1_hd r_mult_2_B_reg_24_ ( .D(n1598), .CK(n1378), .RN(n915), .Q(
        r_mult_2_B[24]) );
  fd2qd1_hd r_mult_2_B_reg_23_ ( .D(n1597), .CK(n1378), .RN(n915), .Q(
        r_mult_2_B[23]) );
  fd2qd1_hd r_mult_2_B_reg_22_ ( .D(n1596), .CK(n1378), .RN(n616), .Q(
        r_mult_2_B[22]) );
  fd2qd1_hd r_mult_2_B_reg_21_ ( .D(n1595), .CK(n1378), .RN(n633), .Q(
        r_mult_2_B[21]) );
  fd2qd1_hd r_mult_2_B_reg_20_ ( .D(n1594), .CK(n1378), .RN(n857), .Q(
        r_mult_2_B[20]) );
  fd2qd1_hd r_mult_2_B_reg_19_ ( .D(n1593), .CK(n1378), .RN(n602), .Q(
        r_mult_2_B[19]) );
  fd2qd1_hd r_mult_2_B_reg_18_ ( .D(n1592), .CK(n1378), .RN(n864), .Q(
        r_mult_2_B[18]) );
  fd2qd1_hd r_mult_2_B_reg_17_ ( .D(n1591), .CK(n1378), .RN(n733), .Q(
        r_mult_2_B[17]) );
  fd2qd1_hd r_mult_2_B_reg_16_ ( .D(n1590), .CK(n1378), .RN(n633), .Q(
        r_mult_2_B[16]) );
  fd2qd1_hd r_mult_2_B_reg_15_ ( .D(n1589), .CK(n1378), .RN(n665), .Q(
        r_mult_2_B[15]) );
  fd2qd1_hd r_mult_2_B_reg_14_ ( .D(n1588), .CK(n1378), .RN(n579), .Q(
        r_mult_2_B[14]) );
  fd2qd1_hd r_mult_2_B_reg_13_ ( .D(n1587), .CK(n1378), .RN(n579), .Q(
        r_mult_2_B[13]) );
  fd2qd1_hd r_mult_2_B_reg_12_ ( .D(n1586), .CK(n1378), .RN(n172), .Q(
        r_mult_2_B[12]) );
  fd2qd1_hd r_mult_2_B_reg_11_ ( .D(n1585), .CK(n1378), .RN(n602), .Q(
        r_mult_2_B[11]) );
  fd2qd1_hd r_mult_2_B_reg_10_ ( .D(n1584), .CK(n1378), .RN(n864), .Q(
        r_mult_2_B[10]) );
  fd2qd1_hd r_mult_2_B_reg_9_ ( .D(n1583), .CK(n1378), .RN(n665), .Q(
        r_mult_2_B[9]) );
  fd2qd1_hd r_mult_2_B_reg_8_ ( .D(n1582), .CK(n1378), .RN(n733), .Q(
        r_mult_2_B[8]) );
  fd2qd1_hd r_mult_2_B_reg_7_ ( .D(n1581), .CK(n1378), .RN(n631), .Q(
        r_mult_2_B[7]) );
  fd2qd1_hd r_mult_2_B_reg_6_ ( .D(n1580), .CK(n1378), .RN(n632), .Q(
        r_mult_2_B[6]) );
  fd2qd1_hd r_mult_2_B_reg_5_ ( .D(n1579), .CK(n1378), .RN(n633), .Q(
        r_mult_2_B[5]) );
  fd2qd1_hd r_mult_2_B_reg_4_ ( .D(n1578), .CK(n1378), .RN(n634), .Q(
        r_mult_2_B[4]) );
  fd2qd1_hd r_mult_2_B_reg_3_ ( .D(n1577), .CK(n1378), .RN(n915), .Q(
        r_mult_2_B[3]) );
  fd2qd1_hd r_mult_2_B_reg_2_ ( .D(n1576), .CK(n1378), .RN(n636), .Q(
        r_mult_2_B[2]) );
  fd2qd1_hd r_mult_2_B_reg_1_ ( .D(n1575), .CK(n1378), .RN(n668), .Q(
        r_mult_2_B[1]) );
  fd2qd1_hd r_mult_2_B_reg_0_ ( .D(n1574), .CK(n1378), .RN(n599), .Q(
        r_mult_2_B[0]) );
  fd2qd1_hd r_add_B_reg_30_ ( .D(n1533), .CK(n1379), .RN(n634), .Q(r_add_B[30]) );
  fd2qd1_hd r_add_B_reg_29_ ( .D(n1532), .CK(n1379), .RN(w_rstn), .Q(
        r_add_B[29]) );
  fd2qd1_hd r_add_B_reg_27_ ( .D(n1530), .CK(n1379), .RN(n636), .Q(r_add_B[27]) );
  fd2qd1_hd r_add_B_reg_26_ ( .D(n1529), .CK(n1379), .RN(n864), .Q(r_add_B[26]) );
  fd2qd1_hd r_add_B_reg_25_ ( .D(n1528), .CK(n1379), .RN(n636), .Q(r_add_B[25]) );
  fd2qd1_hd r_add_B_reg_22_ ( .D(n1525), .CK(n1379), .RN(n857), .Q(r_add_B[22]) );
  fd2qd1_hd r_add_B_reg_16_ ( .D(n1519), .CK(n1379), .RN(n603), .Q(r_add_B[16]) );
  fd2qd1_hd r_add_B_reg_14_ ( .D(n1517), .CK(n1379), .RN(n915), .Q(r_add_B[14]) );
  fd2qd1_hd r_add_B_reg_12_ ( .D(n1515), .CK(n1379), .RN(n616), .Q(r_add_B[12]) );
  fd2qd1_hd r_add_B_reg_10_ ( .D(n1513), .CK(n1379), .RN(n598), .Q(r_add_B[10]) );
  fd2qd1_hd r_add_B_reg_6_ ( .D(n1509), .CK(n1379), .RN(n599), .Q(r_add_B[6])
         );
  fd2qd1_hd r_add_B_reg_4_ ( .D(n1507), .CK(n1379), .RN(n792), .Q(r_add_B[4])
         );
  fd2qd1_hd r_add_B_reg_2_ ( .D(n1505), .CK(n1379), .RN(n172), .Q(r_add_B[2])
         );
  fd2qd1_hd r_add_B_reg_0_ ( .D(n1503), .CK(n1379), .RN(n172), .Q(r_add_B[0])
         );
  fd2qd1_hd r_mult_Z_ACK_reg ( .D(n1384), .CK(i_CLK), .RN(n665), .Q(
        r_mult_Z_ACK) );
  fd2qd1_hd r_add_A_reg_31_ ( .D(n1501), .CK(n1379), .RN(n603), .Q(r_add_A[31]) );
  fd2qd1_hd r_counter_reg_0_ ( .D(n1386), .CK(i_CLK), .RN(n603), .Q(
        r_counter[0]) );
  fd2qd1_hd r_add_A_reg_30_ ( .D(n1500), .CK(n1379), .RN(n634), .Q(r_add_A[30]) );
  fd2qd1_hd r_add_A_reg_29_ ( .D(n1499), .CK(n1379), .RN(n598), .Q(r_add_A[29]) );
  fd2qd1_hd r_add_A_reg_28_ ( .D(n1498), .CK(n1379), .RN(n668), .Q(r_add_A[28]) );
  fd2qd1_hd r_add_A_reg_27_ ( .D(n1497), .CK(n1379), .RN(n598), .Q(r_add_A[27]) );
  fd2qd1_hd r_add_A_reg_26_ ( .D(n1496), .CK(n1379), .RN(n632), .Q(r_add_A[26]) );
  fd2qd1_hd r_add_A_reg_25_ ( .D(n1495), .CK(n1379), .RN(n616), .Q(r_add_A[25]) );
  fd2qd1_hd r_add_A_reg_24_ ( .D(n1494), .CK(n1379), .RN(n665), .Q(r_add_A[24]) );
  fd2qd1_hd r_add_A_reg_23_ ( .D(n1493), .CK(n1379), .RN(n666), .Q(r_add_A[23]) );
  fd2qd1_hd r_add_A_reg_22_ ( .D(n1492), .CK(n1379), .RN(n668), .Q(r_add_A[22]) );
  fd2qd1_hd r_add_A_reg_21_ ( .D(n1491), .CK(n1379), .RN(n616), .Q(r_add_A[21]) );
  fd2qd1_hd r_add_A_reg_20_ ( .D(n1490), .CK(n1379), .RN(n603), .Q(r_add_A[20]) );
  fd2qd1_hd r_add_A_reg_19_ ( .D(n1489), .CK(n1379), .RN(n603), .Q(r_add_A[19]) );
  fd2qd1_hd r_add_A_reg_18_ ( .D(n1488), .CK(n1379), .RN(n732), .Q(r_add_A[18]) );
  fd2qd1_hd r_add_A_reg_17_ ( .D(n1487), .CK(n1379), .RN(n632), .Q(r_add_A[17]) );
  fd2qd1_hd r_add_A_reg_16_ ( .D(n1486), .CK(n1379), .RN(n665), .Q(r_add_A[16]) );
  fd2qd1_hd r_add_A_reg_15_ ( .D(n1485), .CK(n1379), .RN(n599), .Q(r_add_A[15]) );
  fd2qd1_hd r_add_A_reg_14_ ( .D(n1484), .CK(n1379), .RN(n172), .Q(r_add_A[14]) );
  fd2qd1_hd r_add_A_reg_13_ ( .D(n1483), .CK(n1379), .RN(n732), .Q(r_add_A[13]) );
  fd2qd1_hd r_add_A_reg_12_ ( .D(n1482), .CK(n1379), .RN(n733), .Q(r_add_A[12]) );
  fd2qd1_hd r_add_A_reg_11_ ( .D(n1481), .CK(n1379), .RN(n631), .Q(r_add_A[11]) );
  fd2qd1_hd r_add_A_reg_10_ ( .D(n1480), .CK(n1379), .RN(n633), .Q(r_add_A[10]) );
  fd2qd1_hd r_add_A_reg_9_ ( .D(n1479), .CK(n1379), .RN(n792), .Q(r_add_A[9])
         );
  fd2qd1_hd r_add_A_reg_8_ ( .D(n1478), .CK(n1379), .RN(n598), .Q(r_add_A[8])
         );
  fd2qd1_hd r_add_A_reg_7_ ( .D(n1477), .CK(n1379), .RN(n858), .Q(r_add_A[7])
         );
  fd2qd1_hd r_add_A_reg_6_ ( .D(n1476), .CK(n1379), .RN(n596), .Q(r_add_A[6])
         );
  fd2qd1_hd r_add_A_reg_5_ ( .D(n1475), .CK(n1379), .RN(n632), .Q(r_add_A[5])
         );
  fd2qd1_hd r_add_A_reg_4_ ( .D(n1474), .CK(n1379), .RN(n857), .Q(r_add_A[4])
         );
  fd2qd1_hd r_add_A_reg_3_ ( .D(n1473), .CK(n1379), .RN(n857), .Q(r_add_A[3])
         );
  fd2qd1_hd r_add_A_reg_2_ ( .D(n1472), .CK(n1379), .RN(n634), .Q(r_add_A[2])
         );
  fd2qd1_hd r_add_A_reg_1_ ( .D(n1471), .CK(n1379), .RN(w_rstn), .Q(r_add_A[1]) );
  fd2qd1_hd r_add_A_reg_0_ ( .D(n1470), .CK(n1379), .RN(n733), .Q(r_add_A[0])
         );
  fd2qd1_hd r_mult_2_A_reg_29_ ( .D(n1540), .CK(n1378), .RN(n792), .Q(
        r_mult_2_A[29]) );
  fd2qd1_hd r_mult_2_A_reg_28_ ( .D(n1540), .CK(n1378), .RN(n599), .Q(
        r_mult_2_A[28]) );
  fd2qd1_hd r_mult_2_A_reg_27_ ( .D(n1540), .CK(n1378), .RN(n733), .Q(
        r_mult_2_A[27]) );
  fd2qd1_hd r_mult_2_A_reg_26_ ( .D(n1541), .CK(n1378), .RN(n857), .Q(
        r_mult_2_A[26]) );
  fd2qd1_hd r_mult_2_A_reg_20_ ( .D(n1540), .CK(n1378), .RN(n636), .Q(
        r_mult_2_A[20]) );
  fd2qd1_hd r_mult_2_A_reg_17_ ( .D(n1541), .CK(n1378), .RN(n666), .Q(
        r_mult_2_A[17]) );
  fd2qd1_hd r_mult_2_A_reg_16_ ( .D(n1541), .CK(n1378), .RN(n172), .Q(
        r_mult_2_A[16]) );
  fd2qd1_hd r_mult_2_A_reg_11_ ( .D(n1541), .CK(n1378), .RN(n665), .Q(
        r_mult_2_A[11]) );
  fd2qd1_hd r_mult_2_A_reg_10_ ( .D(n1540), .CK(n1378), .RN(n631), .Q(
        r_mult_2_A[10]) );
  fd2qd1_hd r_mult_2_A_reg_7_ ( .D(n1541), .CK(n1378), .RN(n864), .Q(
        r_mult_2_A[7]) );
  fd2qd1_hd r_mult_2_A_reg_6_ ( .D(n1540), .CK(n1378), .RN(n858), .Q(
        r_mult_2_A[6]) );
  fd2qd1_hd r_mult_2_A_reg_5_ ( .D(n1540), .CK(n1378), .RN(n864), .Q(
        r_mult_2_A[5]) );
  fd2qd1_hd r_mult_2_A_reg_3_ ( .D(n1541), .CK(n1378), .RN(n598), .Q(
        r_mult_2_A[3]) );
  fd2qd1_hd r_mult_2_A_reg_0_ ( .D(n1541), .CK(n1378), .RN(n792), .Q(
        r_mult_2_A[0]) );
  fd2qd1_hd r_mult_1_A_reg_29_ ( .D(n1540), .CK(n1378), .RN(n596), .Q(
        r_mult_1_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_28_ ( .D(n1540), .CK(n1378), .RN(n858), .Q(
        r_mult_1_A[28]) );
  fd2qd1_hd r_mult_1_A_reg_27_ ( .D(n1541), .CK(n1378), .RN(n792), .Q(
        r_mult_1_A[27]) );
  fd2qd1_hd r_mult_1_A_reg_26_ ( .D(n1540), .CK(n1378), .RN(n792), .Q(
        r_mult_1_A[26]) );
  fd2qd1_hd r_mult_1_A_reg_23_ ( .D(n1541), .CK(n1378), .RN(n602), .Q(
        r_mult_1_A[23]) );
  fd2qd1_hd r_mult_1_A_reg_22_ ( .D(n1540), .CK(n1378), .RN(n602), .Q(
        r_mult_1_A[22]) );
  fd2qd1_hd r_mult_1_A_reg_20_ ( .D(n1541), .CK(n1378), .RN(n634), .Q(
        r_mult_1_A[20]) );
  fd2qd1_hd r_mult_1_A_reg_17_ ( .D(n1540), .CK(n1378), .RN(n603), .Q(
        r_mult_1_A[17]) );
  fd2qd1_hd r_mult_1_A_reg_11_ ( .D(n1541), .CK(n1378), .RN(n668), .Q(
        r_mult_1_A[11]) );
  fd2qd1_hd r_mult_1_A_reg_10_ ( .D(n1541), .CK(n1378), .RN(n636), .Q(
        r_mult_1_A[10]) );
  fd2qd1_hd r_mult_1_A_reg_7_ ( .D(n1541), .CK(n1378), .RN(n915), .Q(
        r_mult_1_A[7]) );
  fd2qd1_hd r_mult_1_A_reg_6_ ( .D(n1541), .CK(n1378), .RN(n172), .Q(
        r_mult_1_A[6]) );
  fd2qd1_hd r_mult_1_A_reg_5_ ( .D(n1541), .CK(n1378), .RN(n603), .Q(
        r_mult_1_A[5]) );
  fd2qd1_hd r_mult_1_A_reg_3_ ( .D(n1540), .CK(n1378), .RN(n864), .Q(
        r_mult_1_A[3]) );
  clknd2d1_hd U1 ( .A(n255), .B(n1462), .Y(n1460) );
  ivd2_hd U2 ( .A(n167), .Y(n292) );
  clknd2d1_hd U3 ( .A(n982), .B(n969), .Y(n1391) );
  clknd2d1_hd U4 ( .A(r_pstate[1]), .B(n968), .Y(n1392) );
  ivd3_hd U5 ( .A(n964), .Y(n185) );
  ad2bd2_hd U7 ( .B(n965), .AN(n185), .Y(n165) );
  ad2d1_hd U8 ( .A(n970), .B(alt20_n15), .Y(N817) );
  mx2d1_hd U10 ( .D0(r_counter[0]), .D1(N564), .S(N806), .Y(n1386) );
  mx2d1_hd U12 ( .D0(r_mult_Z_ACK), .D1(n964), .S(N812), .Y(n1384) );
  scg2d1_hd U13 ( .A(r_y_data[32]), .B(n978), .C(n1537), .D(w_add_Z[0]), .Y(
        n1574) );
  scg2d1_hd U14 ( .A(r_y_data[33]), .B(n978), .C(n1538), .D(w_add_Z[1]), .Y(
        n1575) );
  scg2d1_hd U15 ( .A(r_y_data[34]), .B(n978), .C(n1537), .D(w_add_Z[2]), .Y(
        n1576) );
  scg2d1_hd U16 ( .A(r_y_data[35]), .B(n978), .C(n1537), .D(w_add_Z[3]), .Y(
        n1577) );
  scg2d1_hd U17 ( .A(r_y_data[36]), .B(n978), .C(n1538), .D(w_add_Z[4]), .Y(
        n1578) );
  scg2d1_hd U18 ( .A(r_y_data[37]), .B(n978), .C(n1539), .D(w_add_Z[5]), .Y(
        n1579) );
  scg2d1_hd U19 ( .A(r_y_data[38]), .B(n978), .C(n1539), .D(w_add_Z[6]), .Y(
        n1580) );
  scg2d1_hd U20 ( .A(r_y_data[39]), .B(n978), .C(n1537), .D(w_add_Z[7]), .Y(
        n1581) );
  scg2d1_hd U21 ( .A(r_y_data[40]), .B(n978), .C(n1538), .D(w_add_Z[8]), .Y(
        n1582) );
  scg2d1_hd U22 ( .A(r_y_data[41]), .B(n978), .C(n1537), .D(w_add_Z[9]), .Y(
        n1583) );
  scg2d1_hd U23 ( .A(r_y_data[42]), .B(n978), .C(n1538), .D(w_add_Z[10]), .Y(
        n1584) );
  scg2d1_hd U24 ( .A(r_y_data[43]), .B(n978), .C(n1539), .D(w_add_Z[11]), .Y(
        n1585) );
  scg2d1_hd U25 ( .A(r_y_data[44]), .B(n978), .C(n1537), .D(w_add_Z[12]), .Y(
        n1586) );
  scg2d1_hd U26 ( .A(r_y_data[45]), .B(n978), .C(n1538), .D(w_add_Z[13]), .Y(
        n1587) );
  scg2d1_hd U27 ( .A(r_y_data[46]), .B(n978), .C(n1539), .D(w_add_Z[14]), .Y(
        n1588) );
  scg2d1_hd U29 ( .A(r_y_data[47]), .B(n979), .C(n1537), .D(w_add_Z[15]), .Y(
        n1589) );
  scg2d1_hd U32 ( .A(r_y_data[48]), .B(n980), .C(n1538), .D(w_add_Z[16]), .Y(
        n1590) );
  scg2d1_hd U33 ( .A(r_y_data[49]), .B(n980), .C(n1539), .D(w_add_Z[17]), .Y(
        n1591) );
  scg2d1_hd U36 ( .A(r_y_data[50]), .B(n254), .C(n1537), .D(w_add_Z[18]), .Y(
        n1592) );
  scg2d1_hd U37 ( .A(r_y_data[51]), .B(n979), .C(n1539), .D(w_add_Z[19]), .Y(
        n1593) );
  scg2d1_hd U38 ( .A(r_y_data[52]), .B(n254), .C(n1537), .D(w_add_Z[20]), .Y(
        n1594) );
  scg2d1_hd U39 ( .A(r_y_data[53]), .B(n978), .C(n1537), .D(w_add_Z[21]), .Y(
        n1595) );
  scg2d1_hd U40 ( .A(r_y_data[54]), .B(n978), .C(n1538), .D(w_add_Z[22]), .Y(
        n1596) );
  scg2d1_hd U41 ( .A(r_y_data[55]), .B(n254), .C(n1539), .D(w_add_Z[23]), .Y(
        n1597) );
  scg2d1_hd U42 ( .A(r_y_data[56]), .B(n254), .C(n1538), .D(w_add_Z[24]), .Y(
        n1598) );
  scg2d1_hd U43 ( .A(r_y_data[57]), .B(n254), .C(n1539), .D(w_add_Z[25]), .Y(
        n1599) );
  scg2d1_hd U44 ( .A(r_y_data[58]), .B(n254), .C(n1538), .D(w_add_Z[26]), .Y(
        n1600) );
  scg2d1_hd U45 ( .A(r_y_data[59]), .B(n254), .C(n1537), .D(w_add_Z[27]), .Y(
        n1601) );
  scg2d1_hd U46 ( .A(r_y_data[60]), .B(n254), .C(n1538), .D(w_add_Z[28]), .Y(
        n1602) );
  scg2d1_hd U47 ( .A(r_y_data[61]), .B(n254), .C(n1539), .D(w_add_Z[29]), .Y(
        n1603) );
  scg2d1_hd U49 ( .A(r_y_data[62]), .B(n254), .C(n1539), .D(w_add_Z[30]), .Y(
        n1604) );
  scg2d1_hd U50 ( .A(n964), .B(r_x_data[32]), .C(r_y_data[0]), .D(n979), .Y(
        n1542) );
  scg2d1_hd U51 ( .A(n964), .B(r_x_data[34]), .C(r_y_data[2]), .D(n979), .Y(
        n1544) );
  scg2d1_hd U52 ( .A(n964), .B(r_x_data[36]), .C(r_y_data[4]), .D(n979), .Y(
        n1546) );
  scg2d1_hd U53 ( .A(n964), .B(r_x_data[38]), .C(r_y_data[6]), .D(n979), .Y(
        n1548) );
  scg2d1_hd U54 ( .A(n964), .B(r_x_data[40]), .C(r_y_data[8]), .D(n979), .Y(
        n1550) );
  scg2d1_hd U55 ( .A(n964), .B(r_x_data[42]), .C(r_y_data[10]), .D(n979), .Y(
        n1552) );
  scg2d1_hd U56 ( .A(n964), .B(r_x_data[44]), .C(r_y_data[12]), .D(n979), .Y(
        n1554) );
  scg2d1_hd U57 ( .A(n964), .B(r_x_data[46]), .C(r_y_data[14]), .D(n979), .Y(
        n1556) );
  scg2d1_hd U58 ( .A(n964), .B(r_x_data[48]), .C(r_y_data[16]), .D(n979), .Y(
        n1558) );
  mx2d1_hd U59 ( .D0(r_pstate[0]), .D1(n1467), .S(n1468), .Y(n1383) );
  clknd2d1_hd U60 ( .A(n1389), .B(n1390), .Y(n1467) );
  mx2d1_hd U61 ( .D0(r_add_Z_ACK), .D1(n964), .S(N813), .Y(n1387) );
  mx2d1_hd U62 ( .D0(o_Y_DATA_VALID), .D1(N561), .S(N804), .Y(n1388) );
  scg2d1_hd U67 ( .A(n964), .B(r_x_data[33]), .C(r_y_data[1]), .D(n980), .Y(
        n1543) );
  scg2d1_hd U69 ( .A(n964), .B(r_x_data[37]), .C(r_y_data[5]), .D(n980), .Y(
        n1547) );
  scg2d1_hd U70 ( .A(n964), .B(r_x_data[43]), .C(r_y_data[11]), .D(n980), .Y(
        n1553) );
  scg2d1_hd U71 ( .A(n964), .B(r_x_data[49]), .C(r_y_data[17]), .D(n980), .Y(
        n1559) );
  scg2d1_hd U72 ( .A(n964), .B(r_x_data[55]), .C(r_y_data[23]), .D(n980), .Y(
        n1565) );
  scg2d1_hd U73 ( .A(n964), .B(r_x_data[58]), .C(r_y_data[26]), .D(n980), .Y(
        n1568) );
  scg2d1_hd U74 ( .A(n964), .B(r_x_data[59]), .C(r_y_data[27]), .D(n980), .Y(
        n1569) );
  scg2d1_hd U75 ( .A(n964), .B(r_x_data[61]), .C(r_y_data[29]), .D(n980), .Y(
        n1571) );
  scg2d1_hd U76 ( .A(n964), .B(r_x_data[63]), .C(r_y_data[31]), .D(n980), .Y(
        n1573) );
  mx2d1_hd U77 ( .D0(r_add_AB_STB), .D1(n967), .S(N802), .Y(n1382) );
  mx2d1_hd U78 ( .D0(r_mult_AB_STB), .D1(N766), .S(N802), .Y(n1381) );
  mx2d1_hd U79 ( .D0(r_counter[1]), .D1(n1465), .S(n1466), .Y(n1385) );
  nr2d1_hd U80 ( .A(n964), .B(n978), .Y(n287) );
  nid2_hd U81 ( .A(w_rst), .Y(n577) );
  ivd3_hd U82 ( .A(n170), .Y(n289) );
  clknd2d1_hd U83 ( .A(N435), .B(n964), .Y(n170) );
  scg2d1_hd U84 ( .A(n964), .B(r_x_data[62]), .C(r_y_data[30]), .D(n981), .Y(
        n1572) );
  scg2d1_hd U85 ( .A(n964), .B(r_x_data[60]), .C(r_y_data[28]), .D(n981), .Y(
        n1570) );
  scg2d1_hd U86 ( .A(n964), .B(r_x_data[57]), .C(r_y_data[25]), .D(n981), .Y(
        n1567) );
  scg2d1_hd U87 ( .A(n964), .B(r_x_data[56]), .C(r_y_data[24]), .D(n981), .Y(
        n1566) );
  scg2d1_hd U88 ( .A(n964), .B(r_x_data[54]), .C(r_y_data[22]), .D(n981), .Y(
        n1564) );
  scg2d1_hd U89 ( .A(n964), .B(r_x_data[53]), .C(r_y_data[21]), .D(n981), .Y(
        n1563) );
  scg2d1_hd U90 ( .A(n964), .B(r_x_data[52]), .C(r_y_data[20]), .D(n981), .Y(
        n1562) );
  scg2d1_hd U91 ( .A(n964), .B(r_x_data[51]), .C(r_y_data[19]), .D(n981), .Y(
        n1561) );
  scg2d1_hd U92 ( .A(n964), .B(r_x_data[50]), .C(r_y_data[18]), .D(n981), .Y(
        n1560) );
  scg2d1_hd U93 ( .A(n964), .B(r_x_data[47]), .C(r_y_data[15]), .D(n981), .Y(
        n1557) );
  scg2d1_hd U94 ( .A(n964), .B(r_x_data[45]), .C(r_y_data[13]), .D(n981), .Y(
        n1555) );
  scg2d1_hd U95 ( .A(n964), .B(r_x_data[41]), .C(r_y_data[9]), .D(n981), .Y(
        n1551) );
  scg2d1_hd U96 ( .A(n964), .B(r_x_data[39]), .C(r_y_data[7]), .D(n981), .Y(
        n1549) );
  scg2d1_hd U99 ( .A(n964), .B(r_x_data[35]), .C(r_y_data[3]), .D(n981), .Y(
        n1545) );
  ivd2_hd U101 ( .A(n170), .Y(n1502) );
  ivd1_hd U102 ( .A(n185), .Y(n1539) );
  ivd1_hd U103 ( .A(n185), .Y(n1538) );
  ivd1_hd U104 ( .A(n185), .Y(n1537) );
  nr2d4_hd U105 ( .A(N39), .B(r_counter[0]), .Y(n965) );
  ivd1_hd U106 ( .A(r_counter[1]), .Y(N39) );
  nr2d4_hd U107 ( .A(r_counter[1]), .B(N40), .Y(n962) );
  ivd1_hd U108 ( .A(n287), .Y(n1541) );
  ivd1_hd U109 ( .A(n287), .Y(n1540) );
  ivd1_hd U110 ( .A(N35), .Y(n982) );
  oa21d1_hd U111 ( .A(n966), .B(n170), .C(n164), .Y(n1374) );
  ivd1_hd U112 ( .A(r_pstate[1]), .Y(N27) );
  nr2d1_hd U113 ( .A(r_counter[1]), .B(n355), .Y(n1465) );
  scg9d1_hd U114 ( .A(r_counter[0]), .B(n355), .C(N806), .Y(n1466) );
  oa211d1_hd U115 ( .A(n968), .B(N28), .C(r_pstate[1]), .D(n1000), .Y(n1390)
         );
  oa211d1_hd U116 ( .A(n969), .B(N28), .C(N35), .D(N27), .Y(n1389) );
  scg10d1_hd U117 ( .A(r_pstate[1]), .B(n1391), .C(n1000), .D(n1392), .Y(n1468) );
  scg4d1_hd U118 ( .A(w_mult_1_Z[0]), .B(n1502), .C(o_Y_DATA[0]), .D(n165), 
        .E(n978), .F(r_x_data[0]), .G(n292), .H(w_mult_2_Z[0]), .Y(n1470) );
  scg4d1_hd U119 ( .A(w_mult_1_Z[1]), .B(n1502), .C(o_Y_DATA[1]), .D(n165), 
        .E(n978), .F(r_x_data[1]), .G(n292), .H(w_mult_2_Z[1]), .Y(n1471) );
  scg4d1_hd U120 ( .A(w_mult_1_Z[2]), .B(n1502), .C(o_Y_DATA[2]), .D(n165), 
        .E(n978), .F(r_x_data[2]), .G(n292), .H(w_mult_2_Z[2]), .Y(n1472) );
  scg4d1_hd U121 ( .A(w_mult_1_Z[3]), .B(n1502), .C(o_Y_DATA[3]), .D(n165), 
        .E(n978), .F(r_x_data[3]), .G(n292), .H(w_mult_2_Z[3]), .Y(n1473) );
  scg4d1_hd U122 ( .A(w_mult_1_Z[4]), .B(n1502), .C(o_Y_DATA[4]), .D(n165), 
        .E(n978), .F(r_x_data[4]), .G(n292), .H(w_mult_2_Z[4]), .Y(n1474) );
  scg4d1_hd U123 ( .A(w_mult_1_Z[5]), .B(n1502), .C(o_Y_DATA[5]), .D(n165), 
        .E(n978), .F(r_x_data[5]), .G(n292), .H(w_mult_2_Z[5]), .Y(n1475) );
  scg4d1_hd U124 ( .A(w_mult_1_Z[6]), .B(n1502), .C(o_Y_DATA[6]), .D(n165), 
        .E(n978), .F(r_x_data[6]), .G(n292), .H(w_mult_2_Z[6]), .Y(n1476) );
  scg4d1_hd U125 ( .A(w_mult_1_Z[7]), .B(n1502), .C(o_Y_DATA[7]), .D(n165), 
        .E(n978), .F(r_x_data[7]), .G(n292), .H(w_mult_2_Z[7]), .Y(n1477) );
  scg4d1_hd U126 ( .A(w_mult_1_Z[8]), .B(n1502), .C(o_Y_DATA[8]), .D(n165), 
        .E(n978), .F(r_x_data[8]), .G(n292), .H(w_mult_2_Z[8]), .Y(n1478) );
  scg4d1_hd U127 ( .A(w_mult_1_Z[9]), .B(n1502), .C(o_Y_DATA[9]), .D(n165), 
        .E(n978), .F(r_x_data[9]), .G(n292), .H(w_mult_2_Z[9]), .Y(n1479) );
  scg4d1_hd U128 ( .A(w_mult_1_Z[10]), .B(n1502), .C(o_Y_DATA[10]), .D(n165), 
        .E(n978), .F(r_x_data[10]), .G(n292), .H(w_mult_2_Z[10]), .Y(n1480) );
  scg4d1_hd U129 ( .A(w_mult_1_Z[11]), .B(n1502), .C(o_Y_DATA[11]), .D(n165), 
        .E(n978), .F(r_x_data[11]), .G(n292), .H(w_mult_2_Z[11]), .Y(n1481) );
  scg4d1_hd U130 ( .A(w_mult_1_Z[12]), .B(n1502), .C(o_Y_DATA[12]), .D(n165), 
        .E(n978), .F(r_x_data[12]), .G(n292), .H(w_mult_2_Z[12]), .Y(n1482) );
  scg4d1_hd U131 ( .A(w_mult_1_Z[13]), .B(n1502), .C(o_Y_DATA[13]), .D(n165), 
        .E(n978), .F(r_x_data[13]), .G(n292), .H(w_mult_2_Z[13]), .Y(n1483) );
  scg4d1_hd U132 ( .A(w_mult_1_Z[14]), .B(n1502), .C(o_Y_DATA[14]), .D(n165), 
        .E(n978), .F(r_x_data[14]), .G(n292), .H(w_mult_2_Z[14]), .Y(n1484) );
  scg4d1_hd U133 ( .A(w_mult_1_Z[15]), .B(n1502), .C(o_Y_DATA[15]), .D(n165), 
        .E(n978), .F(r_x_data[15]), .G(n292), .H(w_mult_2_Z[15]), .Y(n1485) );
  scg4d1_hd U134 ( .A(w_mult_1_Z[16]), .B(n1502), .C(o_Y_DATA[16]), .D(n165), 
        .E(n978), .F(r_x_data[16]), .G(n292), .H(w_mult_2_Z[16]), .Y(n1486) );
  scg4d1_hd U135 ( .A(w_mult_1_Z[17]), .B(n1502), .C(o_Y_DATA[17]), .D(n165), 
        .E(n978), .F(r_x_data[17]), .G(n292), .H(w_mult_2_Z[17]), .Y(n1487) );
  scg4d1_hd U136 ( .A(w_mult_1_Z[18]), .B(n1502), .C(o_Y_DATA[18]), .D(n165), 
        .E(n978), .F(r_x_data[18]), .G(n292), .H(w_mult_2_Z[18]), .Y(n1488) );
  scg4d1_hd U137 ( .A(w_mult_1_Z[19]), .B(n1502), .C(o_Y_DATA[19]), .D(n165), 
        .E(n978), .F(r_x_data[19]), .G(n292), .H(w_mult_2_Z[19]), .Y(n1489) );
  scg4d1_hd U138 ( .A(w_mult_1_Z[20]), .B(n1502), .C(o_Y_DATA[20]), .D(n165), 
        .E(n978), .F(r_x_data[20]), .G(n292), .H(w_mult_2_Z[20]), .Y(n1490) );
  scg4d1_hd U139 ( .A(w_mult_1_Z[21]), .B(n1502), .C(o_Y_DATA[21]), .D(n165), 
        .E(n978), .F(r_x_data[21]), .G(n292), .H(w_mult_2_Z[21]), .Y(n1491) );
  scg4d1_hd U140 ( .A(w_mult_1_Z[22]), .B(n1502), .C(o_Y_DATA[22]), .D(n165), 
        .E(n978), .F(r_x_data[22]), .G(n292), .H(w_mult_2_Z[22]), .Y(n1492) );
  scg4d1_hd U141 ( .A(w_mult_1_Z[23]), .B(n1502), .C(o_Y_DATA[23]), .D(n165), 
        .E(n978), .F(r_x_data[23]), .G(n292), .H(w_mult_2_Z[23]), .Y(n1493) );
  scg4d1_hd U142 ( .A(w_mult_1_Z[24]), .B(n1502), .C(o_Y_DATA[24]), .D(n165), 
        .E(n978), .F(r_x_data[24]), .G(n292), .H(w_mult_2_Z[24]), .Y(n1494) );
  scg4d1_hd U143 ( .A(w_mult_1_Z[25]), .B(n1502), .C(o_Y_DATA[25]), .D(n165), 
        .E(n978), .F(r_x_data[25]), .G(n292), .H(w_mult_2_Z[25]), .Y(n1495) );
  scg4d1_hd U144 ( .A(w_mult_1_Z[26]), .B(n1502), .C(o_Y_DATA[26]), .D(n165), 
        .E(n978), .F(r_x_data[26]), .G(n292), .H(w_mult_2_Z[26]), .Y(n1496) );
  scg4d1_hd U145 ( .A(w_mult_1_Z[27]), .B(n1502), .C(o_Y_DATA[27]), .D(n165), 
        .E(n978), .F(r_x_data[27]), .G(n292), .H(w_mult_2_Z[27]), .Y(n1497) );
  scg4d1_hd U146 ( .A(w_mult_1_Z[28]), .B(n1502), .C(o_Y_DATA[28]), .D(n165), 
        .E(n978), .F(r_x_data[28]), .G(n292), .H(w_mult_2_Z[28]), .Y(n1498) );
  scg4d1_hd U147 ( .A(w_mult_1_Z[29]), .B(n1502), .C(o_Y_DATA[29]), .D(n165), 
        .E(n978), .F(r_x_data[29]), .G(n292), .H(w_mult_2_Z[29]), .Y(n1499) );
  scg4d1_hd U148 ( .A(w_mult_1_Z[30]), .B(n1502), .C(o_Y_DATA[30]), .D(n165), 
        .E(n978), .F(r_x_data[30]), .G(n292), .H(w_mult_2_Z[30]), .Y(n1500) );
  scg4d1_hd U149 ( .A(w_mult_1_Z[31]), .B(n1502), .C(n165), .D(o_Y_DATA[31]), 
        .E(n292), .F(w_mult_2_Z[31]), .G(r_x_data[31]), .H(n978), .Y(n1501) );
  oa21d1_hd U150 ( .A(n185), .B(n1393), .C(n1394), .Y(n1503) );
  ao22d1_hd U151 ( .A(w_mult_2_Z[0]), .B(n289), .C(n979), .D(r_x_data[64]), 
        .Y(n1394) );
  oa21d1_hd U152 ( .A(n965), .B(n962), .C(w_add_Z[0]), .Y(n1393) );
  oa21d1_hd U153 ( .A(n185), .B(n1395), .C(n1396), .Y(n1504) );
  ao22d1_hd U154 ( .A(w_mult_2_Z[1]), .B(n289), .C(n978), .D(r_x_data[65]), 
        .Y(n1396) );
  oa21d1_hd U155 ( .A(n965), .B(n962), .C(w_add_Z[1]), .Y(n1395) );
  oa21d1_hd U156 ( .A(n185), .B(n1397), .C(n1398), .Y(n1505) );
  ao22d1_hd U157 ( .A(w_mult_2_Z[2]), .B(n289), .C(n979), .D(r_x_data[66]), 
        .Y(n1398) );
  oa21d1_hd U158 ( .A(n965), .B(n962), .C(w_add_Z[2]), .Y(n1397) );
  oa21d1_hd U159 ( .A(n185), .B(n1399), .C(n1400), .Y(n1506) );
  ao22d1_hd U160 ( .A(w_mult_2_Z[3]), .B(n289), .C(n980), .D(r_x_data[67]), 
        .Y(n1400) );
  oa21d1_hd U161 ( .A(n965), .B(n962), .C(w_add_Z[3]), .Y(n1399) );
  oa21d1_hd U162 ( .A(n185), .B(n1401), .C(n1402), .Y(n1507) );
  ao22d1_hd U163 ( .A(w_mult_2_Z[4]), .B(n289), .C(n979), .D(r_x_data[68]), 
        .Y(n1402) );
  oa21d1_hd U166 ( .A(n965), .B(n962), .C(w_add_Z[4]), .Y(n1401) );
  oa21d1_hd U167 ( .A(n185), .B(n1403), .C(n1404), .Y(n1508) );
  ao22d1_hd U168 ( .A(w_mult_2_Z[5]), .B(n289), .C(n980), .D(r_x_data[69]), 
        .Y(n1404) );
  oa21d1_hd U169 ( .A(n965), .B(n962), .C(w_add_Z[5]), .Y(n1403) );
  oa21d1_hd U170 ( .A(n185), .B(n1405), .C(n1406), .Y(n1509) );
  ao22d1_hd U171 ( .A(w_mult_2_Z[6]), .B(n289), .C(n979), .D(r_x_data[70]), 
        .Y(n1406) );
  oa21d1_hd U172 ( .A(n965), .B(n962), .C(w_add_Z[6]), .Y(n1405) );
  oa21d1_hd U173 ( .A(n185), .B(n1407), .C(n1408), .Y(n1510) );
  ao22d1_hd U174 ( .A(w_mult_2_Z[7]), .B(n289), .C(n980), .D(r_x_data[71]), 
        .Y(n1408) );
  oa21d1_hd U175 ( .A(n965), .B(n962), .C(w_add_Z[7]), .Y(n1407) );
  oa21d1_hd U176 ( .A(n185), .B(n1409), .C(n1410), .Y(n1511) );
  ao22d1_hd U177 ( .A(w_mult_2_Z[8]), .B(n289), .C(n980), .D(r_x_data[72]), 
        .Y(n1410) );
  oa21d1_hd U178 ( .A(n965), .B(n962), .C(w_add_Z[8]), .Y(n1409) );
  oa21d1_hd U179 ( .A(n185), .B(n1411), .C(n1412), .Y(n1512) );
  ao22d1_hd U180 ( .A(w_mult_2_Z[9]), .B(n289), .C(n980), .D(r_x_data[73]), 
        .Y(n1412) );
  oa21d1_hd U181 ( .A(n965), .B(n962), .C(w_add_Z[9]), .Y(n1411) );
  oa21d1_hd U182 ( .A(n185), .B(n1413), .C(n1414), .Y(n1513) );
  ao22d1_hd U183 ( .A(w_mult_2_Z[10]), .B(n289), .C(n979), .D(r_x_data[74]), 
        .Y(n1414) );
  oa21d1_hd U184 ( .A(n965), .B(n962), .C(w_add_Z[10]), .Y(n1413) );
  oa21d1_hd U185 ( .A(n185), .B(n1415), .C(n1416), .Y(n1514) );
  ao22d1_hd U186 ( .A(w_mult_2_Z[11]), .B(n289), .C(n980), .D(r_x_data[75]), 
        .Y(n1416) );
  oa21d1_hd U187 ( .A(n965), .B(n962), .C(w_add_Z[11]), .Y(n1415) );
  oa21d1_hd U189 ( .A(n185), .B(n1417), .C(n1418), .Y(n1515) );
  ao22d1_hd U190 ( .A(w_mult_2_Z[12]), .B(n289), .C(n979), .D(r_x_data[76]), 
        .Y(n1418) );
  oa21d1_hd U191 ( .A(n965), .B(n962), .C(w_add_Z[12]), .Y(n1417) );
  oa21d1_hd U192 ( .A(n185), .B(n1419), .C(n1420), .Y(n1516) );
  ao22d1_hd U196 ( .A(w_mult_2_Z[13]), .B(n289), .C(n980), .D(r_x_data[77]), 
        .Y(n1420) );
  oa21d1_hd U197 ( .A(n965), .B(n962), .C(w_add_Z[13]), .Y(n1419) );
  oa21d1_hd U198 ( .A(n185), .B(n1421), .C(n1422), .Y(n1517) );
  ao22d1_hd U199 ( .A(w_mult_2_Z[14]), .B(n289), .C(n979), .D(r_x_data[78]), 
        .Y(n1422) );
  oa21d1_hd U201 ( .A(n965), .B(n962), .C(w_add_Z[14]), .Y(n1421) );
  oa21d1_hd U202 ( .A(n185), .B(n1423), .C(n1424), .Y(n1518) );
  ao22d1_hd U203 ( .A(w_mult_2_Z[15]), .B(n289), .C(n980), .D(r_x_data[79]), 
        .Y(n1424) );
  oa21d1_hd U204 ( .A(n965), .B(n962), .C(w_add_Z[15]), .Y(n1423) );
  oa21d1_hd U239 ( .A(n185), .B(n1425), .C(n1426), .Y(n1519) );
  ao22d1_hd U241 ( .A(w_mult_2_Z[16]), .B(n289), .C(n979), .D(r_x_data[80]), 
        .Y(n1426) );
  oa21d1_hd U242 ( .A(n965), .B(n962), .C(w_add_Z[16]), .Y(n1425) );
  oa21d1_hd U244 ( .A(n185), .B(n1427), .C(n1428), .Y(n1520) );
  ao22d1_hd U245 ( .A(w_mult_2_Z[17]), .B(n289), .C(n980), .D(r_x_data[81]), 
        .Y(n1428) );
  oa21d1_hd U247 ( .A(n965), .B(n962), .C(w_add_Z[17]), .Y(n1427) );
  oa21d1_hd U248 ( .A(n185), .B(n1429), .C(n1430), .Y(n1521) );
  ao22d1_hd U250 ( .A(w_mult_2_Z[18]), .B(n289), .C(n980), .D(r_x_data[82]), 
        .Y(n1430) );
  oa21d1_hd U251 ( .A(n965), .B(n962), .C(w_add_Z[18]), .Y(n1429) );
  oa21d1_hd U253 ( .A(n185), .B(n1431), .C(n1432), .Y(n1522) );
  ao22d1_hd U254 ( .A(w_mult_2_Z[19]), .B(n289), .C(n980), .D(r_x_data[83]), 
        .Y(n1432) );
  oa21d1_hd U256 ( .A(n965), .B(n962), .C(w_add_Z[19]), .Y(n1431) );
  oa21d1_hd U257 ( .A(n185), .B(n1433), .C(n1434), .Y(n1523) );
  ao22d1_hd U259 ( .A(w_mult_2_Z[20]), .B(n289), .C(n980), .D(r_x_data[84]), 
        .Y(n1434) );
  oa21d1_hd U260 ( .A(n965), .B(n962), .C(w_add_Z[20]), .Y(n1433) );
  oa21d1_hd U262 ( .A(n185), .B(n1435), .C(n1436), .Y(n1524) );
  ao22d1_hd U263 ( .A(w_mult_2_Z[21]), .B(n289), .C(n980), .D(r_x_data[85]), 
        .Y(n1436) );
  oa21d1_hd U265 ( .A(n965), .B(n962), .C(w_add_Z[21]), .Y(n1435) );
  oa21d1_hd U266 ( .A(n185), .B(n1437), .C(n1438), .Y(n1525) );
  ao22d1_hd U268 ( .A(w_mult_2_Z[22]), .B(n289), .C(n979), .D(r_x_data[86]), 
        .Y(n1438) );
  oa21d1_hd U269 ( .A(n965), .B(n962), .C(w_add_Z[22]), .Y(n1437) );
  oa21d1_hd U271 ( .A(n185), .B(n1439), .C(n1440), .Y(n1526) );
  ao22d1_hd U272 ( .A(w_mult_2_Z[23]), .B(n289), .C(n980), .D(r_x_data[87]), 
        .Y(n1440) );
  oa21d1_hd U274 ( .A(n965), .B(n962), .C(w_add_Z[23]), .Y(n1439) );
  oa21d1_hd U275 ( .A(n185), .B(n1441), .C(n1442), .Y(n1527) );
  ao22d1_hd U277 ( .A(w_mult_2_Z[24]), .B(n289), .C(n980), .D(r_x_data[88]), 
        .Y(n1442) );
  oa21d1_hd U278 ( .A(n965), .B(n962), .C(w_add_Z[24]), .Y(n1441) );
  oa21d1_hd U280 ( .A(n185), .B(n1443), .C(n1444), .Y(n1528) );
  ao22d1_hd U281 ( .A(w_mult_2_Z[25]), .B(n289), .C(n979), .D(r_x_data[89]), 
        .Y(n1444) );
  oa21d1_hd U283 ( .A(n965), .B(n962), .C(w_add_Z[25]), .Y(n1443) );
  oa21d1_hd U284 ( .A(n185), .B(n1445), .C(n1446), .Y(n1529) );
  ao22d1_hd U286 ( .A(w_mult_2_Z[26]), .B(n289), .C(n979), .D(r_x_data[90]), 
        .Y(n1446) );
  oa21d1_hd U287 ( .A(n965), .B(n962), .C(w_add_Z[26]), .Y(n1445) );
  oa21d1_hd U289 ( .A(n185), .B(n1447), .C(n1448), .Y(n1530) );
  ao22d1_hd U290 ( .A(w_mult_2_Z[27]), .B(n289), .C(n979), .D(r_x_data[91]), 
        .Y(n1448) );
  oa21d1_hd U292 ( .A(n965), .B(n962), .C(w_add_Z[27]), .Y(n1447) );
  oa21d1_hd U293 ( .A(n185), .B(n1449), .C(n1450), .Y(n1531) );
  ao22d1_hd U295 ( .A(w_mult_2_Z[28]), .B(n289), .C(n980), .D(r_x_data[92]), 
        .Y(n1450) );
  oa21d1_hd U296 ( .A(n965), .B(n962), .C(w_add_Z[28]), .Y(n1449) );
  oa21d1_hd U298 ( .A(n185), .B(n1451), .C(n1452), .Y(n1532) );
  ao22d1_hd U299 ( .A(w_mult_2_Z[29]), .B(n289), .C(n979), .D(r_x_data[93]), 
        .Y(n1452) );
  oa21d1_hd U301 ( .A(n965), .B(n962), .C(w_add_Z[29]), .Y(n1451) );
  oa21d1_hd U302 ( .A(n185), .B(n1453), .C(n1454), .Y(n1533) );
  ao22d1_hd U304 ( .A(w_mult_2_Z[30]), .B(n289), .C(n979), .D(r_x_data[94]), 
        .Y(n1454) );
  oa21d1_hd U305 ( .A(n965), .B(n962), .C(w_add_Z[30]), .Y(n1453) );
  oa21d1_hd U307 ( .A(n185), .B(n1455), .C(n1456), .Y(n1534) );
  ao22d1_hd U308 ( .A(w_mult_2_Z[31]), .B(n289), .C(n980), .D(r_x_data[95]), 
        .Y(n1456) );
  oa21d1_hd U310 ( .A(n965), .B(n962), .C(w_add_Z[31]), .Y(n1455) );
  oa22d1_hd U311 ( .A(n185), .B(n1457), .C(n972), .D(n1458), .Y(n1536) );
  nr2d1_hd U313 ( .A(n1459), .B(n1460), .Y(n1458) );
  scg12d1_hd U314 ( .A(n962), .B(w_add_Z[31]), .C(n185), .Y(n1459) );
  oa211d1_hd U316 ( .A(w_add_Z[31]), .B(n1460), .C(n965), .D(n1461), .Y(n1457)
         );
  nd2bd1_hd U317 ( .AN(w_add_Z_STB), .B(n972), .Y(n1461) );
  ao22d1_hd U319 ( .A(w_mult_2_Z[31]), .B(n289), .C(n980), .D(r_x_data[95]), 
        .Y(n1462) );
  oa22ad1_hd U320 ( .A(n190), .B(n185), .C(r_y_data[63]), .D(n978), .Y(n1605)
         );
  oa21d1_hd U322 ( .A(n1463), .B(n164), .C(n1464), .Y(n1607) );
  scg13d1_hd U323 ( .A(n966), .B(n170), .C(n164), .Y(n1464) );
  scg20d1_hd U325 ( .A(N818), .B(n969), .C(n979), .Y(n1463) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_notch_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module iir_notch ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   w_rstn, w_rst, w_add_1_AB_ACK, w_add_2_AB_ACK, w_add_AB_ACK,
         w_add_1_Z_STB, w_add_2_Z_STB, w_add_Z_STB, r_add_1_AB_STB,
         r_add_1_Z_ACK, r_add_2_AB_STB, r_add_2_Z_ACK, w_mult_1_Z_STB,
         w_mult_2_Z_STB, w_mult_3_Z_STB, w_mult_Z_STB, w_mult_1_AB_ACK,
         w_mult_2_AB_ACK, w_mult_3_AB_ACK, w_mult_AB_ACK, r_mult_3_AB_STB,
         r_mult_3_Z_ACK, N25, N32, N33, N34, N37, N44, N45, N46, N47, N48, N49,
         N52, N55, N58, N66, N131, N196, N325, N714, N715, N716, N719, N722,
         N723, N725, N730, N731, N739, N743, N754, N1000, N1001, N1003, N1004,
         N1005, N1343, N1376, N1378, N1379, N1382, N1398, N1399, N1401, N1402,
         N1403, N1406, N1407, N1408, N1410, N1411, N1417, N1418, N1419,
         alt59_n44, alt59_n45, alt59_n46, alt59_n73, alt59_n74, alt59_n75,
         alt59_n76, alt59_n135, alt59_n136, add_x_1_n1, n2, n3, n6, n7, n8, n9,
         n298, n303, n304, n306, n309, n311, n312, n314, n316, n317, n318,
         n319, n321, n322, n323, n324, n326, n327, n328, n334, n485, n518,
         n584, n838, n841, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n1500, n1501, n1502, n1503, n1504, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1518, n1543, n1544,
         n1550, n1559, n1560, n302, n308, n888, n889, n893, n895, n899, n938,
         n962, n964, n1021, n1062, n1073, n1097, n1101, n1104, n1117, n1207,
         n1235, n1341, n1353, n1370, n1372, n1384, n1394, n1401, n1420, n1424,
         n1431, n1434, n1442, n1443, n1446, n1447, n1458, n1461, n1463, n1466,
         n1468, n1471, n1647, n1673, n2122, n2178, n2181, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813;
  wire   [31:0] r_add_1_A;
  wire   [31:0] r_add_1_B;
  wire   [31:0] w_add_1_Z;
  wire   [31:0] r_add_2_A;
  wire   [31:0] r_add_2_B;
  wire   [31:0] w_add_2_Z;
  wire   [31:0] r_mult_1_A;
  wire   [31:0] r_mult_1_B;
  wire   [31:0] w_mult_1_Z;
  wire   [29:3] r_mult_2_A;
  wire   [31:0] r_mult_2_B;
  wire   [31:0] w_mult_2_Z;
  wire   [29:3] r_mult_3_A;
  wire   [31:0] r_mult_3_B;
  wire   [31:0] w_mult_3_Z;
  wire   [159:0] r_x_data;
  wire   [127:0] r_y_data;
  wire   [1:0] r_pstate;
  wire   [2:0] r_counter;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  float_adder add_1 ( .i_A(r_add_1_A), .i_B(r_add_1_B), .i_AB_STB(
        r_add_1_AB_STB), .o_AB_ACK(w_add_1_AB_ACK), .o_Z(w_add_1_Z), .o_Z_STB(
        w_add_1_Z_STB), .i_Z_ACK(r_add_1_Z_ACK), .i_CLK(i_CLK), .i_RST(n848)
         );
  float_adder add_2 ( .i_A(r_add_2_A), .i_B(r_add_2_B), .i_AB_STB(
        r_add_2_AB_STB), .o_AB_ACK(w_add_2_AB_ACK), .o_Z(w_add_2_Z), .o_Z_STB(
        w_add_2_Z_STB), .i_Z_ACK(r_add_2_Z_ACK), .i_CLK(i_CLK), .i_RST(n848)
         );
  float_multiplier mult_1 ( .i_A(r_mult_1_A), .i_B(r_mult_1_B), .i_AB_STB(
        n2242), .o_AB_ACK(w_mult_1_AB_ACK), .o_Z(w_mult_1_Z), .o_Z_STB(
        w_mult_1_Z_STB), .i_Z_ACK(n2241), .i_CLK(i_CLK), .i_RST(n848) );
  float_multiplier mult_2 ( .i_A({n2244, 1'b0, r_mult_2_A[29:25], n2245, 1'b0, 
        r_mult_2_A[22:21], n2243, n2244, n2240, n2245, 1'b0, n2245, n2244, 
        n2243, n2240, 1'b0, r_mult_2_A[10:8], n2244, r_mult_2_A[6:5], n2243, 
        r_mult_2_A[3], 1'b0, n2243, n2245}), .i_B(r_mult_2_B), .i_AB_STB(n2242), .o_AB_ACK(w_mult_2_AB_ACK), .o_Z(w_mult_2_Z), .o_Z_STB(w_mult_2_Z_STB), 
        .i_Z_ACK(n2241), .i_CLK(i_CLK), .i_RST(n848) );
  float_multiplier mult_3 ( .i_A({n2247, 1'b0, r_mult_3_A[29:25], n2247, n2247, 
        r_mult_3_A[22], n2247, n2246, n2246, n2247, r_mult_3_A[17], n2246, 
        n2247, n2246, n2246, r_mult_3_A[12], n2247, n2247, n2246, n2247, 
        r_mult_3_A[7], n2246, r_mult_3_A[5:3], n2247, n2246, n2246}), .i_B(
        r_mult_3_B), .i_AB_STB(r_mult_3_AB_STB), .o_AB_ACK(w_mult_3_AB_ACK), 
        .o_Z(w_mult_3_Z), .o_Z_STB(w_mult_3_Z_STB), .i_Z_ACK(r_mult_3_Z_ACK), 
        .i_CLK(i_CLK), .i_RST(n848) );
  had1_hd add_x_1_U2 ( .A(r_counter[1]), .B(r_counter[0]), .CO(add_x_1_n1), 
        .S(N730) );
  nd2bd1_hd U293 ( .AN(N48), .B(n3), .Y(N66) );
  nr4d1_hd U295 ( .A(n1511), .B(n1503), .C(n1501), .D(n1500), .Y(n3) );
  nr2d1_hd U298 ( .A(r_counter[0]), .B(N44), .Y(n6) );
  nr2d1_hd U299 ( .A(r_counter[0]), .B(N739), .Y(n7) );
  oa211d1_hd U300 ( .A(w_add_Z_STB), .B(N46), .C(r_counter[1]), .D(N44), .Y(n8) );
  ao22d1_hd U301 ( .A(N25), .B(N44), .C(w_add_1_Z_STB), .D(n6), .Y(n9) );
  oa22d1_hd U302 ( .A(n7), .B(n8), .C(n9), .D(r_counter[1]), .Y(N754) );
  scg6d1_hd U311 ( .A(n298), .B(N66), .C(n2235), .Y(N1401) );
  nr2d1_hd U312 ( .A(n321), .B(n1508), .Y(n298) );
  scg12d1_hd U315 ( .A(n1504), .B(w_add_1_Z_STB), .C(n2234), .Y(n304) );
  scg4d1_hd U327 ( .A(n317), .B(n1513), .C(n318), .D(n309), .E(N743), .F(n311), 
        .G(n2235), .H(N1411), .Y(n316) );
  ivd1_hd U328 ( .A(w_add_Z_STB), .Y(n318) );
  nr2bd1_hd U339 ( .AN(N196), .B(n321), .Y(N1379) );
  nr2bd1_hd U340 ( .AN(N131), .B(n321), .Y(N1378) );
  nr2bd1_hd U341 ( .AN(N325), .B(n321), .Y(N1343) );
  ivd1_hd U652 ( .A(n328), .Y(N1376) );
  scg20d1_hd U841 ( .A(n1508), .B(N1410), .C(n321), .Y(n322) );
  nd2d1_hd U843 ( .A(n303), .B(N48), .Y(n326) );
  nr2d1_hd U844 ( .A(n1508), .B(n321), .Y(n303) );
  ivd1_hd U845 ( .A(n1507), .Y(n321) );
  nr2bd1_hd U850 ( .AN(N731), .B(n485), .Y(N1005) );
  nr2bd1_hd U851 ( .AN(N730), .B(n485), .Y(N1004) );
  nr2d1_hd U852 ( .A(n485), .B(r_counter[0]), .Y(N1003) );
  nr3d1_hd U853 ( .A(n309), .B(n311), .C(n317), .Y(n485) );
  ad2d1_hd U863 ( .A(alt59_n136), .B(n1509), .Y(N1000) );
  nd2bd1_hd U1224 ( .AN(n2234), .B(n1502), .Y(n334) );
  clknd2d1_hd U1225 ( .A(N25), .B(n312), .Y(n1515) );
  or2d1_hd U1226 ( .A(n1503), .B(alt59_n75), .Y(alt59_n74) );
  or2d1_hd U1227 ( .A(n1501), .B(alt59_n76), .Y(alt59_n75) );
  or2d1_hd U1228 ( .A(n1500), .B(N48), .Y(alt59_n76) );
  ad2d1_hd U1229 ( .A(w_add_1_AB_ACK), .B(w_add_2_AB_ACK), .Y(w_add_AB_ACK) );
  ad2d1_hd U1230 ( .A(N1418), .B(w_mult_3_AB_ACK), .Y(w_mult_AB_ACK) );
  ad2d1_hd U1231 ( .A(w_mult_1_AB_ACK), .B(w_mult_2_AB_ACK), .Y(N1418) );
  ad2d1_hd U1232 ( .A(N47), .B(N46), .Y(N48) );
  ad2d1_hd U1233 ( .A(N44), .B(N45), .Y(N47) );
  ad2d1_hd U1235 ( .A(N714), .B(N46), .Y(N715) );
  ad2d1_hd U1236 ( .A(N44), .B(N45), .Y(N714) );
  ivd1_hd U1237 ( .A(r_counter[1]), .Y(N45) );
  ad2d1_hd U1238 ( .A(N1419), .B(w_mult_2_Z_STB), .Y(N739) );
  ad2d1_hd U1239 ( .A(w_add_Z_STB), .B(w_mult_1_Z_STB), .Y(N1419) );
  or2d1_hd U1240 ( .A(n1502), .B(N715), .Y(alt59_n46) );
  ad2d1_hd U1241 ( .A(N1417), .B(w_mult_3_Z_STB), .Y(w_mult_Z_STB) );
  ad2d1_hd U1242 ( .A(w_mult_1_Z_STB), .B(w_mult_2_Z_STB), .Y(N1417) );
  clknd2d1_hd U1245 ( .A(w_add_Z_STB), .B(n309), .Y(n1560) );
  clknd2d1_hd U1280 ( .A(n3), .B(alt59_n73), .Y(N1410) );
  or2d1_hd U1281 ( .A(n1511), .B(alt59_n74), .Y(alt59_n73) );
  ad2d1_hd U1282 ( .A(r_pstate[1]), .B(r_pstate[0]), .Y(alt59_n136) );
  or3d1_hd U1283 ( .A(N48), .B(n1500), .C(n1501), .Y(N196) );
  ivd1_hd U1285 ( .A(alt59_n136), .Y(alt59_n135) );
  clknd2d1_hd U1286 ( .A(n306), .B(n319), .Y(N1382) );
  clknd2d1_hd U1287 ( .A(N754), .B(n2235), .Y(n306) );
  ad2d1_hd U1288 ( .A(N32), .B(N33), .Y(N34) );
  ivd1_hd U1289 ( .A(N739), .Y(N743) );
  or2d1_hd U1290 ( .A(n2544), .B(alt59_n45), .Y(alt59_n44) );
  or2d1_hd U1291 ( .A(n1506), .B(alt59_n46), .Y(alt59_n45) );
  ad2d1_hd U1292 ( .A(w_add_1_Z_STB), .B(w_add_2_Z_STB), .Y(w_add_Z_STB) );
  clknd2d1_hd U1293 ( .A(n1514), .B(n334), .Y(n317) );
  mx2d1_hd U1359 ( .D0(r_add_2_Z_ACK), .D1(n2235), .S(N1399), .Y(n518) );
  mx2d1_hd U1575 ( .D0(r_mult_3_Z_ACK), .D1(n2235), .S(n851), .Y(n838) );
  or4d1_hd U1930 ( .A(N48), .B(n1500), .C(n1501), .D(n1503), .Y(N131) );
  mx2d1_hd U1965 ( .D0(r_add_1_Z_ACK), .D1(n2235), .S(N1398), .Y(n584) );
  clknd2d1_hd U1966 ( .A(n321), .B(n306), .Y(N1398) );
  mx2d1_hd U1967 ( .D0(r_counter[0]), .D1(N1003), .S(N1382), .Y(n844) );
  ad2d1_hd U1969 ( .A(N34), .B(w_rstn), .Y(N1402) );
  ad2d1_hd U1970 ( .A(N1401), .B(n888), .Y(N1403) );
  or2d1_hd U1971 ( .A(N48), .B(n1500), .Y(N325) );
  scg9d1_hd U1972 ( .A(n1514), .B(n1513), .C(n321), .Y(n845) );
  scg9d1_hd U1973 ( .A(N743), .B(n1559), .C(n847), .Y(n846) );
  ad2d1_hd U1974 ( .A(n1515), .B(n845), .Y(n847) );
  ivd1_hd U1977 ( .A(n314), .Y(n1514) );
  nid2_hd U1990 ( .A(w_rstn), .Y(n1550) );
  ad2d1_hd U1991 ( .A(w_add_Z_STB), .B(w_mult_Z_STB), .Y(N25) );
  ivd1_hd U1992 ( .A(N25), .Y(n1513) );
  mx2d1_hd U1996 ( .D0(r_counter[2]), .D1(N1005), .S(N1382), .Y(n843) );
  xo2d1_hd U1997 ( .A(add_x_1_n1), .B(r_counter[2]), .Y(N731) );
  or2d1_hd U1998 ( .A(r_counter[2]), .B(N45), .Y(N722) );
  or2d1_hd U1999 ( .A(r_counter[2]), .B(N45), .Y(N719) );
  or2d1_hd U2000 ( .A(r_counter[2]), .B(N45), .Y(N55) );
  or2d1_hd U2001 ( .A(r_counter[2]), .B(N45), .Y(N52) );
  nr2d4_hd U2005 ( .A(n2233), .B(N723), .Y(n309) );
  ivd1_hd U2007 ( .A(n311), .Y(n1559) );
  ivd1_hd U2664 ( .A(r_pstate[0]), .Y(N33) );
  nr2d1_hd U2669 ( .A(N52), .B(r_counter[0]), .Y(n1501) );
  nid4_hd U2670 ( .A(n1516), .Y(n1518) );
  nr2d1_hd U2674 ( .A(N55), .B(N46), .Y(n1503) );
  nr2d1_hd U2688 ( .A(N725), .B(r_counter[0]), .Y(n1504) );
  nr2d1_hd U2698 ( .A(r_pstate[1]), .B(N33), .Y(n1507) );
  clknd2d1_hd U2699 ( .A(w_mult_AB_ACK), .B(w_add_AB_ACK), .Y(n1508) );
  clknd2d1_hd U2700 ( .A(o_Y_DATA_VALID), .B(i_Y_ACK), .Y(n1509) );
  ivd2_hd U2704 ( .A(n2224), .Y(n1543) );
  ivd2_hd U2705 ( .A(n2224), .Y(n1544) );
  nid2_hd U2707 ( .A(n323), .Y(n1516) );
  scg8d1_hd U2708 ( .A(n303), .B(n1500), .C(n304), .D(alt59_n136), .Y(n1510)
         );
  nr2d1_hd U2709 ( .A(N58), .B(r_counter[0]), .Y(n1511) );
  nr2d1_hd U2711 ( .A(n1504), .B(alt59_n44), .Y(n1512) );
  or2d1_hd U2712 ( .A(n1504), .B(n1512), .Y(N1411) );
  ivd1_hd U2713 ( .A(N34), .Y(n319) );
  or2d1_hd U2714 ( .A(N34), .B(alt59_n136), .Y(N1001) );
  mx2d1_hd U2716 ( .D0(r_counter[1]), .D1(N1004), .S(N1382), .Y(n841) );
  or2d1_hd U2717 ( .A(N44), .B(r_counter[1]), .Y(N725) );
  or2d1_hd U2718 ( .A(N44), .B(r_counter[1]), .Y(N58) );
  or2d1_hd U2719 ( .A(r_counter[2]), .B(r_counter[1]), .Y(N49) );
  or2d1_hd U2720 ( .A(r_counter[2]), .B(r_counter[1]), .Y(N716) );
  ivd1_hd U7 ( .A(n2178), .Y(n302) );
  ivd1_hd U10 ( .A(n1647), .Y(n308) );
  ivd1_hd U52 ( .A(n1647), .Y(n888) );
  ivd1_hd U53 ( .A(n2181), .Y(n889) );
  ivd1_hd U57 ( .A(n2178), .Y(n893) );
  ivd1_hd U59 ( .A(n2122), .Y(n895) );
  ivd1_hd U63 ( .A(n2181), .Y(n899) );
  ivd1_hd U102 ( .A(n1647), .Y(n938) );
  ivd1_hd U126 ( .A(n1673), .Y(n962) );
  ivd1_hd U128 ( .A(n1673), .Y(n964) );
  ivd1_hd U185 ( .A(n2122), .Y(n1021) );
  ivd1_hd U226 ( .A(n2181), .Y(n1062) );
  ivd1_hd U237 ( .A(n1673), .Y(n1073) );
  ivd1_hd U261 ( .A(n2178), .Y(n1097) );
  ivd1_hd U265 ( .A(n2181), .Y(n1101) );
  ivd1_hd U268 ( .A(n2178), .Y(n1104) );
  ivd1_hd U281 ( .A(n2122), .Y(n1117) );
  ivd1_hd U754 ( .A(n2122), .Y(n1207) );
  ivd1_hd U857 ( .A(n1673), .Y(n1235) );
  ivd1_hd U964 ( .A(n2122), .Y(n1341) );
  ivd1_hd U976 ( .A(n2181), .Y(n1353) );
  ivd1_hd U993 ( .A(n2178), .Y(n1370) );
  ivd1_hd U995 ( .A(n2122), .Y(n1372) );
  ivd1_hd U1007 ( .A(n2181), .Y(n1384) );
  ivd1_hd U1017 ( .A(n2178), .Y(n1394) );
  ivd1_hd U1024 ( .A(n2181), .Y(n1401) );
  ivd1_hd U1043 ( .A(n2178), .Y(n1420) );
  ivd1_hd U1047 ( .A(n2181), .Y(n1424) );
  ivd1_hd U1054 ( .A(n2122), .Y(n1431) );
  ivd1_hd U1057 ( .A(n2181), .Y(n1434) );
  ivd1_hd U1065 ( .A(n2181), .Y(n1442) );
  ivd1_hd U1066 ( .A(n2122), .Y(n1443) );
  ivd1_hd U1069 ( .A(n2122), .Y(n1446) );
  ivd1_hd U1070 ( .A(n2178), .Y(n1447) );
  ivd1_hd U1081 ( .A(n2122), .Y(n1458) );
  ivd1_hd U1084 ( .A(n2122), .Y(n1461) );
  ivd1_hd U1086 ( .A(n1673), .Y(n1463) );
  ivd1_hd U1089 ( .A(n1673), .Y(n1466) );
  ivd1_hd U1091 ( .A(n2178), .Y(n1468) );
  ivd1_hd U1094 ( .A(n2181), .Y(n1471) );
  ivd1_hd U1212 ( .A(w_rstn), .Y(n1647) );
  ivd1_hd U2034 ( .A(n1420), .Y(n1673) );
  ivd1_hd U2483 ( .A(w_rstn), .Y(n2122) );
  ivd1_hd U2539 ( .A(w_rstn), .Y(n2178) );
  ivd1_hd U2542 ( .A(w_rstn), .Y(n2181) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_12 clk_gate_r_counter_reg_2__0 ( .CLK(i_CLK), 
        .EN(alt59_n135), .ENCLK(n2255), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_14 clk_gate_r_mult_2_AB_STB_reg_0 ( .CLK(
        i_CLK), .EN(N1401), .ENCLK(n2254), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_15 clk_gate_o_Y_DATA_reg_31__0 ( .CLK(i_CLK), 
        .EN(N1406), .ENCLK(n2253), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_16 clk_gate_r_mult_3_B_reg_22__0 ( .CLK(i_CLK), .EN(n2511), .ENCLK(n2252), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_17 clk_gate_r_add_1_B_reg_31__0 ( .CLK(i_CLK), 
        .EN(n2578), .ENCLK(n2251), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_18 clk_gate_r_add_2_B_reg_31__0 ( .CLK(i_CLK), 
        .EN(n2644), .ENCLK(n2250), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_19 clk_gate_r_mult_2_B_reg_31__0 ( .CLK(i_CLK), .EN(n2746), .ENCLK(n2249), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_notch_20 clk_gate_r_y_data_reg_101__0 ( .CLK(i_CLK), 
        .EN(n1543), .ENCLK(n2248), .TE(1'b0) );
  fd1eqd1_hd r_mult_3_AB_STB_reg ( .D(N1343), .E(N1403), .CK(n2254), .Q(
        r_mult_3_AB_STB) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n2), .E(N1402), .CK(n2255), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_counter_reg_2_ ( .D(n843), .CK(n2255), .RN(n1104), .Q(
        r_counter[2]) );
  fd2qd1_hd r_pstate_reg_1_ ( .D(n2256), .CK(i_CLK), .RN(n1104), .Q(
        r_pstate[1]) );
  fd2qd1_hd r_y_data_reg_114_ ( .D(r_y_data[82]), .CK(n2248), .RN(n1353), .Q(
        r_y_data[114]) );
  fd2qd1_hd r_y_data_reg_85_ ( .D(r_y_data[53]), .CK(n2248), .RN(n1117), .Q(
        r_y_data[85]) );
  fd2qd1_hd r_y_data_reg_84_ ( .D(r_y_data[52]), .CK(n2248), .RN(n895), .Q(
        r_y_data[84]) );
  fd2qd1_hd r_y_data_reg_83_ ( .D(r_y_data[51]), .CK(n2248), .RN(n938), .Q(
        r_y_data[83]) );
  fd2qd1_hd r_y_data_reg_82_ ( .D(r_y_data[50]), .CK(n2248), .RN(n1463), .Q(
        r_y_data[82]) );
  fd2qd1_hd r_y_data_reg_52_ ( .D(r_y_data[20]), .CK(n2248), .RN(n962), .Q(
        r_y_data[52]) );
  fd2qd1_hd r_y_data_reg_51_ ( .D(r_y_data[19]), .CK(n2248), .RN(n1447), .Q(
        r_y_data[51]) );
  fd2qd1_hd r_y_data_reg_50_ ( .D(r_y_data[18]), .CK(n2248), .RN(n964), .Q(
        r_y_data[50]) );
  fd2qd1_hd r_y_data_reg_122_ ( .D(r_y_data[90]), .CK(n2248), .RN(n1384), .Q(
        r_y_data[122]) );
  fd2qd1_hd r_y_data_reg_95_ ( .D(r_y_data[63]), .CK(n2248), .RN(n308), .Q(
        r_y_data[95]) );
  fd2qd1_hd r_y_data_reg_94_ ( .D(r_y_data[62]), .CK(n2248), .RN(n1431), .Q(
        r_y_data[94]) );
  fd2qd1_hd r_y_data_reg_63_ ( .D(r_y_data[31]), .CK(n2248), .RN(n1370), .Q(
        r_y_data[63]) );
  fd2qd1_hd r_y_data_reg_62_ ( .D(r_y_data[30]), .CK(n2248), .RN(n302), .Q(
        r_y_data[62]) );
  fd2qd1_hd r_y_data_reg_59_ ( .D(r_y_data[27]), .CK(n2248), .RN(n1073), .Q(
        r_y_data[59]) );
  fd2qd1_hd r_y_data_reg_57_ ( .D(r_y_data[25]), .CK(n2248), .RN(n1550), .Q(
        r_y_data[57]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(o_Y_DATA[29]), .CK(n2248), .RN(n895), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_x_data_reg_154_ ( .D(r_x_data[122]), .CK(n2248), .RN(n1443), .Q(
        r_x_data[154]) );
  fd2qd1_hd r_x_data_reg_153_ ( .D(r_x_data[121]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[153]) );
  fd2qd1_hd r_x_data_reg_152_ ( .D(r_x_data[120]), .CK(n2248), .RN(n1443), .Q(
        r_x_data[152]) );
  fd2qd1_hd r_x_data_reg_151_ ( .D(r_x_data[119]), .CK(n2248), .RN(n1073), .Q(
        r_x_data[151]) );
  fd2qd1_hd r_x_data_reg_150_ ( .D(r_x_data[118]), .CK(n2248), .RN(n1550), .Q(
        r_x_data[150]) );
  fd2qd1_hd r_x_data_reg_149_ ( .D(r_x_data[117]), .CK(n2248), .RN(n899), .Q(
        r_x_data[149]) );
  fd2qd1_hd r_x_data_reg_148_ ( .D(r_x_data[116]), .CK(n2248), .RN(n1101), .Q(
        r_x_data[148]) );
  fd2qd1_hd r_x_data_reg_147_ ( .D(r_x_data[115]), .CK(n2248), .RN(n893), .Q(
        r_x_data[147]) );
  fd2qd1_hd r_x_data_reg_129_ ( .D(r_x_data[97]), .CK(n2248), .RN(n893), .Q(
        r_x_data[129]) );
  fd2qd1_hd r_x_data_reg_121_ ( .D(r_x_data[89]), .CK(n2248), .RN(n1117), .Q(
        r_x_data[121]) );
  fd2qd1_hd r_x_data_reg_120_ ( .D(r_x_data[88]), .CK(n2248), .RN(n1097), .Q(
        r_x_data[120]) );
  fd2qd1_hd r_x_data_reg_119_ ( .D(r_x_data[87]), .CK(n2248), .RN(n1461), .Q(
        r_x_data[119]) );
  fd2qd1_hd r_x_data_reg_118_ ( .D(r_x_data[86]), .CK(n2248), .RN(n938), .Q(
        r_x_data[118]) );
  fd2qd1_hd r_x_data_reg_117_ ( .D(r_x_data[85]), .CK(n2248), .RN(n1384), .Q(
        r_x_data[117]) );
  fd2qd1_hd r_x_data_reg_116_ ( .D(r_x_data[84]), .CK(n2248), .RN(n962), .Q(
        r_x_data[116]) );
  fd2qd1_hd r_x_data_reg_115_ ( .D(r_x_data[83]), .CK(n2248), .RN(n1372), .Q(
        r_x_data[115]) );
  fd2qd1_hd r_x_data_reg_97_ ( .D(r_x_data[65]), .CK(n2248), .RN(n1101), .Q(
        r_x_data[97]) );
  fd2qd1_hd r_x_data_reg_94_ ( .D(r_x_data[62]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[94]) );
  fd2qd1_hd r_x_data_reg_89_ ( .D(r_x_data[57]), .CK(n2248), .RN(n1235), .Q(
        r_x_data[89]) );
  fd2qd1_hd r_x_data_reg_88_ ( .D(r_x_data[56]), .CK(n2248), .RN(n964), .Q(
        r_x_data[88]) );
  fd2qd1_hd r_x_data_reg_87_ ( .D(r_x_data[55]), .CK(n2248), .RN(n1353), .Q(
        r_x_data[87]) );
  fd2qd1_hd r_x_data_reg_86_ ( .D(r_x_data[54]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[86]) );
  fd2qd1_hd r_x_data_reg_85_ ( .D(r_x_data[53]), .CK(n2248), .RN(n1207), .Q(
        r_x_data[85]) );
  fd2qd1_hd r_x_data_reg_84_ ( .D(r_x_data[52]), .CK(n2248), .RN(n308), .Q(
        r_x_data[84]) );
  fd2qd1_hd r_x_data_reg_83_ ( .D(r_x_data[51]), .CK(n2248), .RN(n1420), .Q(
        r_x_data[83]) );
  fd2qd1_hd r_x_data_reg_64_ ( .D(r_x_data[32]), .CK(n2248), .RN(n1073), .Q(
        r_x_data[64]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(r_x_data[25]), .CK(n2248), .RN(n1073), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(r_x_data[24]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(r_x_data[23]), .CK(n2248), .RN(n1442), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(r_x_data[22]), .CK(n2248), .RN(n938), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(r_x_data[21]), .CK(n2248), .RN(n1384), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(r_x_data[20]), .CK(n2248), .RN(n962), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(r_x_data[19]), .CK(n2248), .RN(n889), .Q(
        r_x_data[51]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(n2208), .CK(n2253), .RN(n302), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(n2209), .CK(n2253), .RN(n308), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(n2214), .CK(n2253), .RN(n1443), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(n2213), .CK(n2253), .RN(n1463), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd R_6 ( .D(N1379), .CK(n2254), .RN(n1434), .Q(n2242) );
  fd2qd1_hd r_y_data_reg_117_ ( .D(r_y_data[85]), .CK(n2248), .RN(n1461), .Q(
        r_y_data[117]) );
  fd2qd1_hd r_y_data_reg_99_ ( .D(r_y_data[67]), .CK(n2248), .RN(n1434), .Q(
        r_y_data[99]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(n2201), .CK(n2253), .RN(n1434), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd r_y_data_reg_126_ ( .D(r_y_data[94]), .CK(n2248), .RN(n1458), .Q(
        r_y_data[126]) );
  fd2qd1_hd r_y_data_reg_125_ ( .D(r_y_data[93]), .CK(n2248), .RN(n1466), .Q(
        r_y_data[125]) );
  fd2qd1_hd r_y_data_reg_116_ ( .D(r_y_data[84]), .CK(n2248), .RN(n1446), .Q(
        r_y_data[116]) );
  fd2qd1_hd r_y_data_reg_115_ ( .D(r_y_data[83]), .CK(n2248), .RN(n1463), .Q(
        r_y_data[115]) );
  fd2qd1_hd r_y_data_reg_98_ ( .D(r_y_data[66]), .CK(n2248), .RN(n1424), .Q(
        r_y_data[98]) );
  fd2qd1_hd r_y_data_reg_97_ ( .D(r_y_data[65]), .CK(n2248), .RN(n1461), .Q(
        r_y_data[97]) );
  fd2qd1_hd r_y_data_reg_96_ ( .D(r_y_data[64]), .CK(n2248), .RN(n1431), .Q(
        r_y_data[96]) );
  fd2qd1_hd r_y_data_reg_93_ ( .D(r_y_data[61]), .CK(n2248), .RN(n893), .Q(
        r_y_data[93]) );
  fd2qd1_hd r_y_data_reg_91_ ( .D(r_y_data[59]), .CK(n2248), .RN(n1235), .Q(
        r_y_data[91]) );
  fd2qd1_hd r_y_data_reg_76_ ( .D(r_y_data[44]), .CK(n2248), .RN(n1463), .Q(
        r_y_data[76]) );
  fd2qd1_hd r_y_data_reg_75_ ( .D(r_y_data[43]), .CK(n2248), .RN(n1442), .Q(
        r_y_data[75]) );
  fd2qd1_hd r_y_data_reg_67_ ( .D(r_y_data[35]), .CK(n2248), .RN(n1471), .Q(
        r_y_data[67]) );
  fd2qd1_hd r_y_data_reg_66_ ( .D(r_y_data[34]), .CK(n2248), .RN(n1341), .Q(
        r_y_data[66]) );
  fd2qd1_hd r_y_data_reg_61_ ( .D(r_y_data[29]), .CK(n2248), .RN(n964), .Q(
        r_y_data[61]) );
  fd2qd1_hd r_y_data_reg_45_ ( .D(r_y_data[13]), .CK(n2248), .RN(n899), .Q(
        r_y_data[45]) );
  fd2qd1_hd r_y_data_reg_44_ ( .D(r_y_data[12]), .CK(n2248), .RN(n1341), .Q(
        r_y_data[44]) );
  fd2qd1_hd r_y_data_reg_43_ ( .D(r_y_data[11]), .CK(n2248), .RN(n1550), .Q(
        r_y_data[43]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(o_Y_DATA[22]), .CK(n2248), .RN(n964), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(o_Y_DATA[20]), .CK(n2248), .RN(n1468), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(o_Y_DATA[18]), .CK(n2248), .RN(n1446), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(o_Y_DATA[13]), .CK(n2248), .RN(n1353), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(o_Y_DATA[12]), .CK(n2248), .RN(n1207), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(o_Y_DATA[11]), .CK(n2248), .RN(n1341), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_x_data_reg_69_ ( .D(r_x_data[37]), .CK(n2248), .RN(n1370), .Q(
        r_x_data[69]) );
  fd2qd1_hd r_x_data_reg_67_ ( .D(r_x_data[35]), .CK(n2248), .RN(n964), .Q(
        r_x_data[67]) );
  fd2qd1_hd r_x_data_reg_66_ ( .D(r_x_data[34]), .CK(n2248), .RN(n1420), .Q(
        r_x_data[66]) );
  fd2qd1_hd r_x_data_reg_65_ ( .D(r_x_data[33]), .CK(n2248), .RN(n1458), .Q(
        r_x_data[65]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(r_x_data[4]), .CK(n2248), .RN(n962), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(r_x_data[2]), .CK(n2248), .RN(n938), .Q(
        r_x_data[34]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(n2223), .CK(n2253), .RN(n1446), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(n2210), .CK(n2253), .RN(n1073), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(n2220), .CK(n2253), .RN(n1101), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(n2219), .CK(n2253), .RN(n1101), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(n2218), .CK(n2253), .RN(n1468), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd r_y_data_reg_124_ ( .D(r_y_data[92]), .CK(n2248), .RN(n1443), .Q(
        r_y_data[124]) );
  fd2qd1_hd r_y_data_reg_110_ ( .D(r_y_data[78]), .CK(n2248), .RN(n964), .Q(
        r_y_data[110]) );
  fd2qd1_hd r_y_data_reg_109_ ( .D(r_y_data[77]), .CK(n2248), .RN(n1466), .Q(
        r_y_data[109]) );
  fd2qd1_hd r_y_data_reg_108_ ( .D(r_y_data[76]), .CK(n2248), .RN(n895), .Q(
        r_y_data[108]) );
  fd2qd1_hd r_y_data_reg_107_ ( .D(r_y_data[75]), .CK(n2248), .RN(n1097), .Q(
        r_y_data[107]) );
  fd2qd1_hd r_y_data_reg_77_ ( .D(r_y_data[45]), .CK(n2248), .RN(n1104), .Q(
        r_y_data[77]) );
  fd2qd1_hd r_y_data_reg_65_ ( .D(r_y_data[33]), .CK(n2248), .RN(n888), .Q(
        r_y_data[65]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(o_Y_DATA[30]), .CK(n2248), .RN(n889), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_0_ ( .D(o_Y_DATA[0]), .CK(n2248), .RN(n1443), .Q(
        r_y_data[0]) );
  fd2qd1_hd r_x_data_reg_133_ ( .D(r_x_data[101]), .CK(n2248), .RN(n308), .Q(
        r_x_data[133]) );
  fd2qd1_hd r_x_data_reg_132_ ( .D(r_x_data[100]), .CK(n2248), .RN(n1431), .Q(
        r_x_data[132]) );
  fd2qd1_hd r_x_data_reg_130_ ( .D(r_x_data[98]), .CK(n2248), .RN(n1466), .Q(
        r_x_data[130]) );
  fd2qd1_hd r_x_data_reg_128_ ( .D(r_x_data[96]), .CK(n2248), .RN(n308), .Q(
        r_x_data[128]) );
  fd2qd1_hd r_x_data_reg_101_ ( .D(r_x_data[69]), .CK(n2248), .RN(n1097), .Q(
        r_x_data[101]) );
  fd2qd1_hd r_x_data_reg_68_ ( .D(r_x_data[36]), .CK(n2248), .RN(n1104), .Q(
        r_x_data[68]) );
  fd2qd1_hd r_y_data_reg_127_ ( .D(r_y_data[95]), .CK(n2248), .RN(n899), .Q(
        r_y_data[127]) );
  fd2qd1_hd r_y_data_reg_64_ ( .D(r_y_data[32]), .CK(n2248), .RN(n889), .Q(
        r_y_data[64]) );
  fd2qd1_hd r_y_data_reg_60_ ( .D(r_y_data[28]), .CK(n2248), .RN(n889), .Q(
        r_y_data[60]) );
  fd2qd1_hd r_y_data_reg_35_ ( .D(r_y_data[3]), .CK(n2248), .RN(n1431), .Q(
        r_y_data[35]) );
  fd2qd1_hd r_y_data_reg_34_ ( .D(r_y_data[2]), .CK(n2248), .RN(n893), .Q(
        r_y_data[34]) );
  fd2qd1_hd r_y_data_reg_33_ ( .D(r_y_data[1]), .CK(n2248), .RN(n1370), .Q(
        r_y_data[33]) );
  fd2qd1_hd r_y_data_reg_32_ ( .D(r_y_data[0]), .CK(n2248), .RN(n895), .Q(
        r_y_data[32]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(o_Y_DATA[31]), .CK(n2248), .RN(n1434), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(o_Y_DATA[3]), .CK(n2248), .RN(n1384), .Q(
        r_y_data[3]) );
  fd2qd1_hd r_y_data_reg_2_ ( .D(o_Y_DATA[2]), .CK(n2248), .RN(n899), .Q(
        r_y_data[2]) );
  fd2qd1_hd r_y_data_reg_1_ ( .D(o_Y_DATA[1]), .CK(n2248), .RN(n1471), .Q(
        r_y_data[1]) );
  fd2qd1_hd r_x_data_reg_122_ ( .D(r_x_data[90]), .CK(n2248), .RN(n1370), .Q(
        r_x_data[122]) );
  fd2qd1_hd R_4 ( .D(n2235), .CK(n2249), .RN(n889), .Q(n2244) );
  fd2qd1_hd R_2 ( .D(n2235), .CK(n2252), .RN(n893), .Q(n2246) );
  fd2qd1_hd r_y_data_reg_49_ ( .D(r_y_data[17]), .CK(n2248), .RN(n938), .Q(
        r_y_data[49]) );
  fd2qd1_hd r_y_data_reg_48_ ( .D(r_y_data[16]), .CK(n2248), .RN(n1207), .Q(
        r_y_data[48]) );
  fd2qd1_hd r_y_data_reg_47_ ( .D(r_y_data[15]), .CK(n2248), .RN(n888), .Q(
        r_y_data[47]) );
  fd2qd1_hd r_y_data_reg_46_ ( .D(r_y_data[14]), .CK(n2248), .RN(n1550), .Q(
        r_y_data[46]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(o_Y_DATA[19]), .CK(n2248), .RN(n1207), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(o_Y_DATA[17]), .CK(n2248), .RN(n895), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(o_Y_DATA[16]), .CK(n2248), .RN(n962), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(o_Y_DATA[15]), .CK(n2248), .RN(n1207), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(o_Y_DATA[14]), .CK(n2248), .RN(n964), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_x_data_reg_131_ ( .D(r_x_data[99]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[131]) );
  fd2qd1_hd r_x_data_reg_100_ ( .D(r_x_data[68]), .CK(n2248), .RN(n938), .Q(
        r_x_data[100]) );
  fd2qd1_hd r_x_data_reg_99_ ( .D(r_x_data[67]), .CK(n2248), .RN(n1341), .Q(
        r_x_data[99]) );
  fd2qd1_hd r_x_data_reg_98_ ( .D(r_x_data[66]), .CK(n2248), .RN(n1341), .Q(
        r_x_data[98]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(r_x_data[1]), .CK(n2248), .RN(n308), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_y_data_reg_120_ ( .D(r_y_data[88]), .CK(n2248), .RN(n1468), .Q(
        r_y_data[120]) );
  fd2qd1_hd r_y_data_reg_119_ ( .D(r_y_data[87]), .CK(n2248), .RN(n1372), .Q(
        r_y_data[119]) );
  fd2qd1_hd r_y_data_reg_106_ ( .D(r_y_data[74]), .CK(n2248), .RN(n1104), .Q(
        r_y_data[106]) );
  fd2qd1_hd r_y_data_reg_105_ ( .D(r_y_data[73]), .CK(n2248), .RN(n1235), .Q(
        r_y_data[105]) );
  fd2qd1_hd r_y_data_reg_104_ ( .D(r_y_data[72]), .CK(n2248), .RN(n308), .Q(
        r_y_data[104]) );
  fd2qd1_hd r_y_data_reg_103_ ( .D(r_y_data[71]), .CK(n2248), .RN(n1442), .Q(
        r_y_data[103]) );
  fd2qd1_hd r_y_data_reg_102_ ( .D(r_y_data[70]), .CK(n2248), .RN(n889), .Q(
        r_y_data[102]) );
  fd2qd1_hd r_y_data_reg_101_ ( .D(r_y_data[69]), .CK(n2248), .RN(n1370), .Q(
        r_y_data[101]) );
  fd2qd1_hd r_y_data_reg_100_ ( .D(r_y_data[68]), .CK(n2248), .RN(n1446), .Q(
        r_y_data[100]) );
  fd2qd1_hd r_y_data_reg_89_ ( .D(r_y_data[57]), .CK(n2248), .RN(n1443), .Q(
        r_y_data[89]) );
  fd2qd1_hd r_y_data_reg_88_ ( .D(r_y_data[56]), .CK(n2248), .RN(n1117), .Q(
        r_y_data[88]) );
  fd2qd1_hd r_y_data_reg_87_ ( .D(r_y_data[55]), .CK(n2248), .RN(n1447), .Q(
        r_y_data[87]) );
  fd2qd1_hd r_y_data_reg_74_ ( .D(r_y_data[42]), .CK(n2248), .RN(n1434), .Q(
        r_y_data[74]) );
  fd2qd1_hd r_y_data_reg_73_ ( .D(r_y_data[41]), .CK(n2248), .RN(n964), .Q(
        r_y_data[73]) );
  fd2qd1_hd r_y_data_reg_72_ ( .D(r_y_data[40]), .CK(n2248), .RN(n1353), .Q(
        r_y_data[72]) );
  fd2qd1_hd r_y_data_reg_71_ ( .D(r_y_data[39]), .CK(n2248), .RN(n1372), .Q(
        r_y_data[71]) );
  fd2qd1_hd r_y_data_reg_70_ ( .D(r_y_data[38]), .CK(n2248), .RN(n899), .Q(
        r_y_data[70]) );
  fd2qd1_hd r_y_data_reg_69_ ( .D(r_y_data[37]), .CK(n2248), .RN(n1466), .Q(
        r_y_data[69]) );
  fd2qd1_hd r_y_data_reg_68_ ( .D(r_y_data[36]), .CK(n2248), .RN(n1466), .Q(
        r_y_data[68]) );
  fd2qd1_hd r_y_data_reg_56_ ( .D(r_y_data[24]), .CK(n2248), .RN(n1468), .Q(
        r_y_data[56]) );
  fd2qd1_hd r_y_data_reg_55_ ( .D(r_y_data[23]), .CK(n2248), .RN(n962), .Q(
        r_y_data[55]) );
  fd2qd1_hd r_y_data_reg_42_ ( .D(r_y_data[10]), .CK(n2248), .RN(n1466), .Q(
        r_y_data[42]) );
  fd2qd1_hd r_y_data_reg_41_ ( .D(r_y_data[9]), .CK(n2248), .RN(n1394), .Q(
        r_y_data[41]) );
  fd2qd1_hd r_y_data_reg_40_ ( .D(r_y_data[8]), .CK(n2248), .RN(n1394), .Q(
        r_y_data[40]) );
  fd2qd1_hd r_y_data_reg_39_ ( .D(r_y_data[7]), .CK(n2248), .RN(n1424), .Q(
        r_y_data[39]) );
  fd2qd1_hd r_y_data_reg_38_ ( .D(r_y_data[6]), .CK(n2248), .RN(n1021), .Q(
        r_y_data[38]) );
  fd2qd1_hd r_y_data_reg_37_ ( .D(r_y_data[5]), .CK(n2248), .RN(n899), .Q(
        r_y_data[37]) );
  fd2qd1_hd r_y_data_reg_36_ ( .D(r_y_data[4]), .CK(n2248), .RN(n899), .Q(
        r_y_data[36]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(o_Y_DATA[24]), .CK(n2248), .RN(n1431), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(o_Y_DATA[10]), .CK(n2248), .RN(n895), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(o_Y_DATA[9]), .CK(n2248), .RN(n1468), .Q(
        r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(o_Y_DATA[8]), .CK(n2248), .RN(n1372), .Q(
        r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(o_Y_DATA[7]), .CK(n2248), .RN(n1384), .Q(
        r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(o_Y_DATA[6]), .CK(n2248), .RN(n1073), .Q(
        r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(o_Y_DATA[5]), .CK(n2248), .RN(n893), .Q(
        r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(o_Y_DATA[4]), .CK(n2248), .RN(n1372), .Q(
        r_y_data[4]) );
  fd2qd1_hd r_x_data_reg_156_ ( .D(r_x_data[124]), .CK(n2248), .RN(n1550), .Q(
        r_x_data[156]) );
  fd2qd1_hd r_x_data_reg_127_ ( .D(r_x_data[95]), .CK(n2248), .RN(n1021), .Q(
        r_x_data[127]) );
  fd2qd1_hd r_x_data_reg_125_ ( .D(r_x_data[93]), .CK(n2248), .RN(n1207), .Q(
        r_x_data[125]) );
  fd2qd1_hd r_x_data_reg_95_ ( .D(r_x_data[63]), .CK(n2248), .RN(n1235), .Q(
        r_x_data[95]) );
  fd2qd1_hd r_x_data_reg_91_ ( .D(r_x_data[59]), .CK(n2248), .RN(n1446), .Q(
        r_x_data[91]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(r_x_data[28]), .CK(n2248), .RN(n1420), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_32_ ( .D(r_x_data[0]), .CK(n2248), .RN(n1461), .Q(
        r_x_data[32]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(n2200), .CK(n2253), .RN(n1420), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(n2202), .CK(n2253), .RN(n1341), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(n2203), .CK(n2253), .RN(n1117), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(n2222), .CK(n2253), .RN(n1372), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(n2212), .CK(n2253), .RN(n1446), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(n2211), .CK(n2253), .RN(n1461), .Q(
        o_Y_DATA[8]) );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(n2226), .CK(n2253), .RN(n1073), .Q(
        o_Y_DATA[0]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(n2232), .CK(n2253), .RN(n1401), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(n2231), .CK(n2253), .RN(n302), .Q(o_Y_DATA[9]) );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(n2230), .CK(n2253), .RN(n1207), .Q(
        o_Y_DATA[7]) );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(n2206), .CK(n2253), .RN(n1550), .Q(
        o_Y_DATA[6]) );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(n2229), .CK(n2253), .RN(n1101), .Q(
        o_Y_DATA[5]) );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(n2205), .CK(n2253), .RN(n1341), .Q(
        o_Y_DATA[4]) );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(n2204), .CK(n2253), .RN(n1384), .Q(
        o_Y_DATA[3]) );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(n2228), .CK(n2253), .RN(n1434), .Q(
        o_Y_DATA[2]) );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(n2227), .CK(n2253), .RN(n1550), .Q(
        o_Y_DATA[1]) );
  fd2qd1_hd r_y_data_reg_121_ ( .D(r_y_data[89]), .CK(n2248), .RN(n302), .Q(
        r_y_data[121]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(o_Y_DATA[23]), .CK(n2248), .RN(n1468), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_x_data_reg_96_ ( .D(r_x_data[64]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[96]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(r_x_data[31]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[63]) );
  fd2qd1_hd r_add_1_AB_STB_reg ( .D(n1507), .CK(n2254), .RN(n1431), .Q(
        r_add_1_AB_STB) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(N1376), .CK(n2253), .RN(n1461), .Q(
        o_Y_DATA[31]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(r_x_data[3]), .CK(n2248), .RN(n1207), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_add_2_AB_STB_reg ( .D(N1378), .CK(n2254), .RN(n1447), .Q(
        r_add_2_AB_STB) );
  fd2qd1_hd r_y_data_reg_118_ ( .D(r_y_data[86]), .CK(n2248), .RN(n1461), .Q(
        r_y_data[118]) );
  fd2qd1_hd r_y_data_reg_86_ ( .D(r_y_data[54]), .CK(n2248), .RN(n302), .Q(
        r_y_data[86]) );
  fd2qd1_hd r_y_data_reg_54_ ( .D(r_y_data[22]), .CK(n2248), .RN(n1353), .Q(
        r_y_data[54]) );
  fd2qd1_hd r_y_data_reg_53_ ( .D(r_y_data[21]), .CK(n2248), .RN(n1021), .Q(
        r_y_data[53]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(o_Y_DATA[26]), .CK(n2248), .RN(n1117), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(o_Y_DATA[21]), .CK(n2248), .RN(n1384), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_x_data_reg_126_ ( .D(r_x_data[94]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[126]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(r_x_data[29]), .CK(n2248), .RN(n1442), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(r_x_data[26]), .CK(n2248), .RN(n1341), .Q(
        r_x_data[58]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(n2221), .CK(n2253), .RN(n302), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd r_y_data_reg_90_ ( .D(r_y_data[58]), .CK(n2248), .RN(n1446), .Q(
        r_y_data[90]) );
  fd2qd1_hd r_y_data_reg_58_ ( .D(r_y_data[26]), .CK(n2248), .RN(n1073), .Q(
        r_y_data[58]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(o_Y_DATA[28]), .CK(n2248), .RN(n1434), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(o_Y_DATA[27]), .CK(n2248), .RN(n1442), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(o_Y_DATA[25]), .CK(n2248), .RN(n938), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_x_data_reg_159_ ( .D(r_x_data[127]), .CK(n2248), .RN(n1431), .Q(
        r_x_data[159]) );
  fd2qd1_hd r_x_data_reg_158_ ( .D(r_x_data[126]), .CK(n2248), .RN(n1235), .Q(
        r_x_data[158]) );
  fd2qd1_hd r_x_data_reg_157_ ( .D(r_x_data[125]), .CK(n2248), .RN(n1101), .Q(
        r_x_data[157]) );
  fd2qd1_hd r_x_data_reg_155_ ( .D(r_x_data[123]), .CK(n2248), .RN(n1021), .Q(
        r_x_data[155]) );
  fd2qd1_hd r_x_data_reg_124_ ( .D(r_x_data[92]), .CK(n2248), .RN(n1394), .Q(
        r_x_data[124]) );
  fd2qd1_hd r_x_data_reg_123_ ( .D(r_x_data[91]), .CK(n2248), .RN(n938), .Q(
        r_x_data[123]) );
  fd2qd1_hd r_x_data_reg_93_ ( .D(r_x_data[61]), .CK(n2248), .RN(n1117), .Q(
        r_x_data[93]) );
  fd2qd1_hd r_x_data_reg_92_ ( .D(r_x_data[60]), .CK(n2248), .RN(n1207), .Q(
        r_x_data[92]) );
  fd2qd1_hd r_x_data_reg_90_ ( .D(r_x_data[58]), .CK(n2248), .RN(n1468), .Q(
        r_x_data[90]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(r_x_data[30]), .CK(n2248), .RN(n1104), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(r_x_data[27]), .CK(n2248), .RN(n1468), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_y_data_reg_123_ ( .D(r_y_data[91]), .CK(n2248), .RN(n1104), .Q(
        r_y_data[123]) );
  fd2qd1_hd r_y_data_reg_113_ ( .D(r_y_data[81]), .CK(n2248), .RN(n1372), .Q(
        r_y_data[113]) );
  fd2qd1_hd r_y_data_reg_112_ ( .D(r_y_data[80]), .CK(n2248), .RN(n1434), .Q(
        r_y_data[112]) );
  fd2qd1_hd r_y_data_reg_111_ ( .D(r_y_data[79]), .CK(n2248), .RN(n1370), .Q(
        r_y_data[111]) );
  fd2qd1_hd r_y_data_reg_92_ ( .D(r_y_data[60]), .CK(n2248), .RN(n1458), .Q(
        r_y_data[92]) );
  fd2qd1_hd r_y_data_reg_81_ ( .D(r_y_data[49]), .CK(n2248), .RN(n1372), .Q(
        r_y_data[81]) );
  fd2qd1_hd r_y_data_reg_80_ ( .D(r_y_data[48]), .CK(n2248), .RN(n302), .Q(
        r_y_data[80]) );
  fd2qd1_hd r_y_data_reg_79_ ( .D(r_y_data[47]), .CK(n2248), .RN(n1420), .Q(
        r_y_data[79]) );
  fd2qd1_hd r_y_data_reg_78_ ( .D(r_y_data[46]), .CK(n2248), .RN(n1370), .Q(
        r_y_data[78]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(n2217), .CK(n2253), .RN(n888), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(n2216), .CK(n2253), .RN(n889), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(n2207), .CK(n2253), .RN(n895), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(n2215), .CK(n2253), .RN(n893), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd r_mult_2_A_reg_5_ ( .D(n314), .CK(n2249), .RN(n962), .Q(
        r_mult_2_A[5]) );
  fd2qd1_hd r_add_1_Z_ACK_reg ( .D(n584), .CK(n2255), .RN(n1447), .Q(
        r_add_1_Z_ACK) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(i_X_DATA[31]), .CK(n2248), .RN(n1073), .Q(
        r_x_data[31]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(i_X_DATA[30]), .CK(n2248), .RN(n1235), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(i_X_DATA[29]), .CK(n2248), .RN(n895), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(i_X_DATA[28]), .CK(n2248), .RN(n1104), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(i_X_DATA[27]), .CK(n2248), .RN(n1207), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(i_X_DATA[26]), .CK(n2248), .RN(n1550), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(i_X_DATA[25]), .CK(n2248), .RN(n1073), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(i_X_DATA[24]), .CK(n2248), .RN(n964), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(i_X_DATA[23]), .CK(n2248), .RN(n1446), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(i_X_DATA[22]), .CK(n2248), .RN(n1062), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(i_X_DATA[21]), .CK(n2248), .RN(n1442), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(i_X_DATA[20]), .CK(n2248), .RN(n1424), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(i_X_DATA[19]), .CK(n2248), .RN(n1341), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(i_X_DATA[18]), .CK(n2248), .RN(n302), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(i_X_DATA[4]), .CK(n2248), .RN(n1370), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(i_X_DATA[3]), .CK(n2248), .RN(n1235), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(i_X_DATA[2]), .CK(n2248), .RN(n1431), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(i_X_DATA[1]), .CK(n2248), .RN(n1446), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(i_X_DATA[0]), .CK(n2248), .RN(n1117), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_mult_1_A_reg_18_ ( .D(n2663), .CK(n2249), .RN(n1117), .Q(
        r_mult_1_A[18]) );
  fd2qd1_hd r_mult_1_A_reg_17_ ( .D(n2662), .CK(n2249), .RN(n1394), .Q(
        r_mult_1_A[17]) );
  fd2qd1_hd r_mult_1_A_reg_15_ ( .D(n2660), .CK(n2249), .RN(n1442), .Q(
        r_mult_1_A[15]) );
  fd2qd1_hd r_mult_1_A_reg_11_ ( .D(n2656), .CK(n2249), .RN(n1117), .Q(
        r_mult_1_A[11]) );
  fd2qd1_hd r_mult_1_A_reg_10_ ( .D(n2655), .CK(n2249), .RN(n1384), .Q(
        r_mult_1_A[10]) );
  fd2qd1_hd r_mult_1_A_reg_4_ ( .D(n2649), .CK(n2249), .RN(n1394), .Q(
        r_mult_1_A[4]) );
  fd2qd1_hd r_mult_1_A_reg_2_ ( .D(n2647), .CK(n2249), .RN(n1117), .Q(
        r_mult_1_A[2]) );
  fd2qd1_hd r_mult_1_B_reg_19_ ( .D(n2698), .CK(n2249), .RN(n1235), .Q(
        r_mult_1_B[19]) );
  fd2qd1_hd r_mult_1_B_reg_18_ ( .D(n2697), .CK(n2249), .RN(n899), .Q(
        r_mult_1_B[18]) );
  fd2qd1_hd r_mult_1_B_reg_17_ ( .D(n2696), .CK(n2249), .RN(n1062), .Q(
        r_mult_1_B[17]) );
  fd2qd1_hd r_mult_1_B_reg_16_ ( .D(n2695), .CK(n2249), .RN(n962), .Q(
        r_mult_1_B[16]) );
  fd2qd1_hd r_mult_1_B_reg_15_ ( .D(n2694), .CK(n2249), .RN(n1443), .Q(
        r_mult_1_B[15]) );
  fd2qd1_hd r_mult_1_B_reg_14_ ( .D(n2693), .CK(n2249), .RN(n1372), .Q(
        r_mult_1_B[14]) );
  fd2qd1_hd r_mult_1_B_reg_13_ ( .D(n2692), .CK(n2249), .RN(n308), .Q(
        r_mult_1_B[13]) );
  fd2qd1_hd r_mult_1_B_reg_12_ ( .D(n2691), .CK(n2249), .RN(n1434), .Q(
        r_mult_1_B[12]) );
  fd2qd1_hd r_mult_1_B_reg_11_ ( .D(n2690), .CK(n2249), .RN(n1401), .Q(
        r_mult_1_B[11]) );
  fd2qd1_hd r_mult_1_B_reg_10_ ( .D(n2689), .CK(n2249), .RN(n1458), .Q(
        r_mult_1_B[10]) );
  fd2qd1_hd r_mult_1_B_reg_8_ ( .D(n2687), .CK(n2249), .RN(n1463), .Q(
        r_mult_1_B[8]) );
  fd2qd1_hd r_mult_1_B_reg_29_ ( .D(n2708), .CK(n2249), .RN(n1104), .Q(
        r_mult_1_B[29]) );
  fd2qd1_hd r_mult_1_B_reg_9_ ( .D(n2688), .CK(n2249), .RN(n1341), .Q(
        r_mult_1_B[9]) );
  fd2qd1_hd r_mult_1_B_reg_7_ ( .D(n2686), .CK(n2249), .RN(n1235), .Q(
        r_mult_1_B[7]) );
  fd2qd1_hd r_mult_1_B_reg_6_ ( .D(n2685), .CK(n2249), .RN(n1420), .Q(
        r_mult_1_B[6]) );
  fd2qd1_hd r_mult_1_B_reg_5_ ( .D(n2684), .CK(n2249), .RN(n964), .Q(
        r_mult_1_B[5]) );
  fd2qd1_hd r_mult_1_B_reg_4_ ( .D(n2683), .CK(n2249), .RN(n893), .Q(
        r_mult_1_B[4]) );
  fd2qd1_hd r_mult_1_B_reg_3_ ( .D(n2682), .CK(n2249), .RN(n1471), .Q(
        r_mult_1_B[3]) );
  fd2qd1_hd r_mult_1_B_reg_2_ ( .D(n2681), .CK(n2249), .RN(n888), .Q(
        r_mult_1_B[2]) );
  fd2qd1_hd r_mult_1_B_reg_1_ ( .D(n2680), .CK(n2249), .RN(n889), .Q(
        r_mult_1_B[1]) );
  fd2qd1_hd r_mult_1_B_reg_0_ ( .D(n2679), .CK(n2249), .RN(n1420), .Q(
        r_mult_1_B[0]) );
  fd2qd1_hd r_mult_2_B_reg_11_ ( .D(n2724), .CK(n2249), .RN(n938), .Q(
        r_mult_2_B[11]) );
  fd2qd1_hd r_mult_3_B_reg_22_ ( .D(n2509), .CK(n2252), .RN(n1401), .Q(
        r_mult_3_B[22]) );
  fd2qd1_hd r_mult_3_B_reg_15_ ( .D(n2508), .CK(n2252), .RN(n1097), .Q(
        r_mult_3_B[15]) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n2258), .CK(i_CLK), .RN(n1447), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_mult_2_A_reg_21_ ( .D(n2225), .CK(n2249), .RN(n938), .Q(
        r_mult_2_A[21]) );
  fd2qd1_hd r_mult_2_A_reg_9_ ( .D(n2225), .CK(n2249), .RN(n1434), .Q(
        r_mult_2_A[9]) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(n2257), .CK(i_CLK), .RN(n302), .Q(r_pstate[0]) );
  fd2qd1_hd r_x_data_reg_146_ ( .D(n2813), .CK(n2248), .RN(n1447), .Q(
        r_x_data[146]) );
  fd2qd1_hd r_x_data_reg_145_ ( .D(n2812), .CK(n2248), .RN(n1372), .Q(
        r_x_data[145]) );
  fd2qd1_hd r_x_data_reg_144_ ( .D(n2811), .CK(n2248), .RN(n1447), .Q(
        r_x_data[144]) );
  fd2qd1_hd r_x_data_reg_143_ ( .D(n2810), .CK(n2248), .RN(n893), .Q(
        r_x_data[143]) );
  fd2qd1_hd r_x_data_reg_142_ ( .D(n2809), .CK(n2248), .RN(n1401), .Q(
        r_x_data[142]) );
  fd2qd1_hd r_x_data_reg_141_ ( .D(n2808), .CK(n2248), .RN(n1424), .Q(
        r_x_data[141]) );
  fd2qd1_hd r_x_data_reg_140_ ( .D(n2807), .CK(n2248), .RN(n1021), .Q(
        r_x_data[140]) );
  fd2qd1_hd r_x_data_reg_139_ ( .D(n2806), .CK(n2248), .RN(n1550), .Q(
        r_x_data[139]) );
  fd2qd1_hd r_x_data_reg_138_ ( .D(n2805), .CK(n2248), .RN(n1550), .Q(
        r_x_data[138]) );
  fd2qd1_hd r_x_data_reg_137_ ( .D(n2804), .CK(n2248), .RN(n1550), .Q(
        r_x_data[137]) );
  fd2qd1_hd r_x_data_reg_136_ ( .D(n2803), .CK(n2248), .RN(n1550), .Q(
        r_x_data[136]) );
  fd2qd1_hd r_x_data_reg_135_ ( .D(n2802), .CK(n2248), .RN(n1550), .Q(
        r_x_data[135]) );
  fd2qd1_hd r_x_data_reg_134_ ( .D(n2801), .CK(n2248), .RN(n1104), .Q(
        r_x_data[134]) );
  fd2qd1_hd r_x_data_reg_114_ ( .D(n2800), .CK(n2248), .RN(n1431), .Q(
        r_x_data[114]) );
  fd2qd1_hd r_x_data_reg_113_ ( .D(n2799), .CK(n2248), .RN(n1097), .Q(
        r_x_data[113]) );
  fd2qd1_hd r_x_data_reg_112_ ( .D(n2798), .CK(n2248), .RN(n1446), .Q(
        r_x_data[112]) );
  fd2qd1_hd r_x_data_reg_111_ ( .D(n2797), .CK(n2248), .RN(n1101), .Q(
        r_x_data[111]) );
  fd2qd1_hd r_x_data_reg_110_ ( .D(n2796), .CK(n2248), .RN(n1458), .Q(
        r_x_data[110]) );
  fd2qd1_hd r_x_data_reg_109_ ( .D(n2795), .CK(n2248), .RN(n1401), .Q(
        r_x_data[109]) );
  fd2qd1_hd r_x_data_reg_108_ ( .D(n2794), .CK(n2248), .RN(n1461), .Q(
        r_x_data[108]) );
  fd2qd1_hd r_x_data_reg_107_ ( .D(n2793), .CK(n2248), .RN(n1550), .Q(
        r_x_data[107]) );
  fd2qd1_hd r_x_data_reg_106_ ( .D(n2792), .CK(n2248), .RN(n1550), .Q(
        r_x_data[106]) );
  fd2qd1_hd r_x_data_reg_105_ ( .D(n2791), .CK(n2248), .RN(n1550), .Q(
        r_x_data[105]) );
  fd2qd1_hd r_x_data_reg_104_ ( .D(n2790), .CK(n2248), .RN(n1550), .Q(
        r_x_data[104]) );
  fd2qd1_hd r_x_data_reg_103_ ( .D(n2789), .CK(n2248), .RN(n1550), .Q(
        r_x_data[103]) );
  fd2qd1_hd r_x_data_reg_102_ ( .D(n2788), .CK(n2248), .RN(n1104), .Q(
        r_x_data[102]) );
  fd2qd1_hd r_x_data_reg_82_ ( .D(n2787), .CK(n2248), .RN(n889), .Q(
        r_x_data[82]) );
  fd2qd1_hd r_x_data_reg_81_ ( .D(n2786), .CK(n2248), .RN(n1021), .Q(
        r_x_data[81]) );
  fd2qd1_hd r_x_data_reg_80_ ( .D(n2785), .CK(n2248), .RN(n1431), .Q(
        r_x_data[80]) );
  fd2qd1_hd r_x_data_reg_79_ ( .D(n2784), .CK(n2248), .RN(n1471), .Q(
        r_x_data[79]) );
  fd2qd1_hd r_x_data_reg_78_ ( .D(n2783), .CK(n2248), .RN(n1463), .Q(
        r_x_data[78]) );
  fd2qd1_hd r_x_data_reg_77_ ( .D(n2782), .CK(n2248), .RN(n1424), .Q(
        r_x_data[77]) );
  fd2qd1_hd r_x_data_reg_76_ ( .D(n2781), .CK(n2248), .RN(n1466), .Q(
        r_x_data[76]) );
  fd2qd1_hd r_x_data_reg_75_ ( .D(n2780), .CK(n2248), .RN(n1446), .Q(
        r_x_data[75]) );
  fd2qd1_hd r_x_data_reg_74_ ( .D(n2779), .CK(n2248), .RN(n1550), .Q(
        r_x_data[74]) );
  fd2qd1_hd r_x_data_reg_73_ ( .D(n2778), .CK(n2248), .RN(n1550), .Q(
        r_x_data[73]) );
  fd2qd1_hd r_x_data_reg_72_ ( .D(n2777), .CK(n2248), .RN(n1550), .Q(
        r_x_data[72]) );
  fd2qd1_hd r_x_data_reg_71_ ( .D(n2776), .CK(n2248), .RN(n1550), .Q(
        r_x_data[71]) );
  fd2qd1_hd r_x_data_reg_70_ ( .D(n2775), .CK(n2248), .RN(n1550), .Q(
        r_x_data[70]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(n2774), .CK(n2248), .RN(n1341), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(n2773), .CK(n2248), .RN(n1062), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(n2772), .CK(n2248), .RN(n308), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(n2771), .CK(n2248), .RN(n1468), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(n2770), .CK(n2248), .RN(n1458), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(n2769), .CK(n2248), .RN(n1471), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(n2768), .CK(n2248), .RN(n1461), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(n2767), .CK(n2248), .RN(n1207), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(n2766), .CK(n2248), .RN(n1550), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(n2765), .CK(n2248), .RN(n1550), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(n2764), .CK(n2248), .RN(n1550), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(n2763), .CK(n2248), .RN(n1550), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(n2762), .CK(n2248), .RN(n1550), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(n2761), .CK(n2248), .RN(n1463), .Q(
        r_x_data[37]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(n2760), .CK(n2248), .RN(n889), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(n2759), .CK(n2248), .RN(n1372), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(n2758), .CK(n2248), .RN(n1463), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(n2757), .CK(n2248), .RN(n1207), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(n2756), .CK(n2248), .RN(n1466), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(n2755), .CK(n2248), .RN(n1341), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(n2754), .CK(n2248), .RN(n1468), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(n2753), .CK(n2248), .RN(n1550), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(n2752), .CK(n2248), .RN(n1550), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(n2751), .CK(n2248), .RN(n1550), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(n2750), .CK(n2248), .RN(n1550), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(n2749), .CK(n2248), .RN(n1550), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(n2748), .CK(n2248), .RN(n1207), .Q(
        r_x_data[5]) );
  fd2qd1_hd R_3 ( .D(n312), .CK(n2249), .RN(n1021), .Q(n2245) );
  fd2qd1_hd r_mult_3_A_reg_29_ ( .D(n2477), .CK(n2252), .RN(n1394), .Q(
        r_mult_3_A[29]) );
  fd2qd1_hd r_mult_3_A_reg_28_ ( .D(n2476), .CK(n2252), .RN(n1104), .Q(
        r_mult_3_A[28]) );
  fd2qd1_hd r_mult_3_A_reg_27_ ( .D(n2477), .CK(n2252), .RN(n1104), .Q(
        r_mult_3_A[27]) );
  fd2qd1_hd r_mult_3_A_reg_26_ ( .D(n2476), .CK(n2252), .RN(n1424), .Q(
        r_mult_3_A[26]) );
  fd2qd1_hd r_mult_3_A_reg_25_ ( .D(n2476), .CK(n2252), .RN(n895), .Q(
        r_mult_3_A[25]) );
  fd2qd1_hd r_mult_3_A_reg_22_ ( .D(n2476), .CK(n2252), .RN(n1424), .Q(
        r_mult_3_A[22]) );
  fd2qd1_hd r_mult_3_A_reg_17_ ( .D(n2477), .CK(n2252), .RN(n1447), .Q(
        r_mult_3_A[17]) );
  fd2qd1_hd r_mult_3_A_reg_12_ ( .D(n2477), .CK(n2252), .RN(n1353), .Q(
        r_mult_3_A[12]) );
  fd2qd1_hd r_mult_3_A_reg_7_ ( .D(n2476), .CK(n2252), .RN(n1424), .Q(
        r_mult_3_A[7]) );
  fd2qd1_hd r_mult_3_A_reg_5_ ( .D(n2477), .CK(n2252), .RN(n1468), .Q(
        r_mult_3_A[5]) );
  fd2qd1_hd r_mult_3_A_reg_4_ ( .D(n2477), .CK(n2252), .RN(n1461), .Q(
        r_mult_3_A[4]) );
  fd2qd1_hd r_mult_3_A_reg_3_ ( .D(n2476), .CK(n2252), .RN(n1097), .Q(
        r_mult_3_A[3]) );
  fd2qd1_hd r_mult_2_A_reg_29_ ( .D(n2476), .CK(n2249), .RN(n1434), .Q(
        r_mult_2_A[29]) );
  fd2qd1_hd r_mult_2_A_reg_28_ ( .D(n2476), .CK(n2249), .RN(n889), .Q(
        r_mult_2_A[28]) );
  fd2qd1_hd r_mult_2_A_reg_27_ ( .D(n2477), .CK(n2249), .RN(n1458), .Q(
        r_mult_2_A[27]) );
  fd2qd1_hd r_mult_2_A_reg_26_ ( .D(n2477), .CK(n2249), .RN(n893), .Q(
        r_mult_2_A[26]) );
  fd2qd1_hd r_mult_2_A_reg_25_ ( .D(n2477), .CK(n2249), .RN(n1446), .Q(
        r_mult_2_A[25]) );
  fd2qd1_hd r_mult_2_A_reg_22_ ( .D(n2477), .CK(n2249), .RN(n895), .Q(
        r_mult_2_A[22]) );
  fd2qd1_hd r_mult_2_A_reg_10_ ( .D(n2476), .CK(n2249), .RN(n899), .Q(
        r_mult_2_A[10]) );
  fd2qd1_hd r_mult_2_A_reg_8_ ( .D(n2477), .CK(n2249), .RN(n1394), .Q(
        r_mult_2_A[8]) );
  fd2qd1_hd r_mult_2_A_reg_6_ ( .D(n2476), .CK(n2249), .RN(n1424), .Q(
        r_mult_2_A[6]) );
  fd2qd1_hd r_mult_2_A_reg_3_ ( .D(n2477), .CK(n2249), .RN(n1466), .Q(
        r_mult_2_A[3]) );
  fd2qd1_hd R_5 ( .D(n1518), .CK(n2249), .RN(n1466), .Q(n2243) );
  fd2qd1_hd R_1 ( .D(n1518), .CK(n2252), .RN(n888), .Q(n2247) );
  fd2qd1_hd R_8 ( .D(n2712), .CK(n2249), .RN(n308), .Q(n2240) );
  fd2qd1_hd r_mult_1_A_reg_31_ ( .D(n2678), .CK(n2249), .RN(n1443), .Q(
        r_mult_1_A[31]) );
  fd2qd1_hd r_mult_1_A_reg_30_ ( .D(n2677), .CK(n2249), .RN(n1442), .Q(
        r_mult_1_A[30]) );
  fd2qd1_hd r_mult_1_A_reg_20_ ( .D(n2665), .CK(n2249), .RN(n1463), .Q(
        r_mult_1_A[20]) );
  fd2qd1_hd r_mult_1_A_reg_16_ ( .D(n2661), .CK(n2249), .RN(n1073), .Q(
        r_mult_1_A[16]) );
  fd2qd1_hd r_mult_1_A_reg_12_ ( .D(n2657), .CK(n2249), .RN(n1341), .Q(
        r_mult_1_A[12]) );
  fd2qd1_hd r_mult_1_A_reg_9_ ( .D(n2654), .CK(n2249), .RN(n1447), .Q(
        r_mult_1_A[9]) );
  fd2qd1_hd r_mult_1_A_reg_8_ ( .D(n2653), .CK(n2249), .RN(n1394), .Q(
        r_mult_1_A[8]) );
  fd2qd1_hd r_mult_1_A_reg_6_ ( .D(n2651), .CK(n2249), .RN(n1207), .Q(
        r_mult_1_A[6]) );
  fd2qd1_hd r_mult_1_A_reg_1_ ( .D(n2646), .CK(n2249), .RN(n1424), .Q(
        r_mult_1_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_23_ ( .D(n2668), .CK(n2249), .RN(n1466), .Q(
        r_mult_1_A[23]) );
  fd2qd1_hd r_mult_1_A_reg_19_ ( .D(n2664), .CK(n2249), .RN(n1458), .Q(
        r_mult_1_A[19]) );
  fd2qd1_hd r_mult_1_A_reg_14_ ( .D(n2659), .CK(n2249), .RN(n1370), .Q(
        r_mult_1_A[14]) );
  fd2qd1_hd r_mult_1_A_reg_13_ ( .D(n2658), .CK(n2249), .RN(n1021), .Q(
        r_mult_1_A[13]) );
  fd2qd1_hd r_mult_1_A_reg_5_ ( .D(n2650), .CK(n2249), .RN(n1021), .Q(
        r_mult_1_A[5]) );
  fd2qd1_hd r_mult_1_A_reg_0_ ( .D(n2645), .CK(n2249), .RN(n1353), .Q(
        r_mult_1_A[0]) );
  fd2qd1_hd r_mult_1_B_reg_20_ ( .D(n2699), .CK(n2249), .RN(n889), .Q(
        r_mult_1_B[20]) );
  fd2qd1_hd r_mult_1_B_reg_30_ ( .D(n2709), .CK(n2249), .RN(n1097), .Q(
        r_mult_1_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_22_ ( .D(n2701), .CK(n2249), .RN(n1097), .Q(
        r_mult_1_B[22]) );
  fd2qd1_hd r_mult_1_B_reg_21_ ( .D(n2700), .CK(n2249), .RN(n895), .Q(
        r_mult_1_B[21]) );
  fd2qd1_hd r_mult_1_B_reg_28_ ( .D(n2707), .CK(n2249), .RN(n1353), .Q(
        r_mult_1_B[28]) );
  fd2qd1_hd r_mult_1_B_reg_27_ ( .D(n2706), .CK(n2249), .RN(n1384), .Q(
        r_mult_1_B[27]) );
  fd2qd1_hd r_mult_1_B_reg_26_ ( .D(n2705), .CK(n2249), .RN(n1353), .Q(
        r_mult_1_B[26]) );
  fd2qd1_hd r_mult_1_B_reg_25_ ( .D(n2704), .CK(n2249), .RN(n1401), .Q(
        r_mult_1_B[25]) );
  fd2qd1_hd r_mult_1_B_reg_24_ ( .D(n2703), .CK(n2249), .RN(n1104), .Q(
        r_mult_1_B[24]) );
  fd2qd1_hd r_mult_1_B_reg_23_ ( .D(n2702), .CK(n2249), .RN(n962), .Q(
        r_mult_1_B[23]) );
  fd2qd1_hd r_mult_3_B_reg_31_ ( .D(n2482), .CK(n2252), .RN(n1458), .Q(
        r_mult_3_B[31]) );
  fd2qd1_hd r_mult_3_B_reg_30_ ( .D(n2507), .CK(n2252), .RN(n1443), .Q(
        r_mult_3_B[30]) );
  fd2qd1_hd r_mult_3_B_reg_29_ ( .D(n2506), .CK(n2252), .RN(n893), .Q(
        r_mult_3_B[29]) );
  fd2qd1_hd r_mult_3_B_reg_28_ ( .D(n2494), .CK(n2252), .RN(n962), .Q(
        r_mult_3_B[28]) );
  fd2qd1_hd r_mult_3_B_reg_27_ ( .D(n2505), .CK(n2252), .RN(n1021), .Q(
        r_mult_3_B[27]) );
  fd2qd1_hd r_mult_3_B_reg_26_ ( .D(n2504), .CK(n2252), .RN(n893), .Q(
        r_mult_3_B[26]) );
  fd2qd1_hd r_mult_3_B_reg_25_ ( .D(n2503), .CK(n2252), .RN(n1463), .Q(
        r_mult_3_B[25]) );
  fd2qd1_hd r_mult_3_B_reg_24_ ( .D(n2502), .CK(n2252), .RN(n1370), .Q(
        r_mult_3_B[24]) );
  fd2qd1_hd r_mult_3_B_reg_23_ ( .D(n2493), .CK(n2252), .RN(n308), .Q(
        r_mult_3_B[23]) );
  fd2qd1_hd r_mult_3_B_reg_21_ ( .D(n2492), .CK(n2252), .RN(n1384), .Q(
        r_mult_3_B[21]) );
  fd2qd1_hd r_mult_3_B_reg_20_ ( .D(n2501), .CK(n2252), .RN(n1021), .Q(
        r_mult_3_B[20]) );
  fd2qd1_hd r_mult_3_B_reg_19_ ( .D(n2491), .CK(n2252), .RN(n1073), .Q(
        r_mult_3_B[19]) );
  fd2qd1_hd r_mult_3_B_reg_18_ ( .D(n2490), .CK(n2252), .RN(n1097), .Q(
        r_mult_3_B[18]) );
  fd2qd1_hd r_mult_3_B_reg_17_ ( .D(n2489), .CK(n2252), .RN(n964), .Q(
        r_mult_3_B[17]) );
  fd2qd1_hd r_mult_3_B_reg_16_ ( .D(n2500), .CK(n2252), .RN(n1458), .Q(
        r_mult_3_B[16]) );
  fd2qd1_hd r_mult_3_B_reg_14_ ( .D(n2488), .CK(n2252), .RN(n1401), .Q(
        r_mult_3_B[14]) );
  fd2qd1_hd r_mult_3_B_reg_13_ ( .D(n2487), .CK(n2252), .RN(n302), .Q(
        r_mult_3_B[13]) );
  fd2qd1_hd r_mult_3_B_reg_12_ ( .D(n2486), .CK(n2252), .RN(n1101), .Q(
        r_mult_3_B[12]) );
  fd2qd1_hd r_mult_3_B_reg_11_ ( .D(n2485), .CK(n2252), .RN(n1384), .Q(
        r_mult_3_B[11]) );
  fd2qd1_hd r_mult_3_B_reg_10_ ( .D(n2484), .CK(n2252), .RN(n1401), .Q(
        r_mult_3_B[10]) );
  fd2qd1_hd r_mult_3_B_reg_9_ ( .D(n2499), .CK(n2252), .RN(n1384), .Q(
        r_mult_3_B[9]) );
  fd2qd1_hd r_mult_3_B_reg_8_ ( .D(n2498), .CK(n2252), .RN(n889), .Q(
        r_mult_3_B[8]) );
  fd2qd1_hd r_mult_3_B_reg_7_ ( .D(n2497), .CK(n2252), .RN(n1372), .Q(
        r_mult_3_B[7]) );
  fd2qd1_hd r_mult_3_B_reg_5_ ( .D(n2496), .CK(n2252), .RN(n1097), .Q(
        r_mult_3_B[5]) );
  fd2qd1_hd r_mult_3_B_reg_3_ ( .D(n2495), .CK(n2252), .RN(n1021), .Q(
        r_mult_3_B[3]) );
  fd2qd1_hd r_mult_3_B_reg_1_ ( .D(n2483), .CK(n2252), .RN(n1471), .Q(
        r_mult_3_B[1]) );
  fd2qd1_hd r_mult_3_B_reg_6_ ( .D(n2481), .CK(n2252), .RN(n889), .Q(
        r_mult_3_B[6]) );
  fd2qd1_hd r_mult_3_B_reg_4_ ( .D(n2480), .CK(n2252), .RN(n1073), .Q(
        r_mult_3_B[4]) );
  fd2qd1_hd r_mult_3_B_reg_2_ ( .D(n2479), .CK(n2252), .RN(n1401), .Q(
        r_mult_3_B[2]) );
  fd2qd1_hd r_mult_3_B_reg_0_ ( .D(n2478), .CK(n2252), .RN(n302), .Q(
        r_mult_3_B[0]) );
  fd2qd1_hd r_mult_2_B_reg_30_ ( .D(n2743), .CK(n2249), .RN(n1384), .Q(
        r_mult_2_B[30]) );
  fd2qd1_hd r_mult_2_B_reg_26_ ( .D(n2739), .CK(n2249), .RN(n1353), .Q(
        r_mult_2_B[26]) );
  fd2qd1_hd r_mult_2_B_reg_25_ ( .D(n2738), .CK(n2249), .RN(n1101), .Q(
        r_mult_2_B[25]) );
  fd2qd1_hd r_mult_2_B_reg_22_ ( .D(n2735), .CK(n2249), .RN(n1443), .Q(
        r_mult_2_B[22]) );
  fd2qd1_hd r_mult_2_B_reg_20_ ( .D(n2733), .CK(n2249), .RN(n962), .Q(
        r_mult_2_B[20]) );
  fd2qd1_hd r_mult_2_B_reg_18_ ( .D(n2731), .CK(n2249), .RN(n308), .Q(
        r_mult_2_B[18]) );
  fd2qd1_hd r_mult_2_B_reg_15_ ( .D(n2728), .CK(n2249), .RN(n888), .Q(
        r_mult_2_B[15]) );
  fd2qd1_hd r_mult_2_B_reg_14_ ( .D(n2727), .CK(n2249), .RN(n1466), .Q(
        r_mult_2_B[14]) );
  fd2qd1_hd r_mult_2_B_reg_12_ ( .D(n2725), .CK(n2249), .RN(n308), .Q(
        r_mult_2_B[12]) );
  fd2qd1_hd r_mult_2_B_reg_10_ ( .D(n2723), .CK(n2249), .RN(n964), .Q(
        r_mult_2_B[10]) );
  fd2qd1_hd r_mult_2_B_reg_9_ ( .D(n2722), .CK(n2249), .RN(n1370), .Q(
        r_mult_2_B[9]) );
  fd2qd1_hd r_mult_2_B_reg_6_ ( .D(n2719), .CK(n2249), .RN(n888), .Q(
        r_mult_2_B[6]) );
  fd2qd1_hd r_mult_2_B_reg_5_ ( .D(n2718), .CK(n2249), .RN(n899), .Q(
        r_mult_2_B[5]) );
  fd2qd1_hd r_mult_2_B_reg_4_ ( .D(n2717), .CK(n2249), .RN(n888), .Q(
        r_mult_2_B[4]) );
  fd2qd1_hd r_mult_2_B_reg_2_ ( .D(n2715), .CK(n2249), .RN(n1447), .Q(
        r_mult_2_B[2]) );
  fd2qd1_hd r_mult_2_B_reg_1_ ( .D(n2714), .CK(n2249), .RN(n1372), .Q(
        r_mult_2_B[1]) );
  fd2qd1_hd r_mult_2_B_reg_0_ ( .D(n2713), .CK(n2249), .RN(n1434), .Q(
        r_mult_2_B[0]) );
  fd2qd1_hd r_mult_1_B_reg_31_ ( .D(n2710), .CK(n2249), .RN(n1101), .Q(
        r_mult_1_B[31]) );
  fd2qd1_hd r_mult_2_B_reg_31_ ( .D(n2744), .CK(n2249), .RN(n302), .Q(
        r_mult_2_B[31]) );
  fd2qd1_hd r_mult_2_B_reg_29_ ( .D(n2742), .CK(n2249), .RN(n938), .Q(
        r_mult_2_B[29]) );
  fd2qd1_hd r_mult_2_B_reg_28_ ( .D(n2741), .CK(n2249), .RN(n1384), .Q(
        r_mult_2_B[28]) );
  fd2qd1_hd r_mult_2_B_reg_27_ ( .D(n2740), .CK(n2249), .RN(n1235), .Q(
        r_mult_2_B[27]) );
  fd2qd1_hd r_mult_2_B_reg_24_ ( .D(n2737), .CK(n2249), .RN(n1468), .Q(
        r_mult_2_B[24]) );
  fd2qd1_hd r_mult_2_B_reg_23_ ( .D(n2736), .CK(n2249), .RN(n1117), .Q(
        r_mult_2_B[23]) );
  fd2qd1_hd r_mult_2_B_reg_21_ ( .D(n2734), .CK(n2249), .RN(n1420), .Q(
        r_mult_2_B[21]) );
  fd2qd1_hd r_mult_2_B_reg_19_ ( .D(n2732), .CK(n2249), .RN(n962), .Q(
        r_mult_2_B[19]) );
  fd2qd1_hd r_mult_2_B_reg_17_ ( .D(n2730), .CK(n2249), .RN(n1062), .Q(
        r_mult_2_B[17]) );
  fd2qd1_hd r_mult_2_B_reg_16_ ( .D(n2729), .CK(n2249), .RN(n1442), .Q(
        r_mult_2_B[16]) );
  fd2qd1_hd r_mult_2_B_reg_13_ ( .D(n2726), .CK(n2249), .RN(n1458), .Q(
        r_mult_2_B[13]) );
  fd2qd1_hd r_mult_2_B_reg_8_ ( .D(n2721), .CK(n2249), .RN(n1353), .Q(
        r_mult_2_B[8]) );
  fd2qd1_hd r_mult_2_B_reg_7_ ( .D(n2720), .CK(n2249), .RN(n888), .Q(
        r_mult_2_B[7]) );
  fd2qd1_hd r_mult_2_B_reg_3_ ( .D(n2716), .CK(n2249), .RN(n962), .Q(
        r_mult_2_B[3]) );
  fd2qd1_hd r_counter_reg_1_ ( .D(n841), .CK(n2255), .RN(n1401), .Q(
        r_counter[1]) );
  fd2qd1_hd r_add_1_B_reg_0_ ( .D(n2545), .CK(n2251), .RN(n1471), .Q(
        r_add_1_B[0]) );
  fd2qd1_hd r_add_1_A_reg_0_ ( .D(n2512), .CK(n2251), .RN(n1471), .Q(
        r_add_1_A[0]) );
  fd2qd1_hd r_add_1_B_reg_31_ ( .D(n2576), .CK(n2251), .RN(n1550), .Q(
        r_add_1_B[31]) );
  fd2qd1_hd r_add_1_B_reg_30_ ( .D(n2575), .CK(n2251), .RN(n1420), .Q(
        r_add_1_B[30]) );
  fd2qd1_hd r_add_1_B_reg_29_ ( .D(n2574), .CK(n2251), .RN(n1424), .Q(
        r_add_1_B[29]) );
  fd2qd1_hd r_add_1_B_reg_28_ ( .D(n2573), .CK(n2251), .RN(n1424), .Q(
        r_add_1_B[28]) );
  fd2qd1_hd r_add_1_B_reg_27_ ( .D(n2572), .CK(n2251), .RN(n1471), .Q(
        r_add_1_B[27]) );
  fd2qd1_hd r_add_1_B_reg_26_ ( .D(n2571), .CK(n2251), .RN(n1431), .Q(
        r_add_1_B[26]) );
  fd2qd1_hd r_add_1_B_reg_25_ ( .D(n2570), .CK(n2251), .RN(n1097), .Q(
        r_add_1_B[25]) );
  fd2qd1_hd r_add_1_B_reg_24_ ( .D(n2569), .CK(n2251), .RN(n1073), .Q(
        r_add_1_B[24]) );
  fd2qd1_hd r_add_1_B_reg_23_ ( .D(n2568), .CK(n2251), .RN(n893), .Q(
        r_add_1_B[23]) );
  fd2qd1_hd r_add_1_B_reg_22_ ( .D(n2567), .CK(n2251), .RN(n1370), .Q(
        r_add_1_B[22]) );
  fd2qd1_hd r_add_1_B_reg_21_ ( .D(n2566), .CK(n2251), .RN(n1431), .Q(
        r_add_1_B[21]) );
  fd2qd1_hd r_add_1_B_reg_20_ ( .D(n2565), .CK(n2251), .RN(n938), .Q(
        r_add_1_B[20]) );
  fd2qd1_hd r_add_1_B_reg_19_ ( .D(n2564), .CK(n2251), .RN(n964), .Q(
        r_add_1_B[19]) );
  fd2qd1_hd r_add_1_B_reg_18_ ( .D(n2563), .CK(n2251), .RN(n1434), .Q(
        r_add_1_B[18]) );
  fd2qd1_hd r_add_1_B_reg_17_ ( .D(n2562), .CK(n2251), .RN(n1353), .Q(
        r_add_1_B[17]) );
  fd2qd1_hd r_add_1_B_reg_16_ ( .D(n2561), .CK(n2251), .RN(n1424), .Q(
        r_add_1_B[16]) );
  fd2qd1_hd r_add_1_B_reg_15_ ( .D(n2560), .CK(n2251), .RN(n1424), .Q(
        r_add_1_B[15]) );
  fd2qd1_hd r_add_1_B_reg_14_ ( .D(n2559), .CK(n2251), .RN(n1420), .Q(
        r_add_1_B[14]) );
  fd2qd1_hd r_add_1_B_reg_13_ ( .D(n2558), .CK(n2251), .RN(n1394), .Q(
        r_add_1_B[13]) );
  fd2qd1_hd r_add_1_B_reg_12_ ( .D(n2557), .CK(n2251), .RN(n1443), .Q(
        r_add_1_B[12]) );
  fd2qd1_hd r_add_1_B_reg_11_ ( .D(n2556), .CK(n2251), .RN(n895), .Q(
        r_add_1_B[11]) );
  fd2qd1_hd r_add_1_B_reg_10_ ( .D(n2555), .CK(n2251), .RN(n1442), .Q(
        r_add_1_B[10]) );
  fd2qd1_hd r_add_1_B_reg_9_ ( .D(n2554), .CK(n2251), .RN(n1443), .Q(
        r_add_1_B[9]) );
  fd2qd1_hd r_add_1_B_reg_8_ ( .D(n2553), .CK(n2251), .RN(n895), .Q(
        r_add_1_B[8]) );
  fd2qd1_hd r_add_1_B_reg_7_ ( .D(n2552), .CK(n2251), .RN(n899), .Q(
        r_add_1_B[7]) );
  fd2qd1_hd r_add_1_B_reg_6_ ( .D(n2551), .CK(n2251), .RN(n1446), .Q(
        r_add_1_B[6]) );
  fd2qd1_hd r_add_1_B_reg_5_ ( .D(n2550), .CK(n2251), .RN(n1447), .Q(
        r_add_1_B[5]) );
  fd2qd1_hd r_add_1_B_reg_4_ ( .D(n2549), .CK(n2251), .RN(n1341), .Q(
        r_add_1_B[4]) );
  fd2qd1_hd r_add_1_B_reg_3_ ( .D(n2548), .CK(n2251), .RN(n1471), .Q(
        r_add_1_B[3]) );
  fd2qd1_hd r_add_1_B_reg_2_ ( .D(n2547), .CK(n2251), .RN(n1235), .Q(
        r_add_1_B[2]) );
  fd2qd1_hd r_add_1_B_reg_1_ ( .D(n2546), .CK(n2251), .RN(n1235), .Q(
        r_add_1_B[1]) );
  fd2qd1_hd r_add_1_A_reg_31_ ( .D(n2543), .CK(n2251), .RN(n1235), .Q(
        r_add_1_A[31]) );
  fd2qd1_hd r_add_1_A_reg_30_ ( .D(n2542), .CK(n2251), .RN(n888), .Q(
        r_add_1_A[30]) );
  fd2qd1_hd r_add_1_A_reg_29_ ( .D(n2541), .CK(n2251), .RN(n888), .Q(
        r_add_1_A[29]) );
  fd2qd1_hd r_add_1_A_reg_28_ ( .D(n2540), .CK(n2251), .RN(n1370), .Q(
        r_add_1_A[28]) );
  fd2qd1_hd r_add_1_A_reg_27_ ( .D(n2539), .CK(n2251), .RN(n1458), .Q(
        r_add_1_A[27]) );
  fd2qd1_hd r_add_1_A_reg_26_ ( .D(n2538), .CK(n2251), .RN(n1458), .Q(
        r_add_1_A[26]) );
  fd2qd1_hd r_add_1_A_reg_25_ ( .D(n2537), .CK(n2251), .RN(n1117), .Q(
        r_add_1_A[25]) );
  fd2qd1_hd r_add_1_A_reg_24_ ( .D(n2536), .CK(n2251), .RN(n1461), .Q(
        r_add_1_A[24]) );
  fd2qd1_hd r_add_1_A_reg_23_ ( .D(n2535), .CK(n2251), .RN(n1461), .Q(
        r_add_1_A[23]) );
  fd2qd1_hd r_add_1_A_reg_22_ ( .D(n2534), .CK(n2251), .RN(n1463), .Q(
        r_add_1_A[22]) );
  fd2qd1_hd r_add_1_A_reg_21_ ( .D(n2533), .CK(n2251), .RN(n1463), .Q(
        r_add_1_A[21]) );
  fd2qd1_hd r_add_1_A_reg_20_ ( .D(n2532), .CK(n2251), .RN(n1353), .Q(
        r_add_1_A[20]) );
  fd2qd1_hd r_add_1_A_reg_19_ ( .D(n2531), .CK(n2251), .RN(n1466), .Q(
        r_add_1_A[19]) );
  fd2qd1_hd r_add_1_A_reg_18_ ( .D(n2530), .CK(n2251), .RN(n1466), .Q(
        r_add_1_A[18]) );
  fd2qd1_hd r_add_1_A_reg_17_ ( .D(n2529), .CK(n2251), .RN(n1468), .Q(
        r_add_1_A[17]) );
  fd2qd1_hd r_add_1_A_reg_16_ ( .D(n2528), .CK(n2251), .RN(n1468), .Q(
        r_add_1_A[16]) );
  fd2qd1_hd r_add_1_A_reg_15_ ( .D(n2527), .CK(n2251), .RN(n888), .Q(
        r_add_1_A[15]) );
  fd2qd1_hd r_add_1_A_reg_14_ ( .D(n2526), .CK(n2251), .RN(n1471), .Q(
        r_add_1_A[14]) );
  fd2qd1_hd r_add_1_A_reg_13_ ( .D(n2525), .CK(n2251), .RN(n1471), .Q(
        r_add_1_A[13]) );
  fd2qd1_hd r_add_1_A_reg_12_ ( .D(n2524), .CK(n2251), .RN(n1021), .Q(
        r_add_1_A[12]) );
  fd2qd1_hd r_add_1_A_reg_11_ ( .D(n2523), .CK(n2251), .RN(n308), .Q(
        r_add_1_A[11]) );
  fd2qd1_hd r_add_1_A_reg_10_ ( .D(n2522), .CK(n2251), .RN(n1394), .Q(
        r_add_1_A[10]) );
  fd2qd1_hd r_add_1_A_reg_9_ ( .D(n2521), .CK(n2251), .RN(n895), .Q(
        r_add_1_A[9]) );
  fd2qd1_hd r_add_1_A_reg_8_ ( .D(n2520), .CK(n2251), .RN(n1550), .Q(
        r_add_1_A[8]) );
  fd2qd1_hd r_add_1_A_reg_7_ ( .D(n2519), .CK(n2251), .RN(n1117), .Q(
        r_add_1_A[7]) );
  fd2qd1_hd r_add_1_A_reg_6_ ( .D(n2518), .CK(n2251), .RN(n1550), .Q(
        r_add_1_A[6]) );
  fd2qd1_hd r_add_1_A_reg_5_ ( .D(n2517), .CK(n2251), .RN(n1442), .Q(
        r_add_1_A[5]) );
  fd2qd1_hd r_add_1_A_reg_4_ ( .D(n2516), .CK(n2251), .RN(n1447), .Q(
        r_add_1_A[4]) );
  fd2qd1_hd r_add_1_A_reg_3_ ( .D(n2515), .CK(n2251), .RN(n1550), .Q(
        r_add_1_A[3]) );
  fd2qd1_hd r_add_1_A_reg_2_ ( .D(n2514), .CK(n2251), .RN(n899), .Q(
        r_add_1_A[2]) );
  fd2qd1_hd r_add_1_A_reg_1_ ( .D(n2513), .CK(n2251), .RN(n1550), .Q(
        r_add_1_A[1]) );
  fd2qd1_hd r_add_2_A_reg_31_ ( .D(n2610), .CK(n2250), .RN(n1401), .Q(
        r_add_2_A[31]) );
  fd2qd1_hd r_add_2_A_reg_30_ ( .D(n2609), .CK(n2250), .RN(n1062), .Q(
        r_add_2_A[30]) );
  fd2qd1_hd r_add_2_A_reg_29_ ( .D(n2608), .CK(n2250), .RN(n1235), .Q(
        r_add_2_A[29]) );
  fd2qd1_hd r_add_2_A_reg_28_ ( .D(n2607), .CK(n2250), .RN(n964), .Q(
        r_add_2_A[28]) );
  fd2qd1_hd r_add_2_A_reg_27_ ( .D(n2606), .CK(n2250), .RN(n1471), .Q(
        r_add_2_A[27]) );
  fd2qd1_hd r_add_2_A_reg_26_ ( .D(n2605), .CK(n2250), .RN(n1442), .Q(
        r_add_2_A[26]) );
  fd2qd1_hd r_add_2_A_reg_25_ ( .D(n2604), .CK(n2250), .RN(n1394), .Q(
        r_add_2_A[25]) );
  fd2qd1_hd r_add_2_A_reg_24_ ( .D(n2603), .CK(n2250), .RN(n1458), .Q(
        r_add_2_A[24]) );
  fd2qd1_hd r_add_2_A_reg_23_ ( .D(n2602), .CK(n2250), .RN(n893), .Q(
        r_add_2_A[23]) );
  fd2qd1_hd r_add_2_A_reg_22_ ( .D(n2601), .CK(n2250), .RN(n888), .Q(
        r_add_2_A[22]) );
  fd2qd1_hd r_add_2_A_reg_21_ ( .D(n2600), .CK(n2250), .RN(n1101), .Q(
        r_add_2_A[21]) );
  fd2qd1_hd r_add_2_A_reg_20_ ( .D(n2599), .CK(n2250), .RN(n888), .Q(
        r_add_2_A[20]) );
  fd2qd1_hd r_add_2_A_reg_19_ ( .D(n2598), .CK(n2250), .RN(n1062), .Q(
        r_add_2_A[19]) );
  fd2qd1_hd r_add_2_A_reg_18_ ( .D(n2597), .CK(n2250), .RN(n1401), .Q(
        r_add_2_A[18]) );
  fd2qd1_hd r_add_2_A_reg_17_ ( .D(n2596), .CK(n2250), .RN(n302), .Q(
        r_add_2_A[17]) );
  fd2qd1_hd r_add_2_A_reg_16_ ( .D(n2595), .CK(n2250), .RN(n1458), .Q(
        r_add_2_A[16]) );
  fd2qd1_hd r_add_2_A_reg_15_ ( .D(n2594), .CK(n2250), .RN(n1062), .Q(
        r_add_2_A[15]) );
  fd2qd1_hd r_add_2_A_reg_14_ ( .D(n2593), .CK(n2250), .RN(n895), .Q(
        r_add_2_A[14]) );
  fd2qd1_hd r_add_2_A_reg_13_ ( .D(n2592), .CK(n2250), .RN(n308), .Q(
        r_add_2_A[13]) );
  fd2qd1_hd r_add_2_A_reg_12_ ( .D(n2591), .CK(n2250), .RN(n1235), .Q(
        r_add_2_A[12]) );
  fd2qd1_hd r_add_2_A_reg_11_ ( .D(n2590), .CK(n2250), .RN(n938), .Q(
        r_add_2_A[11]) );
  fd2qd1_hd r_add_2_A_reg_10_ ( .D(n2589), .CK(n2250), .RN(n1468), .Q(
        r_add_2_A[10]) );
  fd2qd1_hd r_add_2_A_reg_9_ ( .D(n2588), .CK(n2250), .RN(n1401), .Q(
        r_add_2_A[9]) );
  fd2qd1_hd r_add_2_A_reg_8_ ( .D(n2587), .CK(n2250), .RN(n1207), .Q(
        r_add_2_A[8]) );
  fd2qd1_hd r_add_2_A_reg_7_ ( .D(n2586), .CK(n2250), .RN(n1431), .Q(
        r_add_2_A[7]) );
  fd2qd1_hd r_add_2_A_reg_6_ ( .D(n2585), .CK(n2250), .RN(n1550), .Q(
        r_add_2_A[6]) );
  fd2qd1_hd r_add_2_A_reg_5_ ( .D(n2584), .CK(n2250), .RN(n1461), .Q(
        r_add_2_A[5]) );
  fd2qd1_hd r_add_2_A_reg_4_ ( .D(n2583), .CK(n2250), .RN(n962), .Q(
        r_add_2_A[4]) );
  fd2qd1_hd r_add_2_A_reg_3_ ( .D(n2582), .CK(n2250), .RN(n964), .Q(
        r_add_2_A[3]) );
  fd2qd1_hd r_add_2_A_reg_2_ ( .D(n2581), .CK(n2250), .RN(n938), .Q(
        r_add_2_A[2]) );
  fd2qd1_hd r_add_2_A_reg_1_ ( .D(n2580), .CK(n2250), .RN(n1461), .Q(
        r_add_2_A[1]) );
  fd2qd1_hd r_add_2_A_reg_0_ ( .D(n2579), .CK(n2250), .RN(n1446), .Q(
        r_add_2_A[0]) );
  fd2qd1_hd r_add_2_B_reg_0_ ( .D(n2611), .CK(n2250), .RN(n899), .Q(
        r_add_2_B[0]) );
  fd2qd1_hd r_mult_1_A_reg_29_ ( .D(n2674), .CK(n2249), .RN(n1424), .Q(
        r_mult_1_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_28_ ( .D(n2673), .CK(n2249), .RN(n1443), .Q(
        r_mult_1_A[28]) );
  fd2qd1_hd r_mult_1_A_reg_27_ ( .D(n2672), .CK(n2249), .RN(n1442), .Q(
        r_mult_1_A[27]) );
  fd2qd1_hd r_mult_1_A_reg_26_ ( .D(n2671), .CK(n2249), .RN(n893), .Q(
        r_mult_1_A[26]) );
  fd2qd1_hd r_mult_1_A_reg_25_ ( .D(n2670), .CK(n2249), .RN(n1463), .Q(
        r_mult_1_A[25]) );
  fd2qd1_hd r_mult_1_A_reg_24_ ( .D(n2669), .CK(n2249), .RN(n1394), .Q(
        r_mult_1_A[24]) );
  fd2qd1_hd r_mult_1_A_reg_22_ ( .D(n2667), .CK(n2249), .RN(n1104), .Q(
        r_mult_1_A[22]) );
  fd2qd1_hd r_mult_1_A_reg_21_ ( .D(n2666), .CK(n2249), .RN(n1471), .Q(
        r_mult_1_A[21]) );
  fd2qd1_hd r_mult_1_A_reg_7_ ( .D(n2652), .CK(n2249), .RN(n1463), .Q(
        r_mult_1_A[7]) );
  fd2qd1_hd r_mult_1_A_reg_3_ ( .D(n2648), .CK(n2249), .RN(n1370), .Q(
        r_mult_1_A[3]) );
  fd2qd1_hd r_add_2_B_reg_31_ ( .D(n2642), .CK(n2250), .RN(n1101), .Q(
        r_add_2_B[31]) );
  fd2qd1_hd r_add_2_B_reg_30_ ( .D(n2641), .CK(n2250), .RN(n1434), .Q(
        r_add_2_B[30]) );
  fd2qd1_hd r_add_2_B_reg_29_ ( .D(n2640), .CK(n2250), .RN(n1443), .Q(
        r_add_2_B[29]) );
  fd2qd1_hd r_add_2_B_reg_28_ ( .D(n2639), .CK(n2250), .RN(n1447), .Q(
        r_add_2_B[28]) );
  fd2qd1_hd r_add_2_B_reg_27_ ( .D(n2638), .CK(n2250), .RN(n1446), .Q(
        r_add_2_B[27]) );
  fd2qd1_hd r_add_2_B_reg_26_ ( .D(n2637), .CK(n2250), .RN(n1447), .Q(
        r_add_2_B[26]) );
  fd2qd1_hd r_add_2_B_reg_25_ ( .D(n2636), .CK(n2250), .RN(n1420), .Q(
        r_add_2_B[25]) );
  fd2qd1_hd r_add_2_B_reg_24_ ( .D(n2635), .CK(n2250), .RN(n1443), .Q(
        r_add_2_B[24]) );
  fd2qd1_hd r_add_2_B_reg_23_ ( .D(n2634), .CK(n2250), .RN(n1442), .Q(
        r_add_2_B[23]) );
  fd2qd1_hd r_add_2_B_reg_22_ ( .D(n2633), .CK(n2250), .RN(n1463), .Q(
        r_add_2_B[22]) );
  fd2qd1_hd r_add_2_B_reg_21_ ( .D(n2632), .CK(n2250), .RN(n1466), .Q(
        r_add_2_B[21]) );
  fd2qd1_hd r_add_2_B_reg_20_ ( .D(n2631), .CK(n2250), .RN(n1394), .Q(
        r_add_2_B[20]) );
  fd2qd1_hd r_add_2_B_reg_19_ ( .D(n2630), .CK(n2250), .RN(n889), .Q(
        r_add_2_B[19]) );
  fd2qd1_hd r_add_2_B_reg_18_ ( .D(n2629), .CK(n2250), .RN(n1372), .Q(
        r_add_2_B[18]) );
  fd2qd1_hd r_add_2_B_reg_17_ ( .D(n2628), .CK(n2250), .RN(n1370), .Q(
        r_add_2_B[17]) );
  fd2qd1_hd r_add_2_B_reg_16_ ( .D(n2627), .CK(n2250), .RN(n1394), .Q(
        r_add_2_B[16]) );
  fd2qd1_hd r_add_2_B_reg_15_ ( .D(n2626), .CK(n2250), .RN(n1372), .Q(
        r_add_2_B[15]) );
  fd2qd1_hd r_add_2_B_reg_14_ ( .D(n2625), .CK(n2250), .RN(n1442), .Q(
        r_add_2_B[14]) );
  fd2qd1_hd r_add_2_B_reg_13_ ( .D(n2624), .CK(n2250), .RN(n1461), .Q(
        r_add_2_B[13]) );
  fd2qd1_hd r_add_2_B_reg_12_ ( .D(n2623), .CK(n2250), .RN(n1097), .Q(
        r_add_2_B[12]) );
  fd2qd1_hd r_add_2_B_reg_11_ ( .D(n2622), .CK(n2250), .RN(n1434), .Q(
        r_add_2_B[11]) );
  fd2qd1_hd r_add_2_B_reg_10_ ( .D(n2621), .CK(n2250), .RN(n1097), .Q(
        r_add_2_B[10]) );
  fd2qd1_hd r_add_2_B_reg_9_ ( .D(n2620), .CK(n2250), .RN(n1471), .Q(
        r_add_2_B[9]) );
  fd2qd1_hd r_add_2_B_reg_8_ ( .D(n2619), .CK(n2250), .RN(n1401), .Q(
        r_add_2_B[8]) );
  fd2qd1_hd r_add_2_B_reg_7_ ( .D(n2618), .CK(n2250), .RN(n1420), .Q(
        r_add_2_B[7]) );
  fd2qd1_hd r_add_2_B_reg_6_ ( .D(n2617), .CK(n2250), .RN(n1447), .Q(
        r_add_2_B[6]) );
  fd2qd1_hd r_add_2_B_reg_5_ ( .D(n2616), .CK(n2250), .RN(n1073), .Q(
        r_add_2_B[5]) );
  fd2qd1_hd r_add_2_B_reg_4_ ( .D(n2615), .CK(n2250), .RN(n938), .Q(
        r_add_2_B[4]) );
  fd2qd1_hd r_add_2_B_reg_3_ ( .D(n2614), .CK(n2250), .RN(n1384), .Q(
        r_add_2_B[3]) );
  fd2qd1_hd r_add_2_B_reg_2_ ( .D(n2613), .CK(n2250), .RN(n1341), .Q(
        r_add_2_B[2]) );
  fd2qd1_hd r_add_2_B_reg_1_ ( .D(n2612), .CK(n2250), .RN(n1101), .Q(
        r_add_2_B[1]) );
  fd2qd1_hd R_7 ( .D(n2239), .CK(i_CLK), .RN(n1097), .Q(n2241) );
  fd2qd1_hd r_add_2_Z_ACK_reg ( .D(n518), .CK(n2255), .RN(n1420), .Q(
        r_add_2_Z_ACK) );
  fd2qd1_hd r_mult_3_Z_ACK_reg ( .D(n2238), .CK(i_CLK), .RN(n1401), .Q(
        r_mult_3_Z_ACK) );
  fd2qd1_hd r_counter_reg_0_ ( .D(n844), .CK(n2255), .RN(n1394), .Q(
        r_counter[0]) );
  nr2bd1_hd U1 ( .AN(n1506), .B(n2234), .Y(n311) );
  ivd1_hd U2 ( .A(r_counter[2]), .Y(N44) );
  ivd1_hd U3 ( .A(n847), .Y(n851) );
  ivd1_hd U4 ( .A(n846), .Y(n850) );
  clknd2d1_hd U5 ( .A(r_pstate[1]), .B(n1509), .Y(n2262) );
  ivd2_hd U6 ( .A(r_counter[0]), .Y(N46) );
  clknd2d1_hd U8 ( .A(w_add_1_Z[31]), .B(n2236), .Y(n328) );
  nr2d1_hd U9 ( .A(N49), .B(N46), .Y(n1500) );
  ivd1_hd U11 ( .A(n845), .Y(n849) );
  ad2d1_hd U12 ( .A(n1510), .B(alt59_n135), .Y(N1406) );
  mx2d1_hd U13 ( .D0(r_mult_3_Z_ACK), .D1(n838), .S(n850), .Y(n2238) );
  clknd2d1_hd U14 ( .A(n846), .B(n1560), .Y(N1399) );
  mx2d1_hd U15 ( .D0(n2241), .D1(n2235), .S(n850), .Y(n2239) );
  mx2d1_hd U16 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[3]), .Y(n2648) );
  mx2d1_hd U17 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[7]), .Y(n2652) );
  mx2d1_hd U18 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[21]), .Y(n2666) );
  mx2d1_hd U19 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[22]), .Y(n2667) );
  mx2d1_hd U20 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[24]), .Y(n2669) );
  mx2d1_hd U21 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[25]), .Y(n2670) );
  mx2d1_hd U22 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[26]), .Y(n2671) );
  mx2d1_hd U23 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[27]), .Y(n2672) );
  mx2d1_hd U24 ( .D0(n2676), .D1(n2675), .S(w_mult_1_Z[28]), .Y(n2673) );
  scg2d1_hd U25 ( .A(n2237), .B(r_y_data[64]), .C(r_y_data[32]), .D(n1518), 
        .Y(n2478) );
  scg2d1_hd U26 ( .A(n2237), .B(r_y_data[66]), .C(r_y_data[34]), .D(n1518), 
        .Y(n2479) );
  scg2d1_hd U27 ( .A(n2237), .B(r_y_data[68]), .C(r_y_data[36]), .D(n1518), 
        .Y(n2480) );
  scg2d1_hd U28 ( .A(n2237), .B(r_y_data[70]), .C(r_y_data[38]), .D(n1518), 
        .Y(n2481) );
  scg2d1_hd U29 ( .A(n2235), .B(r_y_data[65]), .C(r_y_data[33]), .D(n1518), 
        .Y(n2483) );
  scg2d1_hd U30 ( .A(n2236), .B(r_y_data[67]), .C(r_y_data[35]), .D(n1518), 
        .Y(n2495) );
  scg2d1_hd U31 ( .A(n2236), .B(r_y_data[69]), .C(r_y_data[37]), .D(n1518), 
        .Y(n2496) );
  scg2d1_hd U32 ( .A(n2236), .B(r_y_data[71]), .C(r_y_data[39]), .D(n1518), 
        .Y(n2497) );
  scg2d1_hd U33 ( .A(n2236), .B(r_y_data[72]), .C(r_y_data[40]), .D(n1518), 
        .Y(n2498) );
  scg2d1_hd U34 ( .A(n2236), .B(r_y_data[73]), .C(r_y_data[41]), .D(n1518), 
        .Y(n2499) );
  scg2d1_hd U35 ( .A(n2236), .B(r_y_data[74]), .C(r_y_data[42]), .D(n1518), 
        .Y(n2484) );
  scg2d1_hd U36 ( .A(n2235), .B(r_y_data[75]), .C(r_y_data[43]), .D(n1518), 
        .Y(n2485) );
  scg2d1_hd U37 ( .A(n2236), .B(r_y_data[76]), .C(r_y_data[44]), .D(n1518), 
        .Y(n2486) );
  scg2d1_hd U38 ( .A(n2235), .B(r_y_data[77]), .C(r_y_data[45]), .D(n1518), 
        .Y(n2487) );
  scg2d1_hd U39 ( .A(n2236), .B(r_y_data[78]), .C(r_y_data[46]), .D(n1518), 
        .Y(n2488) );
  scg2d1_hd U40 ( .A(n2236), .B(r_y_data[80]), .C(r_y_data[48]), .D(n1518), 
        .Y(n2500) );
  scg2d1_hd U41 ( .A(n2235), .B(r_y_data[81]), .C(r_y_data[49]), .D(n1518), 
        .Y(n2489) );
  scg2d1_hd U42 ( .A(n2236), .B(r_y_data[82]), .C(r_y_data[50]), .D(n1518), 
        .Y(n2490) );
  scg2d1_hd U43 ( .A(n2236), .B(r_y_data[83]), .C(r_y_data[51]), .D(n1518), 
        .Y(n2491) );
  scg2d1_hd U44 ( .A(n2236), .B(r_y_data[84]), .C(r_y_data[52]), .D(n1518), 
        .Y(n2501) );
  scg2d1_hd U45 ( .A(n2236), .B(r_y_data[85]), .C(r_y_data[53]), .D(n1518), 
        .Y(n2492) );
  scg2d1_hd U46 ( .A(n2236), .B(r_y_data[87]), .C(r_y_data[55]), .D(n1518), 
        .Y(n2493) );
  scg2d1_hd U47 ( .A(n2236), .B(r_y_data[88]), .C(r_y_data[56]), .D(n1518), 
        .Y(n2502) );
  scg2d1_hd U48 ( .A(n2236), .B(r_y_data[89]), .C(r_y_data[57]), .D(n1518), 
        .Y(n2503) );
  scg2d1_hd U49 ( .A(n2236), .B(r_y_data[90]), .C(r_y_data[58]), .D(n1518), 
        .Y(n2504) );
  scg2d1_hd U50 ( .A(n2236), .B(r_y_data[91]), .C(r_y_data[59]), .D(n1518), 
        .Y(n2505) );
  scg2d1_hd U51 ( .A(n2236), .B(r_y_data[92]), .C(r_y_data[60]), .D(n1518), 
        .Y(n2494) );
  scg2d1_hd U54 ( .A(n2236), .B(r_y_data[93]), .C(r_y_data[61]), .D(n1518), 
        .Y(n2506) );
  scg2d1_hd U55 ( .A(n2236), .B(r_y_data[94]), .C(r_y_data[62]), .D(n1518), 
        .Y(n2507) );
  scg2d1_hd U56 ( .A(n2236), .B(r_y_data[95]), .C(r_y_data[63]), .D(n1518), 
        .Y(n2482) );
  scg2d1_hd U58 ( .A(n1518), .B(r_x_data[87]), .C(n2415), .D(n2416), .Y(n2702)
         );
  clknd2d1_hd U60 ( .A(w_add_1_Z[23]), .B(N714), .Y(n2417) );
  scg2d1_hd U61 ( .A(n1518), .B(r_x_data[88]), .C(n2418), .D(n2419), .Y(n2703)
         );
  clknd2d1_hd U62 ( .A(w_add_1_Z[24]), .B(N714), .Y(n2420) );
  scg2d1_hd U64 ( .A(n1518), .B(r_x_data[89]), .C(n2421), .D(n2422), .Y(n2704)
         );
  clknd2d1_hd U65 ( .A(w_add_1_Z[25]), .B(N714), .Y(n2423) );
  scg2d1_hd U66 ( .A(n1518), .B(r_x_data[90]), .C(n2424), .D(n2425), .Y(n2705)
         );
  clknd2d1_hd U67 ( .A(w_add_1_Z[26]), .B(N714), .Y(n2426) );
  scg2d1_hd U68 ( .A(n1518), .B(r_x_data[91]), .C(n2427), .D(n2428), .Y(n2706)
         );
  clknd2d1_hd U69 ( .A(w_add_1_Z[27]), .B(N714), .Y(n2429) );
  scg2d1_hd U70 ( .A(n1518), .B(r_x_data[92]), .C(n2430), .D(n2431), .Y(n2707)
         );
  clknd2d1_hd U71 ( .A(w_add_1_Z[28]), .B(N714), .Y(n2432) );
  scg2d1_hd U72 ( .A(r_x_data[85]), .B(n1518), .C(n2711), .D(n2221), .Y(n2700)
         );
  scg2d1_hd U73 ( .A(r_x_data[86]), .B(n1518), .C(n2711), .D(n2222), .Y(n2701)
         );
  scg2d1_hd U74 ( .A(r_x_data[94]), .B(n1518), .C(n2711), .D(n2223), .Y(n2709)
         );
  scg2d1_hd U75 ( .A(r_x_data[84]), .B(n323), .C(n2711), .D(n2220), .Y(n2699)
         );
  ivd4_hd U76 ( .A(n334), .Y(n312) );
  mx2d1_hd U77 ( .D0(r_pstate[0]), .D1(n2468), .S(n2469), .Y(n2257) );
  clknd2d1_hd U78 ( .A(n2259), .B(n2260), .Y(n2468) );
  clknd2d1_hd U79 ( .A(n2), .B(n1508), .Y(n2261) );
  mx2d1_hd U80 ( .D0(o_Y_DATA_VALID), .D1(N1000), .S(N1001), .Y(n2258) );
  scg2d1_hd U81 ( .A(n2236), .B(r_y_data[79]), .C(r_y_data[47]), .D(n323), .Y(
        n2508) );
  scg2d1_hd U82 ( .A(n2236), .B(r_y_data[86]), .C(r_y_data[54]), .D(n323), .Y(
        n2509) );
  scg2d1_hd U83 ( .A(r_x_data[64]), .B(n323), .C(n2711), .D(n2226), .Y(n2679)
         );
  scg2d1_hd U84 ( .A(r_x_data[65]), .B(n323), .C(n2711), .D(n2227), .Y(n2680)
         );
  scg2d1_hd U85 ( .A(r_x_data[66]), .B(n323), .C(n2711), .D(n2228), .Y(n2681)
         );
  scg2d1_hd U86 ( .A(r_x_data[67]), .B(n323), .C(n2711), .D(n2204), .Y(n2682)
         );
  scg2d1_hd U87 ( .A(r_x_data[68]), .B(n323), .C(n2711), .D(n2205), .Y(n2683)
         );
  scg2d1_hd U88 ( .A(r_x_data[69]), .B(n323), .C(n2711), .D(n2229), .Y(n2684)
         );
  scg2d1_hd U89 ( .A(r_x_data[70]), .B(n323), .C(n2711), .D(n2206), .Y(n2685)
         );
  scg2d1_hd U90 ( .A(r_x_data[71]), .B(n323), .C(n2711), .D(n2230), .Y(n2686)
         );
  scg2d1_hd U91 ( .A(r_x_data[73]), .B(n323), .C(n2711), .D(n2231), .Y(n2688)
         );
  scg2d1_hd U92 ( .A(n1516), .B(r_x_data[93]), .C(n2433), .D(n2434), .Y(n2708)
         );
  clknd2d1_hd U93 ( .A(w_add_1_Z[29]), .B(N714), .Y(n2435) );
  scg2d1_hd U94 ( .A(r_x_data[72]), .B(n1516), .C(n2711), .D(n2211), .Y(n2687)
         );
  scg2d1_hd U95 ( .A(r_x_data[74]), .B(n1516), .C(n2711), .D(n2212), .Y(n2689)
         );
  scg2d1_hd U96 ( .A(r_x_data[75]), .B(n1516), .C(n2711), .D(n2232), .Y(n2690)
         );
  scg2d1_hd U97 ( .A(r_x_data[76]), .B(n1516), .C(n2711), .D(n2213), .Y(n2691)
         );
  scg2d1_hd U98 ( .A(r_x_data[77]), .B(n1516), .C(n2711), .D(n2214), .Y(n2692)
         );
  scg2d1_hd U99 ( .A(r_x_data[78]), .B(n1516), .C(n2711), .D(n2215), .Y(n2693)
         );
  scg2d1_hd U100 ( .A(r_x_data[79]), .B(n1516), .C(n2711), .D(n2207), .Y(n2694) );
  scg2d1_hd U101 ( .A(r_x_data[80]), .B(n1516), .C(n2711), .D(n2216), .Y(n2695) );
  scg2d1_hd U103 ( .A(r_x_data[81]), .B(n1516), .C(n2711), .D(n2217), .Y(n2696) );
  scg2d1_hd U104 ( .A(r_x_data[82]), .B(n1516), .C(n2711), .D(n2218), .Y(n2697) );
  scg2d1_hd U105 ( .A(r_x_data[83]), .B(n1516), .C(n2711), .D(n2219), .Y(n2698) );
  clknd2d1_hd U106 ( .A(w_mult_1_Z[18]), .B(n1502), .Y(n2414) );
  nr2d1_hd U107 ( .A(n2233), .B(n327), .Y(n314) );
  mx2d1_hd U108 ( .D0(r_pstate[1]), .D1(n2470), .S(n2471), .Y(n2256) );
  nr2d1_hd U109 ( .A(n2236), .B(n323), .Y(n324) );
  nr2d1_hd U110 ( .A(N715), .B(n1506), .Y(n2196) );
  ivd2_hd U111 ( .A(N715), .Y(n327) );
  ivd1_hd U112 ( .A(n2196), .Y(n2197) );
  ivd1_hd U113 ( .A(n2196), .Y(n2198) );
  ivd1_hd U114 ( .A(n2196), .Y(n2199) );
  ivd2_hd U115 ( .A(n327), .Y(n2711) );
  or2d4_hd U116 ( .A(n1502), .B(n1506), .Y(N1407) );
  scg2d1_hd U117 ( .A(N1407), .B(N1376), .C(r_x_data[159]), .D(n323), .Y(n2333) );
  clknd2d1_hd U118 ( .A(r_x_data[127]), .B(n323), .Y(n2407) );
  ivd6_hd U119 ( .A(n326), .Y(n323) );
  ivd1_hd U120 ( .A(n324), .Y(n2477) );
  ivd1_hd U121 ( .A(n324), .Y(n2476) );
  ivd3_hd U122 ( .A(N723), .Y(n2544) );
  or2d1_hd U123 ( .A(N722), .B(N46), .Y(N723) );
  or2d4_hd U124 ( .A(N715), .B(n1502), .Y(N1408) );
  nid4_hd U125 ( .A(w_rst), .Y(n848) );
  nr2d4_hd U127 ( .A(N719), .B(r_counter[0]), .Y(n1506) );
  nr2d6_hd U129 ( .A(N716), .B(N46), .Y(n1502) );
  ad2d1_hd U130 ( .A(w_add_1_Z[28]), .B(n2237), .Y(n2200) );
  ad2d1_hd U131 ( .A(w_add_1_Z[27]), .B(n2237), .Y(n2201) );
  ad2d1_hd U132 ( .A(w_add_1_Z[24]), .B(n2237), .Y(n2202) );
  ad2d1_hd U133 ( .A(w_add_1_Z[23]), .B(n2237), .Y(n2203) );
  or2d1_hd U134 ( .A(N32), .B(r_pstate[0]), .Y(N37) );
  ivd2_hd U135 ( .A(N37), .Y(n2237) );
  ad2d1_hd U136 ( .A(w_add_1_Z[3]), .B(n2235), .Y(n2204) );
  ad2d1_hd U137 ( .A(w_add_1_Z[4]), .B(n2235), .Y(n2205) );
  ad2d1_hd U138 ( .A(w_add_1_Z[6]), .B(n2235), .Y(n2206) );
  ad2d1_hd U139 ( .A(w_add_1_Z[15]), .B(n2235), .Y(n2207) );
  ad2d1_hd U140 ( .A(w_add_1_Z[29]), .B(n2237), .Y(n2208) );
  ad2d1_hd U141 ( .A(w_add_1_Z[26]), .B(n2237), .Y(n2209) );
  ad2d1_hd U142 ( .A(w_add_1_Z[25]), .B(n2237), .Y(n2210) );
  ivd6_hd U143 ( .A(n2236), .Y(n2233) );
  ad2d1_hd U144 ( .A(w_add_1_Z[8]), .B(n2237), .Y(n2211) );
  ad2d1_hd U145 ( .A(w_add_1_Z[10]), .B(n2237), .Y(n2212) );
  ad2d1_hd U146 ( .A(w_add_1_Z[12]), .B(n2237), .Y(n2213) );
  ad2d1_hd U147 ( .A(w_add_1_Z[13]), .B(n2237), .Y(n2214) );
  ad2d1_hd U148 ( .A(w_add_1_Z[14]), .B(n2237), .Y(n2215) );
  ad2d1_hd U149 ( .A(w_add_1_Z[16]), .B(n2237), .Y(n2216) );
  ad2d1_hd U150 ( .A(w_add_1_Z[17]), .B(n2237), .Y(n2217) );
  ad2d1_hd U151 ( .A(w_add_1_Z[18]), .B(n2237), .Y(n2218) );
  ad2d1_hd U152 ( .A(w_add_1_Z[19]), .B(n2237), .Y(n2219) );
  ad2d1_hd U153 ( .A(w_add_1_Z[20]), .B(n2237), .Y(n2220) );
  ad2d1_hd U154 ( .A(w_add_1_Z[21]), .B(n2237), .Y(n2221) );
  ad2d1_hd U155 ( .A(w_add_1_Z[22]), .B(n2237), .Y(n2222) );
  ad2d1_hd U156 ( .A(w_add_1_Z[30]), .B(n2237), .Y(n2223) );
  clknd2d1_hd U157 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(n2224) );
  or2d1_hd U158 ( .A(n314), .B(n323), .Y(n2225) );
  clknd2d1_hd U159 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(n2) );
  ad2d1_hd U160 ( .A(w_add_1_Z[0]), .B(n2235), .Y(n2226) );
  ad2d1_hd U161 ( .A(w_add_1_Z[1]), .B(n2235), .Y(n2227) );
  ad2d1_hd U162 ( .A(w_add_1_Z[2]), .B(n2235), .Y(n2228) );
  ad2d1_hd U163 ( .A(w_add_1_Z[5]), .B(n2235), .Y(n2229) );
  ad2d1_hd U164 ( .A(w_add_1_Z[7]), .B(n2235), .Y(n2230) );
  ad2d1_hd U165 ( .A(w_add_1_Z[9]), .B(n2235), .Y(n2231) );
  ad2d1_hd U166 ( .A(w_add_1_Z[11]), .B(n2235), .Y(n2232) );
  nid2_hd U167 ( .A(n2237), .Y(n2235) );
  ivd1_hd U168 ( .A(r_pstate[1]), .Y(N32) );
  ivd6_hd U169 ( .A(n2237), .Y(n2234) );
  ivd2_hd U170 ( .A(N37), .Y(n2236) );
  oa211d1_hd U171 ( .A(n1509), .B(N33), .C(r_pstate[1]), .D(N754), .Y(n2260)
         );
  oa211d1_hd U172 ( .A(n1508), .B(N33), .C(n1544), .D(N32), .Y(n2259) );
  scg10d1_hd U173 ( .A(r_pstate[1]), .B(n2261), .C(N754), .D(n2262), .Y(n2469)
         );
  nd2bd1_hd U174 ( .AN(n316), .B(n2263), .Y(n2470) );
  oa211d1_hd U175 ( .A(n1509), .B(N32), .C(r_pstate[0]), .D(n2472), .Y(n2263)
         );
  nd3d1_hd U176 ( .A(r_pstate[0]), .B(n1509), .C(n2264), .Y(n2471) );
  nr2d1_hd U177 ( .A(n316), .B(n2472), .Y(n2264) );
  ivd1_hd U178 ( .A(n1508), .Y(n2472) );
  ivd1_hd U179 ( .A(n2265), .Y(n2511) );
  scg16d1_hd U180 ( .A(n322), .B(n2235), .C(n849), .Y(n2265) );
  oa21d1_hd U181 ( .A(n2233), .B(n2266), .C(n2267), .Y(n2512) );
  ao22d1_hd U182 ( .A(r_x_data[0]), .B(n323), .C(n312), .D(w_mult_2_Z[0]), .Y(
        n2267) );
  ao22d1_hd U183 ( .A(w_mult_1_Z[0]), .B(n2198), .C(n2544), .D(w_add_1_Z[0]), 
        .Y(n2266) );
  oa21d1_hd U184 ( .A(n2234), .B(n2268), .C(n2269), .Y(n2513) );
  ao22d1_hd U186 ( .A(r_x_data[1]), .B(n323), .C(n312), .D(w_mult_2_Z[1]), .Y(
        n2269) );
  ao22d1_hd U187 ( .A(n2197), .B(w_mult_1_Z[1]), .C(n2544), .D(w_add_1_Z[1]), 
        .Y(n2268) );
  oa21d1_hd U188 ( .A(n2234), .B(n2270), .C(n2271), .Y(n2514) );
  ao22d1_hd U189 ( .A(r_x_data[2]), .B(n1518), .C(n312), .D(w_mult_2_Z[2]), 
        .Y(n2271) );
  ao22d1_hd U190 ( .A(n2198), .B(w_mult_1_Z[2]), .C(n2544), .D(w_add_1_Z[2]), 
        .Y(n2270) );
  oa21d1_hd U191 ( .A(n2234), .B(n2272), .C(n2273), .Y(n2515) );
  ao22d1_hd U192 ( .A(r_x_data[3]), .B(n323), .C(n312), .D(w_mult_2_Z[3]), .Y(
        n2273) );
  ao22d1_hd U193 ( .A(n2199), .B(w_mult_1_Z[3]), .C(n2544), .D(w_add_1_Z[3]), 
        .Y(n2272) );
  oa21d1_hd U194 ( .A(n2234), .B(n2274), .C(n2275), .Y(n2516) );
  ao22d1_hd U195 ( .A(r_x_data[4]), .B(n1518), .C(n312), .D(w_mult_2_Z[4]), 
        .Y(n2275) );
  ao22d1_hd U196 ( .A(n2197), .B(w_mult_1_Z[4]), .C(n2544), .D(w_add_1_Z[4]), 
        .Y(n2274) );
  oa21d1_hd U197 ( .A(n2234), .B(n2276), .C(n2277), .Y(n2517) );
  ao22d1_hd U198 ( .A(r_x_data[5]), .B(n1518), .C(n312), .D(w_mult_2_Z[5]), 
        .Y(n2277) );
  ao22d1_hd U199 ( .A(n2198), .B(w_mult_1_Z[5]), .C(n2544), .D(w_add_1_Z[5]), 
        .Y(n2276) );
  oa21d1_hd U200 ( .A(n2234), .B(n2278), .C(n2279), .Y(n2518) );
  ao22d1_hd U201 ( .A(r_x_data[6]), .B(n323), .C(n312), .D(w_mult_2_Z[6]), .Y(
        n2279) );
  ao22d1_hd U202 ( .A(n2199), .B(w_mult_1_Z[6]), .C(n2544), .D(w_add_1_Z[6]), 
        .Y(n2278) );
  oa21d1_hd U203 ( .A(n2234), .B(n2280), .C(n2281), .Y(n2519) );
  ao22d1_hd U204 ( .A(r_x_data[7]), .B(n1518), .C(n312), .D(w_mult_2_Z[7]), 
        .Y(n2281) );
  ao22d1_hd U205 ( .A(n2197), .B(w_mult_1_Z[7]), .C(n2544), .D(w_add_1_Z[7]), 
        .Y(n2280) );
  oa21d1_hd U206 ( .A(n2234), .B(n2282), .C(n2283), .Y(n2520) );
  ao22d1_hd U207 ( .A(r_x_data[8]), .B(n323), .C(n312), .D(w_mult_2_Z[8]), .Y(
        n2283) );
  ao22d1_hd U208 ( .A(n2198), .B(w_mult_1_Z[8]), .C(n2544), .D(w_add_1_Z[8]), 
        .Y(n2282) );
  oa21d1_hd U209 ( .A(n2234), .B(n2284), .C(n2285), .Y(n2521) );
  ao22d1_hd U210 ( .A(r_x_data[9]), .B(n323), .C(n312), .D(w_mult_2_Z[9]), .Y(
        n2285) );
  ao22d1_hd U211 ( .A(n2199), .B(w_mult_1_Z[9]), .C(n2544), .D(w_add_1_Z[9]), 
        .Y(n2284) );
  oa21d1_hd U212 ( .A(n2234), .B(n2286), .C(n2287), .Y(n2522) );
  ao22d1_hd U213 ( .A(r_x_data[10]), .B(n1518), .C(n312), .D(w_mult_2_Z[10]), 
        .Y(n2287) );
  ao22d1_hd U214 ( .A(n2197), .B(w_mult_1_Z[10]), .C(n2544), .D(w_add_1_Z[10]), 
        .Y(n2286) );
  oa21d1_hd U215 ( .A(n2234), .B(n2288), .C(n2289), .Y(n2523) );
  ao22d1_hd U216 ( .A(r_x_data[11]), .B(n1516), .C(n312), .D(w_mult_2_Z[11]), 
        .Y(n2289) );
  ao22d1_hd U217 ( .A(n2198), .B(w_mult_1_Z[11]), .C(n2544), .D(w_add_1_Z[11]), 
        .Y(n2288) );
  oa21d1_hd U218 ( .A(n2234), .B(n2290), .C(n2291), .Y(n2524) );
  ao22d1_hd U219 ( .A(r_x_data[12]), .B(n1516), .C(n312), .D(w_mult_2_Z[12]), 
        .Y(n2291) );
  ao22d1_hd U220 ( .A(n2199), .B(w_mult_1_Z[12]), .C(n2544), .D(w_add_1_Z[12]), 
        .Y(n2290) );
  oa21d1_hd U221 ( .A(n2234), .B(n2292), .C(n2293), .Y(n2525) );
  ao22d1_hd U222 ( .A(r_x_data[13]), .B(n1516), .C(n312), .D(w_mult_2_Z[13]), 
        .Y(n2293) );
  ao22d1_hd U223 ( .A(n2197), .B(w_mult_1_Z[13]), .C(n2544), .D(w_add_1_Z[13]), 
        .Y(n2292) );
  oa21d1_hd U224 ( .A(n2234), .B(n2294), .C(n2295), .Y(n2526) );
  ao22d1_hd U225 ( .A(r_x_data[14]), .B(n1516), .C(n312), .D(w_mult_2_Z[14]), 
        .Y(n2295) );
  ao22d1_hd U227 ( .A(n2198), .B(w_mult_1_Z[14]), .C(n2544), .D(w_add_1_Z[14]), 
        .Y(n2294) );
  oa21d1_hd U228 ( .A(n2234), .B(n2296), .C(n2297), .Y(n2527) );
  ao22d1_hd U229 ( .A(r_x_data[15]), .B(n323), .C(n312), .D(w_mult_2_Z[15]), 
        .Y(n2297) );
  ao22d1_hd U230 ( .A(n2199), .B(w_mult_1_Z[15]), .C(n2544), .D(w_add_1_Z[15]), 
        .Y(n2296) );
  oa21d1_hd U231 ( .A(n2234), .B(n2298), .C(n2299), .Y(n2528) );
  ao22d1_hd U232 ( .A(r_x_data[16]), .B(n323), .C(n312), .D(w_mult_2_Z[16]), 
        .Y(n2299) );
  ao22d1_hd U233 ( .A(n2197), .B(w_mult_1_Z[16]), .C(n2544), .D(w_add_1_Z[16]), 
        .Y(n2298) );
  oa21d1_hd U234 ( .A(n2234), .B(n2300), .C(n2301), .Y(n2529) );
  ao22d1_hd U235 ( .A(r_x_data[17]), .B(n1516), .C(n312), .D(w_mult_2_Z[17]), 
        .Y(n2301) );
  ao22d1_hd U236 ( .A(n2198), .B(w_mult_1_Z[17]), .C(n2544), .D(w_add_1_Z[17]), 
        .Y(n2300) );
  oa21d1_hd U238 ( .A(n2234), .B(n2302), .C(n2303), .Y(n2530) );
  ao22d1_hd U239 ( .A(r_x_data[18]), .B(n1518), .C(n312), .D(w_mult_2_Z[18]), 
        .Y(n2303) );
  ao22d1_hd U240 ( .A(n2199), .B(w_mult_1_Z[18]), .C(n2544), .D(w_add_1_Z[18]), 
        .Y(n2302) );
  oa21d1_hd U241 ( .A(n2234), .B(n2304), .C(n2305), .Y(n2531) );
  ao22d1_hd U242 ( .A(r_x_data[19]), .B(n1518), .C(n312), .D(w_mult_2_Z[19]), 
        .Y(n2305) );
  ao22d1_hd U243 ( .A(n2197), .B(w_mult_1_Z[19]), .C(n2544), .D(w_add_1_Z[19]), 
        .Y(n2304) );
  oa21d1_hd U244 ( .A(n2234), .B(n2306), .C(n2307), .Y(n2532) );
  ao22d1_hd U245 ( .A(r_x_data[20]), .B(n323), .C(n312), .D(w_mult_2_Z[20]), 
        .Y(n2307) );
  ao22d1_hd U246 ( .A(n2198), .B(w_mult_1_Z[20]), .C(n2544), .D(w_add_1_Z[20]), 
        .Y(n2306) );
  oa21d1_hd U247 ( .A(n2234), .B(n2308), .C(n2309), .Y(n2533) );
  ao22d1_hd U248 ( .A(r_x_data[21]), .B(n1518), .C(n312), .D(w_mult_2_Z[21]), 
        .Y(n2309) );
  ao22d1_hd U249 ( .A(n2199), .B(w_mult_1_Z[21]), .C(n2544), .D(w_add_1_Z[21]), 
        .Y(n2308) );
  oa21d1_hd U250 ( .A(n2234), .B(n2310), .C(n2311), .Y(n2534) );
  ao22d1_hd U251 ( .A(r_x_data[22]), .B(n1516), .C(n312), .D(w_mult_2_Z[22]), 
        .Y(n2311) );
  ao22d1_hd U252 ( .A(n2197), .B(w_mult_1_Z[22]), .C(n2544), .D(w_add_1_Z[22]), 
        .Y(n2310) );
  oa21d1_hd U253 ( .A(n2234), .B(n2312), .C(n2313), .Y(n2535) );
  ao22d1_hd U254 ( .A(r_x_data[23]), .B(n1516), .C(n312), .D(w_mult_2_Z[23]), 
        .Y(n2313) );
  ao22d1_hd U255 ( .A(n2198), .B(w_mult_1_Z[23]), .C(n2544), .D(w_add_1_Z[23]), 
        .Y(n2312) );
  oa21d1_hd U256 ( .A(n2234), .B(n2314), .C(n2315), .Y(n2536) );
  ao22d1_hd U257 ( .A(r_x_data[24]), .B(n1516), .C(n312), .D(w_mult_2_Z[24]), 
        .Y(n2315) );
  ao22d1_hd U258 ( .A(n2199), .B(w_mult_1_Z[24]), .C(n2544), .D(w_add_1_Z[24]), 
        .Y(n2314) );
  oa21d1_hd U259 ( .A(n2234), .B(n2316), .C(n2317), .Y(n2537) );
  ao22d1_hd U260 ( .A(r_x_data[25]), .B(n1516), .C(n312), .D(w_mult_2_Z[25]), 
        .Y(n2317) );
  ao22d1_hd U262 ( .A(n2197), .B(w_mult_1_Z[25]), .C(n2544), .D(w_add_1_Z[25]), 
        .Y(n2316) );
  oa21d1_hd U263 ( .A(n2234), .B(n2318), .C(n2319), .Y(n2538) );
  ao22d1_hd U264 ( .A(r_x_data[26]), .B(n1516), .C(n312), .D(w_mult_2_Z[26]), 
        .Y(n2319) );
  ao22d1_hd U266 ( .A(n2198), .B(w_mult_1_Z[26]), .C(n2544), .D(w_add_1_Z[26]), 
        .Y(n2318) );
  oa21d1_hd U267 ( .A(n2234), .B(n2320), .C(n2321), .Y(n2539) );
  ao22d1_hd U269 ( .A(r_x_data[27]), .B(n1516), .C(n312), .D(w_mult_2_Z[27]), 
        .Y(n2321) );
  ao22d1_hd U270 ( .A(n2199), .B(w_mult_1_Z[27]), .C(n2544), .D(w_add_1_Z[27]), 
        .Y(n2320) );
  oa21d1_hd U271 ( .A(n2234), .B(n2322), .C(n2323), .Y(n2540) );
  ao22d1_hd U272 ( .A(r_x_data[28]), .B(n1516), .C(n312), .D(w_mult_2_Z[28]), 
        .Y(n2323) );
  ao22d1_hd U273 ( .A(n2197), .B(w_mult_1_Z[28]), .C(n2544), .D(w_add_1_Z[28]), 
        .Y(n2322) );
  oa21d1_hd U274 ( .A(n2234), .B(n2324), .C(n2325), .Y(n2541) );
  ao22d1_hd U275 ( .A(r_x_data[29]), .B(n1516), .C(n312), .D(w_mult_2_Z[29]), 
        .Y(n2325) );
  ao22d1_hd U276 ( .A(n2198), .B(w_mult_1_Z[29]), .C(n2544), .D(w_add_1_Z[29]), 
        .Y(n2324) );
  oa21d1_hd U277 ( .A(n2234), .B(n2326), .C(n2327), .Y(n2542) );
  ao22d1_hd U278 ( .A(r_x_data[30]), .B(n1516), .C(n312), .D(w_mult_2_Z[30]), 
        .Y(n2327) );
  ao22d1_hd U279 ( .A(n2199), .B(w_mult_1_Z[30]), .C(n2544), .D(w_add_1_Z[30]), 
        .Y(n2326) );
  oa21d1_hd U280 ( .A(n2234), .B(n2328), .C(n2329), .Y(n2543) );
  ao22d1_hd U282 ( .A(r_x_data[31]), .B(n1516), .C(n312), .D(w_mult_2_Z[31]), 
        .Y(n2329) );
  ao22d1_hd U283 ( .A(n2197), .B(w_mult_1_Z[31]), .C(w_add_1_Z[31]), .D(n2544), 
        .Y(n2328) );
  scg5d1_hd U284 ( .A(r_x_data[128]), .B(n323), .C(n2226), .D(N1407), .E(
        w_add_2_Z[0]), .F(n309), .Y(n2545) );
  scg5d1_hd U285 ( .A(N1407), .B(n2227), .C(r_x_data[129]), .D(n323), .E(
        w_add_2_Z[1]), .F(n309), .Y(n2546) );
  scg5d1_hd U286 ( .A(N1407), .B(n2228), .C(r_x_data[130]), .D(n323), .E(
        w_add_2_Z[2]), .F(n309), .Y(n2547) );
  scg5d1_hd U287 ( .A(N1407), .B(n2204), .C(r_x_data[131]), .D(n323), .E(
        w_add_2_Z[3]), .F(n309), .Y(n2548) );
  scg5d1_hd U288 ( .A(N1407), .B(n2205), .C(r_x_data[132]), .D(n323), .E(
        w_add_2_Z[4]), .F(n309), .Y(n2549) );
  scg5d1_hd U289 ( .A(N1407), .B(n2229), .C(r_x_data[133]), .D(n1518), .E(
        w_add_2_Z[5]), .F(n309), .Y(n2550) );
  scg5d1_hd U290 ( .A(N1407), .B(n2206), .C(r_x_data[134]), .D(n323), .E(
        w_add_2_Z[6]), .F(n309), .Y(n2551) );
  scg5d1_hd U291 ( .A(N1407), .B(n2230), .C(r_x_data[135]), .D(n1518), .E(
        w_add_2_Z[7]), .F(n309), .Y(n2552) );
  scg5d1_hd U292 ( .A(N1407), .B(n2211), .C(r_x_data[136]), .D(n323), .E(
        w_add_2_Z[8]), .F(n309), .Y(n2553) );
  scg5d1_hd U294 ( .A(N1407), .B(n2231), .C(r_x_data[137]), .D(n323), .E(
        w_add_2_Z[9]), .F(n309), .Y(n2554) );
  scg5d1_hd U296 ( .A(N1407), .B(n2212), .C(r_x_data[138]), .D(n323), .E(
        w_add_2_Z[10]), .F(n309), .Y(n2555) );
  scg5d1_hd U297 ( .A(N1407), .B(n2232), .C(r_x_data[139]), .D(n1518), .E(
        w_add_2_Z[11]), .F(n309), .Y(n2556) );
  scg5d1_hd U303 ( .A(N1407), .B(n2213), .C(r_x_data[140]), .D(n323), .E(
        w_add_2_Z[12]), .F(n309), .Y(n2557) );
  scg5d1_hd U304 ( .A(N1407), .B(n2214), .C(r_x_data[141]), .D(n1518), .E(
        w_add_2_Z[13]), .F(n309), .Y(n2558) );
  scg5d1_hd U305 ( .A(N1407), .B(n2215), .C(r_x_data[142]), .D(n323), .E(
        w_add_2_Z[14]), .F(n309), .Y(n2559) );
  scg5d1_hd U306 ( .A(N1407), .B(n2207), .C(r_x_data[143]), .D(n1518), .E(
        w_add_2_Z[15]), .F(n309), .Y(n2560) );
  scg5d1_hd U307 ( .A(N1407), .B(n2216), .C(r_x_data[144]), .D(n323), .E(
        w_add_2_Z[16]), .F(n309), .Y(n2561) );
  scg5d1_hd U308 ( .A(N1407), .B(n2217), .C(r_x_data[145]), .D(n1518), .E(
        w_add_2_Z[17]), .F(n309), .Y(n2562) );
  scg5d1_hd U309 ( .A(N1407), .B(n2218), .C(r_x_data[146]), .D(n323), .E(
        w_add_2_Z[18]), .F(n309), .Y(n2563) );
  scg5d1_hd U310 ( .A(N1407), .B(n2219), .C(r_x_data[147]), .D(n323), .E(
        w_add_2_Z[19]), .F(n309), .Y(n2564) );
  scg5d1_hd U313 ( .A(N1407), .B(n2220), .C(r_x_data[148]), .D(n323), .E(
        w_add_2_Z[20]), .F(n309), .Y(n2565) );
  scg5d1_hd U314 ( .A(N1407), .B(n2221), .C(r_x_data[149]), .D(n323), .E(
        w_add_2_Z[21]), .F(n309), .Y(n2566) );
  scg5d1_hd U316 ( .A(N1407), .B(n2222), .C(r_x_data[150]), .D(n323), .E(
        w_add_2_Z[22]), .F(n309), .Y(n2567) );
  scg5d1_hd U317 ( .A(N1407), .B(n2203), .C(r_x_data[151]), .D(n323), .E(
        w_add_2_Z[23]), .F(n309), .Y(n2568) );
  scg5d1_hd U318 ( .A(N1407), .B(n2202), .C(r_x_data[152]), .D(n1516), .E(
        w_add_2_Z[24]), .F(n309), .Y(n2569) );
  scg5d1_hd U319 ( .A(N1407), .B(n2210), .C(r_x_data[153]), .D(n323), .E(
        w_add_2_Z[25]), .F(n309), .Y(n2570) );
  scg5d1_hd U320 ( .A(N1407), .B(n2209), .C(r_x_data[154]), .D(n323), .E(
        w_add_2_Z[26]), .F(n309), .Y(n2571) );
  scg5d1_hd U321 ( .A(N1407), .B(n2201), .C(r_x_data[155]), .D(n323), .E(
        w_add_2_Z[27]), .F(n309), .Y(n2572) );
  scg5d1_hd U322 ( .A(N1407), .B(n2200), .C(r_x_data[156]), .D(n323), .E(
        w_add_2_Z[28]), .F(n309), .Y(n2573) );
  scg5d1_hd U323 ( .A(N1407), .B(n2208), .C(r_x_data[157]), .D(n323), .E(
        w_add_2_Z[29]), .F(n309), .Y(n2574) );
  scg5d1_hd U324 ( .A(N1407), .B(n2223), .C(r_x_data[158]), .D(n323), .E(
        w_add_2_Z[30]), .F(n309), .Y(n2575) );
  scg5d1_hd U325 ( .A(N1407), .B(N1376), .C(r_x_data[159]), .D(n323), .E(
        w_add_2_Z[31]), .F(n309), .Y(n2576) );
  oa22d1_hd U326 ( .A(n2330), .B(n2331), .C(n2332), .D(n846), .Y(n2578) );
  scg16d1_hd U329 ( .A(n846), .B(w_add_Z_STB), .C(n309), .Y(n2331) );
  nr2bd1_hd U330 ( .AN(n2332), .B(w_add_2_Z[31]), .Y(n2330) );
  nr2d1_hd U331 ( .A(n2747), .B(n2333), .Y(n2332) );
  oa22ad1_hd U332 ( .A(n2234), .B(n2334), .C(r_x_data[32]), .D(n323), .Y(n2579) );
  ao22d1_hd U333 ( .A(w_add_2_Z[0]), .B(N1407), .C(w_mult_2_Z[0]), .D(n2335), 
        .Y(n2334) );
  ivd1_hd U334 ( .A(n327), .Y(n2335) );
  oa22ad1_hd U335 ( .A(n2234), .B(n2336), .C(r_x_data[33]), .D(n323), .Y(n2580) );
  ao22d1_hd U336 ( .A(w_add_2_Z[1]), .B(N1407), .C(w_mult_2_Z[1]), .D(n2337), 
        .Y(n2336) );
  ivd1_hd U337 ( .A(n327), .Y(n2337) );
  oa22ad1_hd U338 ( .A(n2234), .B(n2338), .C(r_x_data[34]), .D(n323), .Y(n2581) );
  ao22d1_hd U342 ( .A(w_add_2_Z[2]), .B(N1407), .C(w_mult_2_Z[2]), .D(n2339), 
        .Y(n2338) );
  ivd1_hd U343 ( .A(n327), .Y(n2339) );
  oa22ad1_hd U344 ( .A(n2234), .B(n2340), .C(r_x_data[35]), .D(n323), .Y(n2582) );
  ao22d1_hd U345 ( .A(w_add_2_Z[3]), .B(N1407), .C(w_mult_2_Z[3]), .D(n2341), 
        .Y(n2340) );
  ivd1_hd U346 ( .A(n327), .Y(n2341) );
  oa22ad1_hd U347 ( .A(n2234), .B(n2342), .C(r_x_data[36]), .D(n323), .Y(n2583) );
  ao22d1_hd U348 ( .A(w_add_2_Z[4]), .B(N1407), .C(w_mult_2_Z[4]), .D(n2343), 
        .Y(n2342) );
  ivd1_hd U349 ( .A(n327), .Y(n2343) );
  oa22ad1_hd U350 ( .A(n2234), .B(n2344), .C(r_x_data[37]), .D(n323), .Y(n2584) );
  ao22d1_hd U351 ( .A(w_add_2_Z[5]), .B(N1407), .C(w_mult_2_Z[5]), .D(n2345), 
        .Y(n2344) );
  ivd1_hd U352 ( .A(n327), .Y(n2345) );
  oa22ad1_hd U353 ( .A(n2234), .B(n2346), .C(r_x_data[38]), .D(n323), .Y(n2585) );
  ao22d1_hd U354 ( .A(w_add_2_Z[6]), .B(N1407), .C(w_mult_2_Z[6]), .D(n2347), 
        .Y(n2346) );
  ivd1_hd U355 ( .A(n327), .Y(n2347) );
  oa22ad1_hd U356 ( .A(n2234), .B(n2348), .C(r_x_data[39]), .D(n323), .Y(n2586) );
  ao22d1_hd U357 ( .A(w_add_2_Z[7]), .B(N1407), .C(w_mult_2_Z[7]), .D(n2337), 
        .Y(n2348) );
  oa22ad1_hd U358 ( .A(n2234), .B(n2349), .C(r_x_data[40]), .D(n323), .Y(n2587) );
  ao22d1_hd U359 ( .A(w_add_2_Z[8]), .B(N1407), .C(w_mult_2_Z[8]), .D(n2343), 
        .Y(n2349) );
  oa22ad1_hd U360 ( .A(n2234), .B(n2350), .C(r_x_data[41]), .D(n323), .Y(n2588) );
  ao22d1_hd U361 ( .A(w_add_2_Z[9]), .B(N1407), .C(w_mult_2_Z[9]), .D(n2347), 
        .Y(n2350) );
  oa22ad1_hd U362 ( .A(n2234), .B(n2351), .C(r_x_data[42]), .D(n323), .Y(n2589) );
  ao22d1_hd U363 ( .A(w_add_2_Z[10]), .B(N1407), .C(w_mult_2_Z[10]), .D(n2337), 
        .Y(n2351) );
  oa22ad1_hd U364 ( .A(n2234), .B(n2352), .C(r_x_data[43]), .D(n323), .Y(n2590) );
  ao22d1_hd U365 ( .A(w_add_2_Z[11]), .B(N1407), .C(w_mult_2_Z[11]), .D(n2343), 
        .Y(n2352) );
  oa22ad1_hd U366 ( .A(n2234), .B(n2353), .C(r_x_data[44]), .D(n323), .Y(n2591) );
  ao22d1_hd U367 ( .A(w_add_2_Z[12]), .B(N1407), .C(w_mult_2_Z[12]), .D(n2337), 
        .Y(n2353) );
  oa22ad1_hd U368 ( .A(n2234), .B(n2354), .C(r_x_data[45]), .D(n323), .Y(n2592) );
  ao22d1_hd U369 ( .A(w_add_2_Z[13]), .B(N1407), .C(w_mult_2_Z[13]), .D(n2345), 
        .Y(n2354) );
  oa22ad1_hd U370 ( .A(n2234), .B(n2355), .C(r_x_data[46]), .D(n323), .Y(n2593) );
  ao22d1_hd U371 ( .A(w_add_2_Z[14]), .B(N1407), .C(w_mult_2_Z[14]), .D(n2347), 
        .Y(n2355) );
  oa22ad1_hd U372 ( .A(n2234), .B(n2356), .C(r_x_data[47]), .D(n323), .Y(n2594) );
  ao22d1_hd U373 ( .A(w_add_2_Z[15]), .B(N1407), .C(w_mult_2_Z[15]), .D(n2335), 
        .Y(n2356) );
  oa22ad1_hd U374 ( .A(n2234), .B(n2357), .C(r_x_data[48]), .D(n323), .Y(n2595) );
  ao22d1_hd U375 ( .A(w_add_2_Z[16]), .B(N1407), .C(w_mult_2_Z[16]), .D(n2343), 
        .Y(n2357) );
  oa22ad1_hd U376 ( .A(n2234), .B(n2358), .C(r_x_data[49]), .D(n323), .Y(n2596) );
  ao22d1_hd U377 ( .A(w_add_2_Z[17]), .B(N1407), .C(w_mult_2_Z[17]), .D(n2343), 
        .Y(n2358) );
  oa22ad1_hd U378 ( .A(n2234), .B(n2359), .C(r_x_data[50]), .D(n323), .Y(n2597) );
  ao22d1_hd U379 ( .A(w_add_2_Z[18]), .B(N1407), .C(w_mult_2_Z[18]), .D(n2339), 
        .Y(n2359) );
  oa22ad1_hd U380 ( .A(n2234), .B(n2360), .C(r_x_data[51]), .D(n323), .Y(n2598) );
  ao22d1_hd U381 ( .A(w_add_2_Z[19]), .B(N1407), .C(w_mult_2_Z[19]), .D(n2343), 
        .Y(n2360) );
  oa22ad1_hd U382 ( .A(n2234), .B(n2361), .C(r_x_data[52]), .D(n323), .Y(n2599) );
  ao22d1_hd U383 ( .A(w_add_2_Z[20]), .B(N1407), .C(w_mult_2_Z[20]), .D(n2339), 
        .Y(n2361) );
  oa22ad1_hd U384 ( .A(n2234), .B(n2362), .C(r_x_data[53]), .D(n323), .Y(n2600) );
  ao22d1_hd U385 ( .A(w_add_2_Z[21]), .B(N1407), .C(w_mult_2_Z[21]), .D(n2337), 
        .Y(n2362) );
  oa22ad1_hd U386 ( .A(n2234), .B(n2363), .C(r_x_data[54]), .D(n323), .Y(n2601) );
  ao22d1_hd U387 ( .A(w_add_2_Z[22]), .B(N1407), .C(w_mult_2_Z[22]), .D(n2335), 
        .Y(n2363) );
  oa22ad1_hd U388 ( .A(n2234), .B(n2364), .C(r_x_data[55]), .D(n323), .Y(n2602) );
  ao22d1_hd U389 ( .A(w_add_2_Z[23]), .B(N1407), .C(w_mult_2_Z[23]), .D(n2337), 
        .Y(n2364) );
  oa22ad1_hd U390 ( .A(n2234), .B(n2365), .C(r_x_data[56]), .D(n323), .Y(n2603) );
  ao22d1_hd U391 ( .A(w_add_2_Z[24]), .B(N1407), .C(w_mult_2_Z[24]), .D(n2345), 
        .Y(n2365) );
  oa22ad1_hd U392 ( .A(n2234), .B(n2366), .C(r_x_data[57]), .D(n323), .Y(n2604) );
  ao22d1_hd U393 ( .A(w_add_2_Z[25]), .B(N1407), .C(w_mult_2_Z[25]), .D(n2335), 
        .Y(n2366) );
  oa22ad1_hd U394 ( .A(n2234), .B(n2367), .C(r_x_data[58]), .D(n323), .Y(n2605) );
  ao22d1_hd U395 ( .A(w_add_2_Z[26]), .B(N1407), .C(w_mult_2_Z[26]), .D(n2335), 
        .Y(n2367) );
  oa22ad1_hd U396 ( .A(n2234), .B(n2368), .C(r_x_data[59]), .D(n323), .Y(n2606) );
  ao22d1_hd U397 ( .A(w_add_2_Z[27]), .B(N1407), .C(w_mult_2_Z[27]), .D(n2341), 
        .Y(n2368) );
  oa22ad1_hd U398 ( .A(n2234), .B(n2369), .C(r_x_data[60]), .D(n323), .Y(n2607) );
  ao22d1_hd U399 ( .A(w_add_2_Z[28]), .B(N1407), .C(w_mult_2_Z[28]), .D(n2347), 
        .Y(n2369) );
  oa22ad1_hd U400 ( .A(n2234), .B(n2370), .C(r_x_data[61]), .D(n323), .Y(n2608) );
  ao22d1_hd U401 ( .A(w_add_2_Z[29]), .B(N1407), .C(w_mult_2_Z[29]), .D(n2343), 
        .Y(n2370) );
  oa22ad1_hd U402 ( .A(n2234), .B(n2371), .C(r_x_data[62]), .D(n323), .Y(n2609) );
  ao22d1_hd U403 ( .A(w_add_2_Z[30]), .B(N1407), .C(w_mult_2_Z[30]), .D(n2339), 
        .Y(n2371) );
  oa22ad1_hd U404 ( .A(n2234), .B(n2372), .C(r_x_data[63]), .D(n323), .Y(n2610) );
  ao22d1_hd U405 ( .A(w_add_2_Z[31]), .B(N1407), .C(w_mult_2_Z[31]), .D(n2335), 
        .Y(n2372) );
  oa22ad1_hd U406 ( .A(n2234), .B(n2373), .C(r_x_data[96]), .D(n323), .Y(n2611) );
  ao22d1_hd U407 ( .A(N1408), .B(w_mult_3_Z[0]), .C(w_mult_2_Z[0]), .D(n1506), 
        .Y(n2373) );
  oa22ad1_hd U408 ( .A(n2234), .B(n2374), .C(n323), .D(r_x_data[97]), .Y(n2612) );
  ao22d1_hd U409 ( .A(w_mult_2_Z[1]), .B(n1506), .C(N1408), .D(w_mult_3_Z[1]), 
        .Y(n2374) );
  oa22ad1_hd U410 ( .A(n2234), .B(n2375), .C(n323), .D(r_x_data[98]), .Y(n2613) );
  ao22d1_hd U411 ( .A(w_mult_2_Z[2]), .B(n1506), .C(N1408), .D(w_mult_3_Z[2]), 
        .Y(n2375) );
  oa22ad1_hd U412 ( .A(n2234), .B(n2376), .C(n323), .D(r_x_data[99]), .Y(n2614) );
  ao22d1_hd U413 ( .A(w_mult_2_Z[3]), .B(n1506), .C(N1408), .D(w_mult_3_Z[3]), 
        .Y(n2376) );
  oa22ad1_hd U414 ( .A(n2234), .B(n2377), .C(n323), .D(r_x_data[100]), .Y(
        n2615) );
  ao22d1_hd U415 ( .A(w_mult_2_Z[4]), .B(n1506), .C(N1408), .D(w_mult_3_Z[4]), 
        .Y(n2377) );
  oa22ad1_hd U416 ( .A(n2233), .B(n2378), .C(n323), .D(r_x_data[101]), .Y(
        n2616) );
  ao22d1_hd U417 ( .A(w_mult_2_Z[5]), .B(n1506), .C(N1408), .D(w_mult_3_Z[5]), 
        .Y(n2378) );
  oa22ad1_hd U418 ( .A(n2233), .B(n2379), .C(n323), .D(r_x_data[102]), .Y(
        n2617) );
  ao22d1_hd U419 ( .A(w_mult_2_Z[6]), .B(n1506), .C(N1408), .D(w_mult_3_Z[6]), 
        .Y(n2379) );
  oa22ad1_hd U420 ( .A(n2233), .B(n2380), .C(n323), .D(r_x_data[103]), .Y(
        n2618) );
  ao22d1_hd U421 ( .A(w_mult_2_Z[7]), .B(n1506), .C(N1408), .D(w_mult_3_Z[7]), 
        .Y(n2380) );
  oa22ad1_hd U422 ( .A(n2233), .B(n2381), .C(n323), .D(r_x_data[104]), .Y(
        n2619) );
  ao22d1_hd U423 ( .A(w_mult_2_Z[8]), .B(n1506), .C(N1408), .D(w_mult_3_Z[8]), 
        .Y(n2381) );
  oa22ad1_hd U424 ( .A(n2233), .B(n2382), .C(n323), .D(r_x_data[105]), .Y(
        n2620) );
  ao22d1_hd U425 ( .A(w_mult_2_Z[9]), .B(n1506), .C(N1408), .D(w_mult_3_Z[9]), 
        .Y(n2382) );
  oa22ad1_hd U426 ( .A(n2233), .B(n2383), .C(n323), .D(r_x_data[106]), .Y(
        n2621) );
  ao22d1_hd U427 ( .A(w_mult_2_Z[10]), .B(n1506), .C(N1408), .D(w_mult_3_Z[10]), .Y(n2383) );
  oa22ad1_hd U428 ( .A(n2233), .B(n2384), .C(n323), .D(r_x_data[107]), .Y(
        n2622) );
  ao22d1_hd U429 ( .A(w_mult_2_Z[11]), .B(n1506), .C(N1408), .D(w_mult_3_Z[11]), .Y(n2384) );
  oa22ad1_hd U430 ( .A(n2233), .B(n2385), .C(n323), .D(r_x_data[108]), .Y(
        n2623) );
  ao22d1_hd U431 ( .A(w_mult_2_Z[12]), .B(n1506), .C(N1408), .D(w_mult_3_Z[12]), .Y(n2385) );
  oa22ad1_hd U432 ( .A(n2233), .B(n2386), .C(n323), .D(r_x_data[109]), .Y(
        n2624) );
  ao22d1_hd U433 ( .A(w_mult_2_Z[13]), .B(n1506), .C(N1408), .D(w_mult_3_Z[13]), .Y(n2386) );
  oa22ad1_hd U434 ( .A(n2233), .B(n2387), .C(n1516), .D(r_x_data[110]), .Y(
        n2625) );
  ao22d1_hd U435 ( .A(w_mult_2_Z[14]), .B(n1506), .C(N1408), .D(w_mult_3_Z[14]), .Y(n2387) );
  oa22ad1_hd U436 ( .A(n2233), .B(n2388), .C(n323), .D(r_x_data[111]), .Y(
        n2626) );
  ao22d1_hd U437 ( .A(w_mult_2_Z[15]), .B(n1506), .C(N1408), .D(w_mult_3_Z[15]), .Y(n2388) );
  oa22ad1_hd U438 ( .A(n2233), .B(n2389), .C(n323), .D(r_x_data[112]), .Y(
        n2627) );
  ao22d1_hd U439 ( .A(w_mult_2_Z[16]), .B(n1506), .C(N1408), .D(w_mult_3_Z[16]), .Y(n2389) );
  oa22ad1_hd U440 ( .A(n2233), .B(n2390), .C(n323), .D(r_x_data[113]), .Y(
        n2628) );
  ao22d1_hd U441 ( .A(w_mult_2_Z[17]), .B(n1506), .C(N1408), .D(w_mult_3_Z[17]), .Y(n2390) );
  oa22ad1_hd U442 ( .A(n2233), .B(n2391), .C(n323), .D(r_x_data[114]), .Y(
        n2629) );
  ao22d1_hd U443 ( .A(w_mult_2_Z[18]), .B(n1506), .C(N1408), .D(w_mult_3_Z[18]), .Y(n2391) );
  oa22ad1_hd U444 ( .A(n2233), .B(n2392), .C(n323), .D(r_x_data[115]), .Y(
        n2630) );
  ao22d1_hd U445 ( .A(w_mult_2_Z[19]), .B(n1506), .C(N1408), .D(w_mult_3_Z[19]), .Y(n2392) );
  oa22ad1_hd U446 ( .A(n2233), .B(n2393), .C(n323), .D(r_x_data[116]), .Y(
        n2631) );
  ao22d1_hd U447 ( .A(w_mult_2_Z[20]), .B(n1506), .C(N1408), .D(w_mult_3_Z[20]), .Y(n2393) );
  oa22ad1_hd U448 ( .A(n2233), .B(n2394), .C(n323), .D(r_x_data[117]), .Y(
        n2632) );
  ao22d1_hd U449 ( .A(w_mult_2_Z[21]), .B(n1506), .C(N1408), .D(w_mult_3_Z[21]), .Y(n2394) );
  oa22ad1_hd U450 ( .A(n2233), .B(n2395), .C(n323), .D(r_x_data[118]), .Y(
        n2633) );
  ao22d1_hd U451 ( .A(w_mult_2_Z[22]), .B(n1506), .C(N1408), .D(w_mult_3_Z[22]), .Y(n2395) );
  oa22ad1_hd U452 ( .A(n2233), .B(n2396), .C(n323), .D(r_x_data[119]), .Y(
        n2634) );
  ao22d1_hd U453 ( .A(w_mult_2_Z[23]), .B(n1506), .C(N1408), .D(w_mult_3_Z[23]), .Y(n2396) );
  oa22ad1_hd U454 ( .A(n2233), .B(n2397), .C(n323), .D(r_x_data[120]), .Y(
        n2635) );
  ao22d1_hd U455 ( .A(w_mult_2_Z[24]), .B(n1506), .C(N1408), .D(w_mult_3_Z[24]), .Y(n2397) );
  oa22ad1_hd U456 ( .A(n2233), .B(n2398), .C(n323), .D(r_x_data[121]), .Y(
        n2636) );
  ao22d1_hd U457 ( .A(w_mult_2_Z[25]), .B(n1506), .C(N1408), .D(w_mult_3_Z[25]), .Y(n2398) );
  oa22ad1_hd U458 ( .A(n2233), .B(n2399), .C(n323), .D(r_x_data[122]), .Y(
        n2637) );
  ao22d1_hd U459 ( .A(w_mult_2_Z[26]), .B(n1506), .C(N1408), .D(w_mult_3_Z[26]), .Y(n2399) );
  oa22ad1_hd U460 ( .A(n2233), .B(n2400), .C(n323), .D(r_x_data[123]), .Y(
        n2638) );
  ao22d1_hd U461 ( .A(w_mult_2_Z[27]), .B(n1506), .C(N1408), .D(w_mult_3_Z[27]), .Y(n2400) );
  oa22ad1_hd U462 ( .A(n2233), .B(n2401), .C(n323), .D(r_x_data[124]), .Y(
        n2639) );
  ao22d1_hd U463 ( .A(w_mult_2_Z[28]), .B(n1506), .C(N1408), .D(w_mult_3_Z[28]), .Y(n2401) );
  oa22ad1_hd U464 ( .A(n2233), .B(n2402), .C(n323), .D(r_x_data[125]), .Y(
        n2640) );
  ao22d1_hd U465 ( .A(w_mult_2_Z[29]), .B(n1506), .C(N1408), .D(w_mult_3_Z[29]), .Y(n2402) );
  oa22ad1_hd U466 ( .A(n2233), .B(n2403), .C(n323), .D(r_x_data[126]), .Y(
        n2641) );
  ao22d1_hd U467 ( .A(w_mult_2_Z[30]), .B(n1506), .C(N1408), .D(w_mult_3_Z[30]), .Y(n2403) );
  oa22ad1_hd U468 ( .A(n2233), .B(n2404), .C(n323), .D(r_x_data[127]), .Y(
        n2642) );
  ao22d1_hd U469 ( .A(w_mult_2_Z[31]), .B(n1506), .C(N1408), .D(w_mult_3_Z[31]), .Y(n2404) );
  ad2d1_hd U470 ( .A(n850), .B(n2405), .Y(n2644) );
  oa211d1_hd U471 ( .A(n2233), .B(n2406), .C(n322), .D(n2407), .Y(n2405) );
  ao22d1_hd U472 ( .A(w_mult_2_Z[31]), .B(n1506), .C(N1408), .D(w_mult_3_Z[31]), .Y(n2406) );
  scg14d1_hd U473 ( .A(n312), .B(w_mult_1_Z[0]), .C(n326), .Y(n2645) );
  ad2d1_hd U474 ( .A(n312), .B(w_mult_1_Z[1]), .Y(n2646) );
  oa22d1_hd U475 ( .A(n327), .B(n2233), .C(n2234), .D(n2408), .Y(n2647) );
  nd3d1_hd U476 ( .A(n327), .B(w_mult_1_Z[2]), .C(n1502), .Y(n2408) );
  oa22d1_hd U477 ( .A(n327), .B(n2233), .C(n2234), .D(n2409), .Y(n2649) );
  nd3d1_hd U478 ( .A(n327), .B(w_mult_1_Z[4]), .C(n1502), .Y(n2409) );
  scg14d1_hd U479 ( .A(n312), .B(w_mult_1_Z[5]), .C(n326), .Y(n2650) );
  ad2d1_hd U480 ( .A(n312), .B(w_mult_1_Z[6]), .Y(n2651) );
  ad2d1_hd U481 ( .A(n312), .B(w_mult_1_Z[8]), .Y(n2653) );
  ad2d1_hd U482 ( .A(n312), .B(w_mult_1_Z[9]), .Y(n2654) );
  oa22d1_hd U483 ( .A(n327), .B(n2233), .C(n2234), .D(n2410), .Y(n2655) );
  nd3d1_hd U484 ( .A(n327), .B(w_mult_1_Z[10]), .C(n1502), .Y(n2410) );
  oa22d1_hd U485 ( .A(n327), .B(n2233), .C(n2234), .D(n2411), .Y(n2656) );
  nd3d1_hd U486 ( .A(n327), .B(w_mult_1_Z[11]), .C(n1502), .Y(n2411) );
  ad2d1_hd U487 ( .A(n312), .B(w_mult_1_Z[12]), .Y(n2657) );
  scg14d1_hd U488 ( .A(n312), .B(w_mult_1_Z[13]), .C(n326), .Y(n2658) );
  scg14d1_hd U489 ( .A(n312), .B(w_mult_1_Z[14]), .C(n326), .Y(n2659) );
  oa22d1_hd U490 ( .A(n327), .B(n2233), .C(n2234), .D(n2412), .Y(n2660) );
  nd3d1_hd U491 ( .A(n327), .B(w_mult_1_Z[15]), .C(n1502), .Y(n2412) );
  ad2d1_hd U492 ( .A(n312), .B(w_mult_1_Z[16]), .Y(n2661) );
  oa22d1_hd U493 ( .A(n327), .B(n2233), .C(n2234), .D(n2413), .Y(n2662) );
  nd3d1_hd U494 ( .A(n327), .B(w_mult_1_Z[17]), .C(n1502), .Y(n2413) );
  ao21d1_hd U495 ( .A(n2414), .B(n327), .C(n2234), .Y(n2663) );
  scg14d1_hd U496 ( .A(n312), .B(w_mult_1_Z[19]), .C(n326), .Y(n2664) );
  ad2d1_hd U497 ( .A(n312), .B(w_mult_1_Z[20]), .Y(n2665) );
  scg14d1_hd U498 ( .A(n312), .B(w_mult_1_Z[23]), .C(n326), .Y(n2668) );
  scg6d1_hd U499 ( .A(w_mult_1_Z[29]), .B(n2675), .C(n2676), .Y(n2674) );
  scg6d1_hd U500 ( .A(n1502), .B(n2235), .C(n2676), .Y(n2675) );
  scg6d1_hd U501 ( .A(n2711), .B(n2235), .C(n323), .Y(n2676) );
  ad2d1_hd U502 ( .A(n312), .B(w_mult_1_Z[30]), .Y(n2677) );
  ad2d1_hd U503 ( .A(n312), .B(w_mult_1_Z[31]), .Y(n2678) );
  nd2bd1_hd U504 ( .AN(N46), .B(N716), .Y(n2416) );
  ao21d1_hd U505 ( .A(n2417), .B(N46), .C(n2234), .Y(n2415) );
  nd2bd1_hd U506 ( .AN(N46), .B(N716), .Y(n2419) );
  ao21d1_hd U507 ( .A(n2420), .B(N46), .C(n2234), .Y(n2418) );
  nd2bd1_hd U508 ( .AN(N46), .B(N716), .Y(n2422) );
  ao21d1_hd U509 ( .A(n2423), .B(N46), .C(n2234), .Y(n2421) );
  nd2bd1_hd U510 ( .AN(N46), .B(N716), .Y(n2425) );
  ao21d1_hd U511 ( .A(n2426), .B(N46), .C(n2234), .Y(n2424) );
  nd2bd1_hd U512 ( .AN(N46), .B(N716), .Y(n2428) );
  ao21d1_hd U513 ( .A(n2429), .B(N46), .C(n2234), .Y(n2427) );
  nd2bd1_hd U514 ( .AN(N46), .B(N716), .Y(n2431) );
  ao21d1_hd U515 ( .A(n2432), .B(N46), .C(n2234), .Y(n2430) );
  nd2bd1_hd U516 ( .AN(N46), .B(N716), .Y(n2434) );
  ao21d1_hd U517 ( .A(n2435), .B(N46), .C(n2234), .Y(n2433) );
  oa22ad1_hd U518 ( .A(n328), .B(n327), .C(r_x_data[95]), .D(n1518), .Y(n2710)
         );
  nd2bd1_hd U519 ( .AN(n312), .B(n326), .Y(n2712) );
  oa22ad1_hd U520 ( .A(n2233), .B(n2436), .C(r_y_data[0]), .D(n323), .Y(n2713)
         );
  ao22d1_hd U521 ( .A(n1502), .B(r_y_data[96]), .C(w_add_2_Z[0]), .D(n2337), 
        .Y(n2436) );
  oa22ad1_hd U522 ( .A(n2233), .B(n2437), .C(r_y_data[1]), .D(n323), .Y(n2714)
         );
  ao22d1_hd U523 ( .A(n1502), .B(r_y_data[97]), .C(w_add_2_Z[1]), .D(n2345), 
        .Y(n2437) );
  oa22ad1_hd U524 ( .A(n2233), .B(n2438), .C(r_y_data[2]), .D(n323), .Y(n2715)
         );
  ao22d1_hd U525 ( .A(n1502), .B(r_y_data[98]), .C(w_add_2_Z[2]), .D(n2345), 
        .Y(n2438) );
  oa22ad1_hd U526 ( .A(n2233), .B(n2439), .C(r_y_data[3]), .D(n1518), .Y(n2716) );
  ao22d1_hd U527 ( .A(n1502), .B(r_y_data[99]), .C(w_add_2_Z[3]), .D(n2339), 
        .Y(n2439) );
  oa22ad1_hd U528 ( .A(n2233), .B(n2440), .C(r_y_data[4]), .D(n323), .Y(n2717)
         );
  ao22d1_hd U529 ( .A(n1502), .B(r_y_data[100]), .C(w_add_2_Z[4]), .D(n2347), 
        .Y(n2440) );
  oa22ad1_hd U530 ( .A(n2233), .B(n2441), .C(r_y_data[5]), .D(n323), .Y(n2718)
         );
  ao22d1_hd U531 ( .A(n1502), .B(r_y_data[101]), .C(w_add_2_Z[5]), .D(n2335), 
        .Y(n2441) );
  oa22ad1_hd U532 ( .A(n2233), .B(n2442), .C(r_y_data[6]), .D(n323), .Y(n2719)
         );
  ao22d1_hd U533 ( .A(n1502), .B(r_y_data[102]), .C(w_add_2_Z[6]), .D(n2347), 
        .Y(n2442) );
  oa22ad1_hd U534 ( .A(n2233), .B(n2443), .C(r_y_data[7]), .D(n1518), .Y(n2720) );
  ao22d1_hd U535 ( .A(n1502), .B(r_y_data[103]), .C(w_add_2_Z[7]), .D(n2339), 
        .Y(n2443) );
  oa22ad1_hd U536 ( .A(n2233), .B(n2444), .C(r_y_data[8]), .D(n1518), .Y(n2721) );
  ao22d1_hd U537 ( .A(n1502), .B(r_y_data[104]), .C(w_add_2_Z[8]), .D(n2341), 
        .Y(n2444) );
  oa22ad1_hd U538 ( .A(n2233), .B(n2445), .C(r_y_data[9]), .D(n323), .Y(n2722)
         );
  ao22d1_hd U539 ( .A(n1502), .B(r_y_data[105]), .C(w_add_2_Z[9]), .D(n2345), 
        .Y(n2445) );
  oa22ad1_hd U540 ( .A(n2233), .B(n2446), .C(r_y_data[10]), .D(n323), .Y(n2723) );
  ao22d1_hd U541 ( .A(n1502), .B(r_y_data[106]), .C(w_add_2_Z[10]), .D(n2347), 
        .Y(n2446) );
  oa22ad1_hd U542 ( .A(n2233), .B(n2447), .C(r_y_data[11]), .D(n1516), .Y(
        n2724) );
  ao22d1_hd U543 ( .A(n1502), .B(r_y_data[107]), .C(w_add_2_Z[11]), .D(n2335), 
        .Y(n2447) );
  oa22ad1_hd U544 ( .A(n2233), .B(n2448), .C(r_y_data[12]), .D(n323), .Y(n2725) );
  ao22d1_hd U545 ( .A(n1502), .B(r_y_data[108]), .C(w_add_2_Z[12]), .D(n2335), 
        .Y(n2448) );
  oa22ad1_hd U546 ( .A(n2233), .B(n2449), .C(r_y_data[13]), .D(n1518), .Y(
        n2726) );
  ao22d1_hd U547 ( .A(n1502), .B(r_y_data[109]), .C(w_add_2_Z[13]), .D(n2345), 
        .Y(n2449) );
  oa22ad1_hd U548 ( .A(n2233), .B(n2450), .C(r_y_data[14]), .D(n323), .Y(n2727) );
  ao22d1_hd U549 ( .A(n1502), .B(r_y_data[110]), .C(w_add_2_Z[14]), .D(n2341), 
        .Y(n2450) );
  oa22ad1_hd U550 ( .A(n2233), .B(n2451), .C(r_y_data[15]), .D(n323), .Y(n2728) );
  ao22d1_hd U551 ( .A(n1502), .B(r_y_data[111]), .C(w_add_2_Z[15]), .D(n2337), 
        .Y(n2451) );
  oa22ad1_hd U552 ( .A(n2233), .B(n2452), .C(r_y_data[16]), .D(n1518), .Y(
        n2729) );
  ao22d1_hd U553 ( .A(n1502), .B(r_y_data[112]), .C(w_add_2_Z[16]), .D(n2335), 
        .Y(n2452) );
  oa22ad1_hd U554 ( .A(n2233), .B(n2453), .C(r_y_data[17]), .D(n1518), .Y(
        n2730) );
  ao22d1_hd U555 ( .A(n1502), .B(r_y_data[113]), .C(w_add_2_Z[17]), .D(n2339), 
        .Y(n2453) );
  oa22ad1_hd U556 ( .A(n2233), .B(n2454), .C(r_y_data[18]), .D(n323), .Y(n2731) );
  ao22d1_hd U557 ( .A(n1502), .B(r_y_data[114]), .C(w_add_2_Z[18]), .D(n2343), 
        .Y(n2454) );
  oa22ad1_hd U558 ( .A(n2233), .B(n2455), .C(r_y_data[19]), .D(n1518), .Y(
        n2732) );
  ao22d1_hd U559 ( .A(n1502), .B(r_y_data[115]), .C(w_add_2_Z[19]), .D(n2347), 
        .Y(n2455) );
  oa22ad1_hd U560 ( .A(n2233), .B(n2456), .C(r_y_data[20]), .D(n323), .Y(n2733) );
  ao22d1_hd U561 ( .A(n1502), .B(r_y_data[116]), .C(w_add_2_Z[20]), .D(n2339), 
        .Y(n2456) );
  oa22ad1_hd U562 ( .A(n2233), .B(n2457), .C(r_y_data[21]), .D(n1518), .Y(
        n2734) );
  ao22d1_hd U563 ( .A(n1502), .B(r_y_data[117]), .C(w_add_2_Z[21]), .D(n2341), 
        .Y(n2457) );
  oa22ad1_hd U564 ( .A(n2233), .B(n2458), .C(r_y_data[22]), .D(n323), .Y(n2735) );
  ao22d1_hd U565 ( .A(n1502), .B(r_y_data[118]), .C(w_add_2_Z[22]), .D(n2341), 
        .Y(n2458) );
  oa22ad1_hd U566 ( .A(n2233), .B(n2459), .C(r_y_data[23]), .D(n1518), .Y(
        n2736) );
  ao22d1_hd U567 ( .A(n1502), .B(r_y_data[119]), .C(w_add_2_Z[23]), .D(n2345), 
        .Y(n2459) );
  oa22ad1_hd U568 ( .A(n2233), .B(n2460), .C(r_y_data[24]), .D(n1518), .Y(
        n2737) );
  ao22d1_hd U569 ( .A(n1502), .B(r_y_data[120]), .C(w_add_2_Z[24]), .D(n2337), 
        .Y(n2460) );
  oa22ad1_hd U570 ( .A(n2233), .B(n2461), .C(r_y_data[25]), .D(n323), .Y(n2738) );
  ao22d1_hd U571 ( .A(n1502), .B(r_y_data[121]), .C(w_add_2_Z[25]), .D(n2341), 
        .Y(n2461) );
  oa22ad1_hd U572 ( .A(n2233), .B(n2462), .C(r_y_data[26]), .D(n1518), .Y(
        n2739) );
  ao22d1_hd U573 ( .A(n1502), .B(r_y_data[122]), .C(w_add_2_Z[26]), .D(n2341), 
        .Y(n2462) );
  oa22ad1_hd U574 ( .A(n2233), .B(n2463), .C(r_y_data[27]), .D(n1518), .Y(
        n2740) );
  ao22d1_hd U575 ( .A(n1502), .B(r_y_data[123]), .C(w_add_2_Z[27]), .D(n2345), 
        .Y(n2463) );
  oa22ad1_hd U576 ( .A(n2233), .B(n2464), .C(r_y_data[28]), .D(n1518), .Y(
        n2741) );
  ao22d1_hd U577 ( .A(n1502), .B(r_y_data[124]), .C(w_add_2_Z[28]), .D(n2339), 
        .Y(n2464) );
  oa22ad1_hd U578 ( .A(n2233), .B(n2465), .C(r_y_data[29]), .D(n1518), .Y(
        n2742) );
  ao22d1_hd U579 ( .A(n1502), .B(r_y_data[125]), .C(w_add_2_Z[29]), .D(n2343), 
        .Y(n2465) );
  oa22ad1_hd U580 ( .A(n2233), .B(n2466), .C(r_y_data[30]), .D(n1518), .Y(
        n2743) );
  ao22d1_hd U581 ( .A(n1502), .B(r_y_data[126]), .C(w_add_2_Z[30]), .D(n2347), 
        .Y(n2466) );
  oa22ad1_hd U582 ( .A(n2233), .B(n2467), .C(r_y_data[31]), .D(n1518), .Y(
        n2744) );
  ao22d1_hd U583 ( .A(n1502), .B(r_y_data[127]), .C(w_add_2_Z[31]), .D(n2341), 
        .Y(n2467) );
  scg9d1_hd U584 ( .A(n2235), .B(n2747), .C(n851), .Y(n2746) );
  ivd1_hd U585 ( .A(n322), .Y(n2747) );
  ad2d1_hd U586 ( .A(n1544), .B(i_X_DATA[5]), .Y(n2748) );
  ad2d1_hd U587 ( .A(n1544), .B(i_X_DATA[6]), .Y(n2749) );
  ad2d1_hd U588 ( .A(n1544), .B(i_X_DATA[7]), .Y(n2750) );
  ad2d1_hd U589 ( .A(n1544), .B(i_X_DATA[8]), .Y(n2751) );
  ad2d1_hd U590 ( .A(n1544), .B(i_X_DATA[9]), .Y(n2752) );
  ad2d1_hd U591 ( .A(n1544), .B(i_X_DATA[10]), .Y(n2753) );
  ad2d1_hd U592 ( .A(n1544), .B(i_X_DATA[11]), .Y(n2754) );
  ad2d1_hd U593 ( .A(n1543), .B(i_X_DATA[12]), .Y(n2755) );
  ad2d1_hd U594 ( .A(n1543), .B(i_X_DATA[13]), .Y(n2756) );
  ad2d1_hd U595 ( .A(n1543), .B(i_X_DATA[14]), .Y(n2757) );
  ad2d1_hd U596 ( .A(n1543), .B(i_X_DATA[15]), .Y(n2758) );
  ad2d1_hd U597 ( .A(n1543), .B(i_X_DATA[16]), .Y(n2759) );
  ad2d1_hd U598 ( .A(n1543), .B(i_X_DATA[17]), .Y(n2760) );
  ad2d1_hd U599 ( .A(n1544), .B(r_x_data[5]), .Y(n2761) );
  ad2d1_hd U600 ( .A(n1544), .B(r_x_data[6]), .Y(n2762) );
  ad2d1_hd U601 ( .A(n1544), .B(r_x_data[7]), .Y(n2763) );
  ad2d1_hd U602 ( .A(n1544), .B(r_x_data[8]), .Y(n2764) );
  ad2d1_hd U603 ( .A(n1544), .B(r_x_data[9]), .Y(n2765) );
  ad2d1_hd U604 ( .A(n1544), .B(r_x_data[10]), .Y(n2766) );
  ad2d1_hd U605 ( .A(n1544), .B(r_x_data[11]), .Y(n2767) );
  ad2d1_hd U606 ( .A(n1543), .B(r_x_data[12]), .Y(n2768) );
  ad2d1_hd U607 ( .A(n1543), .B(r_x_data[13]), .Y(n2769) );
  ad2d1_hd U608 ( .A(n1543), .B(r_x_data[14]), .Y(n2770) );
  ad2d1_hd U609 ( .A(n1543), .B(r_x_data[15]), .Y(n2771) );
  ad2d1_hd U610 ( .A(n1543), .B(r_x_data[16]), .Y(n2772) );
  ad2d1_hd U611 ( .A(n1543), .B(r_x_data[17]), .Y(n2773) );
  ad2d1_hd U612 ( .A(n1543), .B(r_x_data[18]), .Y(n2774) );
  ad2d1_hd U613 ( .A(n1544), .B(r_x_data[38]), .Y(n2775) );
  ad2d1_hd U614 ( .A(n1544), .B(r_x_data[39]), .Y(n2776) );
  ad2d1_hd U615 ( .A(n1544), .B(r_x_data[40]), .Y(n2777) );
  ad2d1_hd U616 ( .A(n1544), .B(r_x_data[41]), .Y(n2778) );
  ad2d1_hd U617 ( .A(n1544), .B(r_x_data[42]), .Y(n2779) );
  ad2d1_hd U618 ( .A(n1544), .B(r_x_data[43]), .Y(n2780) );
  ad2d1_hd U619 ( .A(n1543), .B(r_x_data[44]), .Y(n2781) );
  ad2d1_hd U620 ( .A(n1543), .B(r_x_data[45]), .Y(n2782) );
  ad2d1_hd U621 ( .A(n1543), .B(r_x_data[46]), .Y(n2783) );
  ad2d1_hd U622 ( .A(n1543), .B(r_x_data[47]), .Y(n2784) );
  ad2d1_hd U623 ( .A(n1543), .B(r_x_data[48]), .Y(n2785) );
  ad2d1_hd U624 ( .A(n1543), .B(r_x_data[49]), .Y(n2786) );
  ad2d1_hd U625 ( .A(n1543), .B(r_x_data[50]), .Y(n2787) );
  ad2d1_hd U626 ( .A(n1544), .B(r_x_data[70]), .Y(n2788) );
  ad2d1_hd U627 ( .A(n1544), .B(r_x_data[71]), .Y(n2789) );
  ad2d1_hd U628 ( .A(n1544), .B(r_x_data[72]), .Y(n2790) );
  ad2d1_hd U629 ( .A(n1544), .B(r_x_data[73]), .Y(n2791) );
  ad2d1_hd U630 ( .A(n1544), .B(r_x_data[74]), .Y(n2792) );
  ad2d1_hd U631 ( .A(n1544), .B(r_x_data[75]), .Y(n2793) );
  ad2d1_hd U632 ( .A(n1543), .B(r_x_data[76]), .Y(n2794) );
  ad2d1_hd U633 ( .A(n1543), .B(r_x_data[77]), .Y(n2795) );
  ad2d1_hd U634 ( .A(n1543), .B(r_x_data[78]), .Y(n2796) );
  ad2d1_hd U635 ( .A(n1543), .B(r_x_data[79]), .Y(n2797) );
  ad2d1_hd U636 ( .A(n1543), .B(r_x_data[80]), .Y(n2798) );
  ad2d1_hd U637 ( .A(n1543), .B(r_x_data[81]), .Y(n2799) );
  ad2d1_hd U638 ( .A(n1543), .B(r_x_data[82]), .Y(n2800) );
  ad2d1_hd U639 ( .A(n1544), .B(r_x_data[102]), .Y(n2801) );
  ad2d1_hd U640 ( .A(n1544), .B(r_x_data[103]), .Y(n2802) );
  ad2d1_hd U641 ( .A(n1544), .B(r_x_data[104]), .Y(n2803) );
  ad2d1_hd U642 ( .A(n1544), .B(r_x_data[105]), .Y(n2804) );
  ad2d1_hd U643 ( .A(n1544), .B(r_x_data[106]), .Y(n2805) );
  ad2d1_hd U644 ( .A(n1544), .B(r_x_data[107]), .Y(n2806) );
  ad2d1_hd U645 ( .A(n1544), .B(r_x_data[108]), .Y(n2807) );
  ad2d1_hd U646 ( .A(n1543), .B(r_x_data[109]), .Y(n2808) );
  ad2d1_hd U647 ( .A(n1543), .B(r_x_data[110]), .Y(n2809) );
  ad2d1_hd U648 ( .A(n1543), .B(r_x_data[111]), .Y(n2810) );
  ad2d1_hd U649 ( .A(n1543), .B(r_x_data[112]), .Y(n2811) );
  ad2d1_hd U650 ( .A(n1543), .B(r_x_data[113]), .Y(n2812) );
  ad2d1_hd U651 ( .A(n1543), .B(r_x_data[114]), .Y(n2813) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_hpf_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_hpf_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_hpf_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_iir_hpf_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module iir_hpf ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   w_rstn, w_rst, r_add_AB_STB, w_add_AB_ACK, w_add_Z_STB, r_add_Z_ACK,
         r_mult_AB_STB, w_mult_AB_ACK, w_mult_Z_STB, r_mult_Z_ACK, N25, N26,
         N27, N28, N37, N38, N39, N48, N49, N114, N311, N317, N319, N320, N322,
         N371, N374, N376, N511, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N546, N548, N550, N552, N554, N556, N557, N558,
         N559, N562, N563, N564, alt24_n18, alt24_n19, alt24_n58, alt24_n109,
         n100, n101, n102, n103, n104, n106, n107, n108, n109, n111, n112,
         n113, n115, n116, n119, n120, n121, n122, n123, n124, n126, n280,
         n535, n536, n537, n538, n539, n540, n541, n543, n544, n545, n546,
         n547, n554, n287, n294, n305, n306, n307, n308, n318, n378, n379,
         n392, n436, n438, n469, n470, n472, n491, n530, n580, n581, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n931;
  wire   [31:0] r_add_A;
  wire   [31:0] r_add_B;
  wire   [31:0] w_add_Z;
  wire   [29:0] r_mult_A;
  wire   [31:0] r_mult_B;
  wire   [31:0] w_mult_Z;
  wire   [63:0] r_x_data;
  wire   [31:0] r_y_data;
  wire   [1:0] r_pstate;
  wire   [1:0] r_counter;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  float_adder add ( .i_A(r_add_A), .i_B(r_add_B), .i_AB_STB(r_add_AB_STB), 
        .o_AB_ACK(w_add_AB_ACK), .o_Z(w_add_Z), .o_Z_STB(w_add_Z_STB), 
        .i_Z_ACK(r_add_Z_ACK), .i_CLK(i_CLK), .i_RST(w_rst) );
  float_multiplier mult ( .i_A({1'b0, 1'b0, r_mult_A[29:24], 1'b0, 
        r_mult_A[22:21], 1'b0, 1'b0, 1'b0, r_mult_A[17:16], 1'b0, 
        r_mult_A[14:13], 1'b0, r_mult_A[11], 1'b0, r_mult_A[9:5], 1'b0, 1'b0, 
        1'b0, r_mult_A[1:0]}), .i_B(r_mult_B), .i_AB_STB(r_mult_AB_STB), 
        .o_AB_ACK(w_mult_AB_ACK), .o_Z(w_mult_Z), .o_Z_STB(w_mult_Z_STB), 
        .i_Z_ACK(r_mult_Z_ACK), .i_CLK(i_CLK), .i_RST(n806) );
  or2d1_hd U116 ( .A(n102), .B(N556), .Y(N557) );
  nr2d1_hd U120 ( .A(n805), .B(n106), .Y(n102) );
  ao211d1_hd U122 ( .A(n807), .B(N564), .C(n109), .D(N371), .Y(n108) );
  nr2d1_hd U123 ( .A(n539), .B(N28), .Y(n109) );
  ao22d1_hd U124 ( .A(n111), .B(N320), .C(N322), .D(n112), .Y(n107) );
  ao22d1_hd U130 ( .A(N311), .B(N317), .C(n538), .D(w_add_Z_STB), .Y(n116) );
  scg22d1_hd U135 ( .A(n104), .B(N48), .C(n539), .D(n805), .Y(N548) );
  ivd1_hd U141 ( .A(n100), .Y(n120) );
  nr2d1_hd U143 ( .A(N320), .B(n122), .Y(n103) );
  nr2bd1_hd U144 ( .AN(N49), .B(N28), .Y(N546) );
  nr2bd1_hd U178 ( .AN(N114), .B(N28), .Y(N511) );
  scg12d1_hd U297 ( .A(n104), .B(N39), .C(n539), .Y(n119) );
  nr2bd1_hd U300 ( .AN(N319), .B(n126), .Y(N376) );
  nr2d1_hd U301 ( .A(n126), .B(r_counter[0]), .Y(N374) );
  nr2d1_hd U302 ( .A(n111), .B(n112), .Y(n126) );
  ad2d1_hd U303 ( .A(n807), .B(n540), .Y(n112) );
  ad2d1_hd U306 ( .A(alt24_n19), .B(n545), .Y(N371) );
  ivd1_hd U463 ( .A(r_counter[0]), .Y(N38) );
  clknd2d1_hd U465 ( .A(n807), .B(N311), .Y(n122) );
  ad2d1_hd U466 ( .A(N37), .B(N38), .Y(N311) );
  ad2d1_hd U467 ( .A(w_add_Z_STB), .B(w_mult_Z_STB), .Y(N317) );
  clknd2d1_hd U468 ( .A(w_mult_Z_STB), .B(n540), .Y(n106) );
  or2d1_hd U469 ( .A(n544), .B(N39), .Y(alt24_n58) );
  ad2d2_hd U472 ( .A(n807), .B(n538), .Y(n121) );
  ivd1_hd U474 ( .A(alt24_n19), .Y(alt24_n18) );
  ad2d1_hd U475 ( .A(r_pstate[1]), .B(r_pstate[0]), .Y(alt24_n19) );
  clknd2d1_hd U476 ( .A(n121), .B(w_add_Z_STB), .Y(n100) );
  nr2d1_hd U477 ( .A(N37), .B(r_counter[0]), .Y(n541) );
  ad2d1_hd U478 ( .A(N37), .B(N38), .Y(N39) );
  nr2d1_hd U479 ( .A(r_counter[1]), .B(N38), .Y(n544) );
  or2d1_hd U480 ( .A(r_pstate[1]), .B(N26), .Y(N28) );
  or3d1_hd U481 ( .A(N39), .B(n544), .C(n541), .Y(N48) );
  or2d1_hd U482 ( .A(n540), .B(N311), .Y(alt24_n109) );
  ivd2_hd U483 ( .A(n122), .Y(n111) );
  clknd2d1_hd U484 ( .A(w_mult_AB_ACK), .B(w_add_AB_ACK), .Y(n539) );
  ivd1_hd U485 ( .A(N28), .Y(n104) );
  clknd2d1_hd U486 ( .A(n807), .B(n554), .Y(n115) );
  clknd2d1_hd U487 ( .A(n116), .B(n106), .Y(n554) );
  clknd2d1_hd U488 ( .A(n113), .B(n115), .Y(N552) );
  ad2d1_hd U489 ( .A(N25), .B(N26), .Y(N27) );
  scg2d1_hd U704 ( .A(w_mult_Z[0]), .B(n111), .C(w_add_Z[0]), .D(n121), .Y(
        N513) );
  scg2d1_hd U706 ( .A(w_mult_Z[1]), .B(n111), .C(w_add_Z[1]), .D(n121), .Y(
        N514) );
  scg2d1_hd U708 ( .A(w_mult_Z[2]), .B(n111), .C(w_add_Z[2]), .D(n121), .Y(
        N515) );
  scg2d1_hd U710 ( .A(w_mult_Z[3]), .B(n111), .C(w_add_Z[3]), .D(n121), .Y(
        N516) );
  scg2d1_hd U712 ( .A(w_mult_Z[4]), .B(n111), .C(w_add_Z[4]), .D(n121), .Y(
        N517) );
  scg2d1_hd U714 ( .A(w_mult_Z[5]), .B(n111), .C(w_add_Z[5]), .D(n121), .Y(
        N518) );
  scg2d1_hd U716 ( .A(w_mult_Z[6]), .B(n111), .C(w_add_Z[6]), .D(n121), .Y(
        N519) );
  scg2d1_hd U718 ( .A(w_mult_Z[7]), .B(n111), .C(w_add_Z[7]), .D(n121), .Y(
        N520) );
  scg2d1_hd U720 ( .A(w_mult_Z[8]), .B(n111), .C(w_add_Z[8]), .D(n121), .Y(
        N521) );
  scg2d1_hd U722 ( .A(w_mult_Z[9]), .B(n111), .C(w_add_Z[9]), .D(n121), .Y(
        N522) );
  scg2d1_hd U724 ( .A(w_mult_Z[10]), .B(n111), .C(w_add_Z[10]), .D(n121), .Y(
        N523) );
  scg2d1_hd U726 ( .A(w_mult_Z[11]), .B(n111), .C(w_add_Z[11]), .D(n121), .Y(
        N524) );
  scg2d1_hd U728 ( .A(w_mult_Z[12]), .B(n111), .C(w_add_Z[12]), .D(n121), .Y(
        N525) );
  scg2d1_hd U730 ( .A(w_mult_Z[13]), .B(n111), .C(w_add_Z[13]), .D(n121), .Y(
        N526) );
  scg2d1_hd U732 ( .A(w_mult_Z[14]), .B(n111), .C(w_add_Z[14]), .D(n121), .Y(
        N527) );
  scg2d1_hd U734 ( .A(w_mult_Z[15]), .B(n111), .C(w_add_Z[15]), .D(n121), .Y(
        N528) );
  scg2d1_hd U736 ( .A(w_mult_Z[16]), .B(n111), .C(w_add_Z[16]), .D(n121), .Y(
        N529) );
  scg2d1_hd U738 ( .A(w_mult_Z[17]), .B(n111), .C(w_add_Z[17]), .D(n121), .Y(
        N530) );
  scg2d1_hd U740 ( .A(w_mult_Z[18]), .B(n111), .C(w_add_Z[18]), .D(n121), .Y(
        N531) );
  scg2d1_hd U742 ( .A(w_mult_Z[19]), .B(n111), .C(w_add_Z[19]), .D(n121), .Y(
        N532) );
  scg2d1_hd U744 ( .A(w_mult_Z[20]), .B(n111), .C(w_add_Z[20]), .D(n121), .Y(
        N533) );
  scg2d1_hd U746 ( .A(w_mult_Z[21]), .B(n111), .C(w_add_Z[21]), .D(n121), .Y(
        N534) );
  scg2d1_hd U748 ( .A(w_mult_Z[22]), .B(n111), .C(w_add_Z[22]), .D(n121), .Y(
        N535) );
  scg2d1_hd U750 ( .A(w_mult_Z[23]), .B(n111), .C(w_add_Z[23]), .D(n121), .Y(
        N536) );
  scg2d1_hd U752 ( .A(w_mult_Z[24]), .B(n111), .C(w_add_Z[24]), .D(n121), .Y(
        N537) );
  scg2d1_hd U754 ( .A(w_mult_Z[25]), .B(n111), .C(w_add_Z[25]), .D(n121), .Y(
        N538) );
  scg2d1_hd U756 ( .A(w_mult_Z[26]), .B(n111), .C(w_add_Z[26]), .D(n121), .Y(
        N539) );
  scg2d1_hd U758 ( .A(w_mult_Z[27]), .B(n111), .C(w_add_Z[27]), .D(n121), .Y(
        N540) );
  scg2d1_hd U760 ( .A(w_mult_Z[28]), .B(n111), .C(w_add_Z[28]), .D(n121), .Y(
        N541) );
  scg2d1_hd U762 ( .A(w_mult_Z[29]), .B(n111), .C(w_add_Z[29]), .D(n121), .Y(
        N542) );
  scg2d1_hd U764 ( .A(w_mult_Z[30]), .B(n111), .C(w_add_Z[30]), .D(n121), .Y(
        N543) );
  scg2d1_hd U766 ( .A(w_mult_Z[31]), .B(n111), .C(w_add_Z[31]), .D(n121), .Y(
        N544) );
  or2d1_hd U768 ( .A(N27), .B(alt24_n19), .Y(N550) );
  clknd2d1_hd U771 ( .A(n100), .B(n101), .Y(N558) );
  or2d1_hd U773 ( .A(N39), .B(n541), .Y(N49) );
  or2d1_hd U775 ( .A(N39), .B(n544), .Y(N114) );
  clknd2d1_hd U776 ( .A(n107), .B(n108), .Y(N554) );
  ivd1_hd U777 ( .A(w_mult_Z_STB), .Y(N322) );
  mx2d1_hd U779 ( .D0(r_counter[1]), .D1(N376), .S(N552), .Y(n280) );
  xo2d1_hd U780 ( .A(r_counter[0]), .B(r_counter[1]), .Y(N319) );
  ad2d1_hd U782 ( .A(N27), .B(w_rstn), .Y(N559) );
  or3d1_hd U789 ( .A(n544), .B(n541), .C(n537), .Y(N563) );
  nr2d1_hd U791 ( .A(n104), .B(n103), .Y(n101) );
  ivd1_hd U1043 ( .A(n119), .Y(n535) );
  nr2d1_hd U1044 ( .A(n541), .B(alt24_n58), .Y(n537) );
  nr2d1_hd U1045 ( .A(N37), .B(r_counter[0]), .Y(n538) );
  nr2d1_hd U1046 ( .A(r_counter[1]), .B(N38), .Y(n540) );
  or4d1_hd U1050 ( .A(n536), .B(alt24_n19), .C(n103), .D(n120), .Y(n543) );
  clknd2d1_hd U1051 ( .A(o_Y_DATA_VALID), .B(i_Y_ACK), .Y(n545) );
  clknd2d1_hd U1052 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(n546) );
  ivd1_hd U1053 ( .A(N317), .Y(N320) );
  nr2d1_hd U1054 ( .A(n538), .B(alt24_n109), .Y(n547) );
  or2d1_hd U1055 ( .A(n538), .B(n547), .Y(N564) );
  ivd1_hd U1056 ( .A(N27), .Y(n113) );
  ivd1_hd U10 ( .A(n580), .Y(n287) );
  ivd1_hd U17 ( .A(n580), .Y(n294) );
  ivd1_hd U28 ( .A(n580), .Y(n305) );
  ivd1_hd U29 ( .A(n580), .Y(n306) );
  ivd1_hd U30 ( .A(n581), .Y(n307) );
  ivd1_hd U31 ( .A(n581), .Y(n308) );
  ivd1_hd U41 ( .A(n581), .Y(n318) );
  ivd1_hd U101 ( .A(n581), .Y(n378) );
  ivd1_hd U102 ( .A(n581), .Y(n379) );
  ivd1_hd U115 ( .A(n581), .Y(n392) );
  ivd1_hd U170 ( .A(n580), .Y(n436) );
  ivd1_hd U172 ( .A(n581), .Y(n438) );
  ivd1_hd U326 ( .A(n581), .Y(n469) );
  ivd1_hd U327 ( .A(n580), .Y(n470) );
  ivd1_hd U329 ( .A(n580), .Y(n472) );
  ivd1_hd U348 ( .A(n580), .Y(n491) );
  ivd1_hd U387 ( .A(n580), .Y(n530) );
  ivd1_hd U419 ( .A(w_rstn), .Y(n580) );
  ivd1_hd U420 ( .A(w_rstn), .Y(n581) );
  SNPS_CLOCK_GATE_HIGH_iir_hpf_11 clk_gate_o_Y_DATA_reg_31__0 ( .CLK(i_CLK), 
        .EN(N562), .ENCLK(n812), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_hpf_12 clk_gate_r_mult_A_reg_29__0 ( .CLK(i_CLK), 
        .EN(n865), .ENCLK(n811), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_hpf_13 clk_gate_r_add_B_reg_30__0 ( .CLK(i_CLK), 
        .EN(n931), .ENCLK(n810), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_iir_hpf_14 clk_gate_r_y_data_reg_31__0 ( .CLK(i_CLK), 
        .EN(n808), .ENCLK(n809), .TE(1'b0) );
  fd2qd1_hd r_pstate_reg_1_ ( .D(N554), .CK(i_CLK), .RN(n307), .Q(r_pstate[1])
         );
  fd2qd1_hd r_pstate_reg_0_ ( .D(n815), .CK(i_CLK), .RN(n305), .Q(r_pstate[0])
         );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n546), .E(N559), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_counter_reg_1_ ( .D(n280), .CK(i_CLK), .RN(n530), .Q(
        r_counter[1]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(o_Y_DATA[15]), .CK(n809), .RN(n472), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(o_Y_DATA[14]), .CK(n809), .RN(n306), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(o_Y_DATA[13]), .CK(n809), .RN(n436), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(o_Y_DATA[12]), .CK(n809), .RN(n307), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(o_Y_DATA[11]), .CK(n809), .RN(n472), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(o_Y_DATA[10]), .CK(n809), .RN(n438), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(o_Y_DATA[6]), .CK(n809), .RN(n307), .Q(
        r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(o_Y_DATA[5]), .CK(n809), .RN(n305), .Q(
        r_y_data[5]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(r_x_data[31]), .CK(n809), .RN(n308), .Q(
        r_x_data[63]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(r_x_data[30]), .CK(n809), .RN(n305), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(o_Y_DATA[31]), .CK(n809), .RN(n318), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(o_Y_DATA[30]), .CK(n809), .RN(n294), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(o_Y_DATA[29]), .CK(n809), .RN(n472), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(o_Y_DATA[28]), .CK(n809), .RN(n306), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(o_Y_DATA[27]), .CK(n809), .RN(n379), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(o_Y_DATA[26]), .CK(n809), .RN(n306), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(o_Y_DATA[25]), .CK(n809), .RN(n392), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(o_Y_DATA[24]), .CK(n809), .RN(n472), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(r_x_data[4]), .CK(n809), .RN(n306), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(r_x_data[3]), .CK(n809), .RN(n378), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(r_x_data[2]), .CK(n809), .RN(n379), .Q(
        r_x_data[34]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(r_x_data[1]), .CK(n809), .RN(n294), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_x_data_reg_32_ ( .D(r_x_data[0]), .CK(n809), .RN(n470), .Q(
        r_x_data[32]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(o_Y_DATA[9]), .CK(n809), .RN(n469), .Q(
        r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(o_Y_DATA[4]), .CK(n809), .RN(n305), .Q(
        r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(o_Y_DATA[3]), .CK(n809), .RN(n469), .Q(
        r_y_data[3]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(o_Y_DATA[22]), .CK(n809), .RN(n308), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(o_Y_DATA[21]), .CK(n809), .RN(n491), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(o_Y_DATA[20]), .CK(n809), .RN(n307), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(o_Y_DATA[19]), .CK(n809), .RN(n307), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(o_Y_DATA[18]), .CK(n809), .RN(n318), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(o_Y_DATA[17]), .CK(n809), .RN(n379), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(o_Y_DATA[16]), .CK(n809), .RN(n378), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(o_Y_DATA[8]), .CK(n809), .RN(n306), .Q(
        r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(o_Y_DATA[7]), .CK(n809), .RN(n436), .Q(
        r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_2_ ( .D(o_Y_DATA[2]), .CK(n809), .RN(n470), .Q(
        r_y_data[2]) );
  fd2qd1_hd r_y_data_reg_1_ ( .D(o_Y_DATA[1]), .CK(n809), .RN(n294), .Q(
        r_y_data[1]) );
  fd2qd1_hd r_y_data_reg_0_ ( .D(o_Y_DATA[0]), .CK(n809), .RN(n436), .Q(
        r_y_data[0]) );
  fd2qd1_hd r_mult_AB_STB_reg ( .D(n813), .CK(i_CLK), .RN(n305), .Q(
        r_mult_AB_STB) );
  fd2qd1_hd r_add_AB_STB_reg ( .D(n814), .CK(i_CLK), .RN(n378), .Q(
        r_add_AB_STB) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(o_Y_DATA[23]), .CK(n809), .RN(n305), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(r_x_data[29]), .CK(n809), .RN(n318), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(r_x_data[28]), .CK(n809), .RN(n469), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(r_x_data[27]), .CK(n809), .RN(n308), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(r_x_data[26]), .CK(n809), .RN(n491), .Q(
        r_x_data[58]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(r_x_data[25]), .CK(n809), .RN(n305), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(r_x_data[24]), .CK(n809), .RN(n307), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(r_x_data[23]), .CK(n809), .RN(n318), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(r_x_data[22]), .CK(n809), .RN(n469), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(r_x_data[21]), .CK(n809), .RN(n470), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(r_x_data[20]), .CK(n809), .RN(n378), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(r_x_data[19]), .CK(n809), .RN(n379), .Q(
        r_x_data[51]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(r_x_data[18]), .CK(n809), .RN(n287), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(r_x_data[17]), .CK(n809), .RN(n491), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(r_x_data[16]), .CK(n809), .RN(n469), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(r_x_data[15]), .CK(n809), .RN(n307), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(r_x_data[14]), .CK(n809), .RN(n305), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(r_x_data[13]), .CK(n809), .RN(n530), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(r_x_data[12]), .CK(n809), .RN(n287), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(r_x_data[11]), .CK(n809), .RN(n294), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(r_x_data[10]), .CK(n809), .RN(n530), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(r_x_data[9]), .CK(n809), .RN(n472), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(r_x_data[8]), .CK(n809), .RN(n530), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(r_x_data[7]), .CK(n809), .RN(n294), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(r_x_data[6]), .CK(n809), .RN(n470), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(r_x_data[5]), .CK(n809), .RN(n436), .Q(
        r_x_data[37]) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(N544), .CK(n812), .RN(n306), .Q(o_Y_DATA[31]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(N543), .CK(n812), .RN(n287), .Q(o_Y_DATA[30]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(N542), .CK(n812), .RN(n308), .Q(o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(N541), .CK(n812), .RN(n436), .Q(o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(N540), .CK(n812), .RN(n306), .Q(o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(N539), .CK(n812), .RN(n318), .Q(o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(N538), .CK(n812), .RN(n530), .Q(o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(N537), .CK(n812), .RN(n294), .Q(o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(N536), .CK(n812), .RN(n294), .Q(o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(N535), .CK(n812), .RN(n287), .Q(o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(N534), .CK(n812), .RN(n470), .Q(o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(N533), .CK(n812), .RN(n530), .Q(o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(N532), .CK(n812), .RN(n491), .Q(o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(N531), .CK(n812), .RN(n530), .Q(o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(N530), .CK(n812), .RN(n305), .Q(o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(N529), .CK(n812), .RN(n287), .Q(o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(N528), .CK(n812), .RN(n469), .Q(o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(N527), .CK(n812), .RN(n491), .Q(o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(N526), .CK(n812), .RN(n306), .Q(o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(N525), .CK(n812), .RN(n305), .Q(o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(N524), .CK(n812), .RN(n306), .Q(o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(N523), .CK(n812), .RN(n307), .Q(o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(N522), .CK(n812), .RN(n308), .Q(o_Y_DATA[9])
         );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(N521), .CK(n812), .RN(n491), .Q(o_Y_DATA[8])
         );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(N520), .CK(n812), .RN(n392), .Q(o_Y_DATA[7])
         );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(N519), .CK(n812), .RN(n438), .Q(o_Y_DATA[6])
         );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(N518), .CK(n812), .RN(n287), .Q(o_Y_DATA[5])
         );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(N517), .CK(n812), .RN(n294), .Q(o_Y_DATA[4])
         );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(N516), .CK(n812), .RN(n436), .Q(o_Y_DATA[3])
         );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(N515), .CK(n812), .RN(n308), .Q(o_Y_DATA[2])
         );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(N514), .CK(n812), .RN(n470), .Q(o_Y_DATA[1])
         );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(N513), .CK(n812), .RN(n470), .Q(o_Y_DATA[0])
         );
  fd2qd1_hd r_mult_B_reg_31_ ( .D(n861), .CK(n811), .RN(n469), .Q(r_mult_B[31]) );
  fd2qd1_hd r_mult_B_reg_30_ ( .D(n860), .CK(n811), .RN(n436), .Q(r_mult_B[30]) );
  fd2qd1_hd r_mult_B_reg_29_ ( .D(n859), .CK(n811), .RN(n307), .Q(r_mult_B[29]) );
  fd2qd1_hd r_mult_B_reg_28_ ( .D(n858), .CK(n811), .RN(n438), .Q(r_mult_B[28]) );
  fd2qd1_hd r_mult_B_reg_27_ ( .D(n857), .CK(n811), .RN(n287), .Q(r_mult_B[27]) );
  fd2qd1_hd r_mult_B_reg_26_ ( .D(n856), .CK(n811), .RN(n287), .Q(r_mult_B[26]) );
  fd2qd1_hd r_mult_B_reg_25_ ( .D(n855), .CK(n811), .RN(n294), .Q(r_mult_B[25]) );
  fd2qd1_hd r_mult_B_reg_24_ ( .D(n854), .CK(n811), .RN(n378), .Q(r_mult_B[24]) );
  fd2qd1_hd r_mult_B_reg_23_ ( .D(n853), .CK(n811), .RN(n436), .Q(r_mult_B[23]) );
  fd2qd1_hd r_mult_B_reg_22_ ( .D(n852), .CK(n811), .RN(n379), .Q(r_mult_B[22]) );
  fd2qd1_hd r_mult_B_reg_21_ ( .D(n851), .CK(n811), .RN(n530), .Q(r_mult_B[21]) );
  fd2qd1_hd r_mult_B_reg_20_ ( .D(n850), .CK(n811), .RN(n438), .Q(r_mult_B[20]) );
  fd2qd1_hd r_mult_B_reg_19_ ( .D(n849), .CK(n811), .RN(n378), .Q(r_mult_B[19]) );
  fd2qd1_hd r_mult_B_reg_18_ ( .D(n848), .CK(n811), .RN(n392), .Q(r_mult_B[18]) );
  fd2qd1_hd r_mult_B_reg_17_ ( .D(n847), .CK(n811), .RN(n392), .Q(r_mult_B[17]) );
  fd2qd1_hd r_mult_B_reg_16_ ( .D(n846), .CK(n811), .RN(n470), .Q(r_mult_B[16]) );
  fd2qd1_hd r_mult_B_reg_15_ ( .D(n845), .CK(n811), .RN(n378), .Q(r_mult_B[15]) );
  fd2qd1_hd r_mult_B_reg_14_ ( .D(n844), .CK(n811), .RN(n469), .Q(r_mult_B[14]) );
  fd2qd1_hd r_mult_B_reg_13_ ( .D(n843), .CK(n811), .RN(n294), .Q(r_mult_B[13]) );
  fd2qd1_hd r_mult_B_reg_12_ ( .D(n842), .CK(n811), .RN(n305), .Q(r_mult_B[12]) );
  fd2qd1_hd r_mult_B_reg_11_ ( .D(n841), .CK(n811), .RN(n436), .Q(r_mult_B[11]) );
  fd2qd1_hd r_mult_B_reg_10_ ( .D(n840), .CK(n811), .RN(n469), .Q(r_mult_B[10]) );
  fd2qd1_hd r_mult_B_reg_9_ ( .D(n839), .CK(n811), .RN(n308), .Q(r_mult_B[9])
         );
  fd2qd1_hd r_mult_B_reg_8_ ( .D(n838), .CK(n811), .RN(n318), .Q(r_mult_B[8])
         );
  fd2qd1_hd r_mult_B_reg_7_ ( .D(n837), .CK(n811), .RN(n287), .Q(r_mult_B[7])
         );
  fd2qd1_hd r_mult_B_reg_6_ ( .D(n836), .CK(n811), .RN(n469), .Q(r_mult_B[6])
         );
  fd2qd1_hd r_mult_B_reg_5_ ( .D(n835), .CK(n811), .RN(n469), .Q(r_mult_B[5])
         );
  fd2qd1_hd r_mult_B_reg_4_ ( .D(n834), .CK(n811), .RN(n491), .Q(r_mult_B[4])
         );
  fd2qd1_hd r_mult_B_reg_3_ ( .D(n833), .CK(n811), .RN(n491), .Q(r_mult_B[3])
         );
  fd2qd1_hd r_mult_B_reg_2_ ( .D(n832), .CK(n811), .RN(n438), .Q(r_mult_B[2])
         );
  fd2qd1_hd r_mult_B_reg_1_ ( .D(n831), .CK(n811), .RN(n472), .Q(r_mult_B[1])
         );
  fd2qd1_hd r_mult_B_reg_0_ ( .D(n830), .CK(n811), .RN(n392), .Q(r_mult_B[0])
         );
  fd2qd1_hd r_add_B_reg_30_ ( .D(n929), .CK(n810), .RN(n294), .Q(r_add_B[30])
         );
  fd2qd1_hd r_add_B_reg_29_ ( .D(n928), .CK(n810), .RN(n294), .Q(r_add_B[29])
         );
  fd2qd1_hd r_add_B_reg_28_ ( .D(n927), .CK(n810), .RN(n469), .Q(r_add_B[28])
         );
  fd2qd1_hd r_add_B_reg_27_ ( .D(n926), .CK(n810), .RN(n470), .Q(r_add_B[27])
         );
  fd2qd1_hd r_add_B_reg_26_ ( .D(n925), .CK(n810), .RN(n530), .Q(r_add_B[26])
         );
  fd2qd1_hd r_add_B_reg_25_ ( .D(n924), .CK(n810), .RN(n472), .Q(r_add_B[25])
         );
  fd2qd1_hd r_add_B_reg_24_ ( .D(n923), .CK(n810), .RN(n472), .Q(r_add_B[24])
         );
  fd2qd1_hd r_add_B_reg_23_ ( .D(n922), .CK(n810), .RN(n294), .Q(r_add_B[23])
         );
  fd2qd1_hd r_add_B_reg_22_ ( .D(n921), .CK(n810), .RN(n305), .Q(r_add_B[22])
         );
  fd2qd1_hd r_add_B_reg_21_ ( .D(n920), .CK(n810), .RN(n392), .Q(r_add_B[21])
         );
  fd2qd1_hd r_add_B_reg_20_ ( .D(n919), .CK(n810), .RN(n469), .Q(r_add_B[20])
         );
  fd2qd1_hd r_add_B_reg_19_ ( .D(n918), .CK(n810), .RN(n491), .Q(r_add_B[19])
         );
  fd2qd1_hd r_add_B_reg_18_ ( .D(n917), .CK(n810), .RN(n287), .Q(r_add_B[18])
         );
  fd2qd1_hd r_add_B_reg_17_ ( .D(n916), .CK(n810), .RN(n530), .Q(r_add_B[17])
         );
  fd2qd1_hd r_add_B_reg_16_ ( .D(n915), .CK(n810), .RN(n472), .Q(r_add_B[16])
         );
  fd2qd1_hd r_add_B_reg_15_ ( .D(n914), .CK(n810), .RN(n318), .Q(r_add_B[15])
         );
  fd2qd1_hd r_add_B_reg_14_ ( .D(n913), .CK(n810), .RN(n308), .Q(r_add_B[14])
         );
  fd2qd1_hd r_add_B_reg_13_ ( .D(n912), .CK(n810), .RN(n378), .Q(r_add_B[13])
         );
  fd2qd1_hd r_add_B_reg_12_ ( .D(n911), .CK(n810), .RN(n287), .Q(r_add_B[12])
         );
  fd2qd1_hd r_add_B_reg_11_ ( .D(n910), .CK(n810), .RN(n436), .Q(r_add_B[11])
         );
  fd2qd1_hd r_add_B_reg_10_ ( .D(n909), .CK(n810), .RN(n392), .Q(r_add_B[10])
         );
  fd2qd1_hd r_add_B_reg_9_ ( .D(n908), .CK(n810), .RN(n436), .Q(r_add_B[9]) );
  fd2qd1_hd r_add_B_reg_8_ ( .D(n907), .CK(n810), .RN(n472), .Q(r_add_B[8]) );
  fd2qd1_hd r_add_B_reg_7_ ( .D(n906), .CK(n810), .RN(n438), .Q(r_add_B[7]) );
  fd2qd1_hd r_add_B_reg_6_ ( .D(n905), .CK(n810), .RN(n491), .Q(r_add_B[6]) );
  fd2qd1_hd r_add_B_reg_5_ ( .D(n904), .CK(n810), .RN(n469), .Q(r_add_B[5]) );
  fd2qd1_hd r_add_B_reg_4_ ( .D(n903), .CK(n810), .RN(n294), .Q(r_add_B[4]) );
  fd2qd1_hd r_add_B_reg_3_ ( .D(n902), .CK(n810), .RN(n472), .Q(r_add_B[3]) );
  fd2qd1_hd r_add_B_reg_2_ ( .D(n901), .CK(n810), .RN(n392), .Q(r_add_B[2]) );
  fd2qd1_hd r_add_B_reg_1_ ( .D(n900), .CK(n810), .RN(n287), .Q(r_add_B[1]) );
  fd2qd1_hd r_add_B_reg_0_ ( .D(n899), .CK(n810), .RN(n438), .Q(r_add_B[0]) );
  fd2qd1_hd r_add_A_reg_31_ ( .D(n898), .CK(n810), .RN(n491), .Q(r_add_A[31])
         );
  fd2qd1_hd r_add_A_reg_30_ ( .D(n897), .CK(n810), .RN(n306), .Q(r_add_A[30])
         );
  fd2qd1_hd r_add_A_reg_29_ ( .D(n896), .CK(n810), .RN(n308), .Q(r_add_A[29])
         );
  fd2qd1_hd r_add_A_reg_28_ ( .D(n895), .CK(n810), .RN(n287), .Q(r_add_A[28])
         );
  fd2qd1_hd r_add_A_reg_27_ ( .D(n894), .CK(n810), .RN(n308), .Q(r_add_A[27])
         );
  fd2qd1_hd r_add_A_reg_26_ ( .D(n893), .CK(n810), .RN(n438), .Q(r_add_A[26])
         );
  fd2qd1_hd r_add_A_reg_25_ ( .D(n892), .CK(n810), .RN(n438), .Q(r_add_A[25])
         );
  fd2qd1_hd r_add_A_reg_24_ ( .D(n891), .CK(n810), .RN(n379), .Q(r_add_A[24])
         );
  fd2qd1_hd r_add_A_reg_23_ ( .D(n890), .CK(n810), .RN(n491), .Q(r_add_A[23])
         );
  fd2qd1_hd r_add_A_reg_22_ ( .D(n889), .CK(n810), .RN(n436), .Q(r_add_A[22])
         );
  fd2qd1_hd r_add_A_reg_21_ ( .D(n888), .CK(n810), .RN(n470), .Q(r_add_A[21])
         );
  fd2qd1_hd r_add_A_reg_20_ ( .D(n887), .CK(n810), .RN(n378), .Q(r_add_A[20])
         );
  fd2qd1_hd r_add_A_reg_19_ ( .D(n886), .CK(n810), .RN(n379), .Q(r_add_A[19])
         );
  fd2qd1_hd r_add_A_reg_18_ ( .D(n885), .CK(n810), .RN(n305), .Q(r_add_A[18])
         );
  fd2qd1_hd r_add_A_reg_17_ ( .D(n884), .CK(n810), .RN(n470), .Q(r_add_A[17])
         );
  fd2qd1_hd r_add_A_reg_16_ ( .D(n883), .CK(n810), .RN(n379), .Q(r_add_A[16])
         );
  fd2qd1_hd r_add_A_reg_15_ ( .D(n882), .CK(n810), .RN(n378), .Q(r_add_A[15])
         );
  fd2qd1_hd r_add_A_reg_14_ ( .D(n881), .CK(n810), .RN(n308), .Q(r_add_A[14])
         );
  fd2qd1_hd r_add_A_reg_13_ ( .D(n880), .CK(n810), .RN(n379), .Q(r_add_A[13])
         );
  fd2qd1_hd r_add_A_reg_12_ ( .D(n879), .CK(n810), .RN(n305), .Q(r_add_A[12])
         );
  fd2qd1_hd r_add_A_reg_11_ ( .D(n878), .CK(n810), .RN(n378), .Q(r_add_A[11])
         );
  fd2qd1_hd r_add_A_reg_10_ ( .D(n877), .CK(n810), .RN(n306), .Q(r_add_A[10])
         );
  fd2qd1_hd r_add_A_reg_9_ ( .D(n876), .CK(n810), .RN(n379), .Q(r_add_A[9]) );
  fd2qd1_hd r_add_A_reg_8_ ( .D(n875), .CK(n810), .RN(n305), .Q(r_add_A[8]) );
  fd2qd1_hd r_add_A_reg_7_ ( .D(n874), .CK(n810), .RN(n307), .Q(r_add_A[7]) );
  fd2qd1_hd r_add_A_reg_6_ ( .D(n873), .CK(n810), .RN(n318), .Q(r_add_A[6]) );
  fd2qd1_hd r_add_A_reg_5_ ( .D(n872), .CK(n810), .RN(n379), .Q(r_add_A[5]) );
  fd2qd1_hd r_add_A_reg_4_ ( .D(n871), .CK(n810), .RN(n378), .Q(r_add_A[4]) );
  fd2qd1_hd r_add_A_reg_3_ ( .D(n870), .CK(n810), .RN(n306), .Q(r_add_A[3]) );
  fd2qd1_hd r_add_A_reg_2_ ( .D(n869), .CK(n810), .RN(n436), .Q(r_add_A[2]) );
  fd2qd1_hd r_add_A_reg_1_ ( .D(n868), .CK(n810), .RN(n470), .Q(r_add_A[1]) );
  fd2qd1_hd r_add_A_reg_0_ ( .D(n867), .CK(n810), .RN(n294), .Q(r_add_A[0]) );
  fd2qd1_hd r_mult_Z_ACK_reg ( .D(n816), .CK(i_CLK), .RN(n491), .Q(
        r_mult_Z_ACK) );
  fd2qd1_hd r_add_Z_ACK_reg ( .D(n818), .CK(i_CLK), .RN(n438), .Q(r_add_Z_ACK)
         );
  fd2qd1_hd r_add_B_reg_31_ ( .D(n866), .CK(n810), .RN(n530), .Q(r_add_B[31])
         );
  fd2qd1_hd r_x_data_reg_31_ ( .D(i_X_DATA[31]), .CK(n809), .RN(n318), .Q(
        r_x_data[31]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(i_X_DATA[30]), .CK(n809), .RN(n530), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(i_X_DATA[29]), .CK(n809), .RN(n306), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(i_X_DATA[28]), .CK(n809), .RN(n378), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(i_X_DATA[27]), .CK(n809), .RN(n379), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(i_X_DATA[26]), .CK(n809), .RN(n318), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(i_X_DATA[25]), .CK(n809), .RN(n307), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(i_X_DATA[24]), .CK(n809), .RN(n469), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(i_X_DATA[23]), .CK(n809), .RN(n307), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(i_X_DATA[22]), .CK(n809), .RN(n392), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(i_X_DATA[21]), .CK(n809), .RN(n392), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(i_X_DATA[20]), .CK(n809), .RN(n318), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(i_X_DATA[19]), .CK(n809), .RN(n379), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(i_X_DATA[18]), .CK(n809), .RN(n378), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(i_X_DATA[17]), .CK(n809), .RN(n306), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(i_X_DATA[16]), .CK(n809), .RN(n308), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(i_X_DATA[15]), .CK(n809), .RN(n470), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(i_X_DATA[14]), .CK(n809), .RN(n308), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(i_X_DATA[13]), .CK(n809), .RN(n308), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(i_X_DATA[12]), .CK(n809), .RN(n287), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(i_X_DATA[11]), .CK(n809), .RN(n530), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(i_X_DATA[10]), .CK(n809), .RN(n438), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(i_X_DATA[9]), .CK(n809), .RN(n472), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(i_X_DATA[8]), .CK(n809), .RN(n392), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(i_X_DATA[7]), .CK(n809), .RN(n392), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(i_X_DATA[6]), .CK(n809), .RN(n318), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(i_X_DATA[5]), .CK(n809), .RN(n379), .Q(
        r_x_data[5]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(i_X_DATA[4]), .CK(n809), .RN(n472), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(i_X_DATA[3]), .CK(n809), .RN(n491), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(i_X_DATA[2]), .CK(n809), .RN(n530), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(i_X_DATA[1]), .CK(n809), .RN(n318), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(i_X_DATA[0]), .CK(n809), .RN(n307), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_counter_reg_0_ ( .D(n817), .CK(i_CLK), .RN(n470), .Q(
        r_counter[0]) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n819), .CK(i_CLK), .RN(n491), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_mult_A_reg_29_ ( .D(n863), .CK(n811), .RN(n378), .Q(r_mult_A[29]) );
  fd2qd1_hd r_mult_A_reg_28_ ( .D(n863), .CK(n811), .RN(n379), .Q(r_mult_A[28]) );
  fd2qd1_hd r_mult_A_reg_27_ ( .D(n863), .CK(n811), .RN(n530), .Q(r_mult_A[27]) );
  fd2qd1_hd r_mult_A_reg_26_ ( .D(n862), .CK(n811), .RN(n438), .Q(r_mult_A[26]) );
  fd2qd1_hd r_mult_A_reg_25_ ( .D(n863), .CK(n811), .RN(n438), .Q(r_mult_A[25]) );
  fd2qd1_hd r_mult_A_reg_24_ ( .D(n863), .CK(n811), .RN(n392), .Q(r_mult_A[24]) );
  fd2qd1_hd r_mult_A_reg_22_ ( .D(n862), .CK(n811), .RN(n307), .Q(r_mult_A[22]) );
  fd2qd1_hd r_mult_A_reg_21_ ( .D(n862), .CK(n811), .RN(n308), .Q(r_mult_A[21]) );
  fd2qd1_hd r_mult_A_reg_17_ ( .D(n863), .CK(n811), .RN(n287), .Q(r_mult_A[17]) );
  fd2qd1_hd r_mult_A_reg_16_ ( .D(n862), .CK(n811), .RN(n438), .Q(r_mult_A[16]) );
  fd2qd1_hd r_mult_A_reg_14_ ( .D(n863), .CK(n811), .RN(n438), .Q(r_mult_A[14]) );
  fd2qd1_hd r_mult_A_reg_13_ ( .D(n863), .CK(n811), .RN(n472), .Q(r_mult_A[13]) );
  fd2qd1_hd r_mult_A_reg_11_ ( .D(n863), .CK(n811), .RN(n472), .Q(r_mult_A[11]) );
  fd2qd1_hd r_mult_A_reg_9_ ( .D(n863), .CK(n811), .RN(n392), .Q(r_mult_A[9])
         );
  fd2qd1_hd r_mult_A_reg_8_ ( .D(n862), .CK(n811), .RN(n436), .Q(r_mult_A[8])
         );
  fd2qd1_hd r_mult_A_reg_7_ ( .D(n862), .CK(n811), .RN(n470), .Q(r_mult_A[7])
         );
  fd2qd1_hd r_mult_A_reg_6_ ( .D(n862), .CK(n811), .RN(n392), .Q(r_mult_A[6])
         );
  fd2qd1_hd r_mult_A_reg_5_ ( .D(n863), .CK(n811), .RN(n318), .Q(r_mult_A[5])
         );
  fd2qd1_hd r_mult_A_reg_1_ ( .D(n862), .CK(n811), .RN(n318), .Q(r_mult_A[1])
         );
  fd2qd1_hd r_mult_A_reg_0_ ( .D(n862), .CK(n811), .RN(n307), .Q(r_mult_A[0])
         );
  ivd1_hd U1 ( .A(r_counter[1]), .Y(N37) );
  clknd2d1_hd U2 ( .A(r_pstate[1]), .B(n545), .Y(n823) );
  clknd2d1_hd U3 ( .A(n546), .B(n539), .Y(n822) );
  mx2d1_hd U4 ( .D0(n825), .D1(n102), .S(N28), .Y(n931) );
  scg20d1_hd U5 ( .A(n539), .B(N563), .C(N28), .Y(n123) );
  ad2d1_hd U6 ( .A(n543), .B(alt24_n18), .Y(N562) );
  mx2d1_hd U7 ( .D0(o_Y_DATA_VALID), .D1(N371), .S(N550), .Y(n819) );
  mx2d1_hd U8 ( .D0(r_counter[0]), .D1(N374), .S(N552), .Y(n817) );
  scg2d1_hd U9 ( .A(o_Y_DATA[31]), .B(n807), .C(n536), .D(n824), .Y(n866) );
  mx2d1_hd U11 ( .D0(r_add_Z_ACK), .D1(n807), .S(N558), .Y(n818) );
  mx2d1_hd U12 ( .D0(r_mult_Z_ACK), .D1(n807), .S(N557), .Y(n816) );
  scg2d1_hd U13 ( .A(n536), .B(r_x_data[0]), .C(n807), .D(w_mult_Z[0]), .Y(
        n867) );
  scg2d1_hd U14 ( .A(n536), .B(r_x_data[1]), .C(n807), .D(w_mult_Z[1]), .Y(
        n868) );
  scg2d1_hd U15 ( .A(n536), .B(r_x_data[2]), .C(n807), .D(w_mult_Z[2]), .Y(
        n869) );
  scg2d1_hd U16 ( .A(n536), .B(r_x_data[3]), .C(n807), .D(w_mult_Z[3]), .Y(
        n870) );
  scg2d1_hd U18 ( .A(n536), .B(r_x_data[4]), .C(n807), .D(w_mult_Z[4]), .Y(
        n871) );
  scg2d1_hd U19 ( .A(n536), .B(r_x_data[5]), .C(n807), .D(w_mult_Z[5]), .Y(
        n872) );
  scg2d1_hd U20 ( .A(n536), .B(r_x_data[6]), .C(n807), .D(w_mult_Z[6]), .Y(
        n873) );
  scg2d1_hd U21 ( .A(n536), .B(r_x_data[7]), .C(n807), .D(w_mult_Z[7]), .Y(
        n874) );
  scg2d1_hd U22 ( .A(n536), .B(r_x_data[8]), .C(n807), .D(w_mult_Z[8]), .Y(
        n875) );
  scg2d1_hd U23 ( .A(n536), .B(r_x_data[9]), .C(n807), .D(w_mult_Z[9]), .Y(
        n876) );
  scg2d1_hd U24 ( .A(n536), .B(r_x_data[10]), .C(n807), .D(w_mult_Z[10]), .Y(
        n877) );
  scg2d1_hd U25 ( .A(n536), .B(r_x_data[11]), .C(n807), .D(w_mult_Z[11]), .Y(
        n878) );
  scg2d1_hd U26 ( .A(n536), .B(r_x_data[12]), .C(n807), .D(w_mult_Z[12]), .Y(
        n879) );
  scg2d1_hd U27 ( .A(n536), .B(r_x_data[13]), .C(n807), .D(w_mult_Z[13]), .Y(
        n880) );
  scg2d1_hd U32 ( .A(n536), .B(r_x_data[14]), .C(n807), .D(w_mult_Z[14]), .Y(
        n881) );
  scg2d1_hd U33 ( .A(n536), .B(r_x_data[15]), .C(n807), .D(w_mult_Z[15]), .Y(
        n882) );
  scg2d1_hd U34 ( .A(n536), .B(r_x_data[16]), .C(n807), .D(w_mult_Z[16]), .Y(
        n883) );
  scg2d1_hd U35 ( .A(n536), .B(r_x_data[17]), .C(n807), .D(w_mult_Z[17]), .Y(
        n884) );
  scg2d1_hd U36 ( .A(n536), .B(r_x_data[18]), .C(n807), .D(w_mult_Z[18]), .Y(
        n885) );
  scg2d1_hd U37 ( .A(n536), .B(r_x_data[19]), .C(n807), .D(w_mult_Z[19]), .Y(
        n886) );
  scg2d1_hd U38 ( .A(n536), .B(r_x_data[20]), .C(n807), .D(w_mult_Z[20]), .Y(
        n887) );
  scg2d1_hd U39 ( .A(n536), .B(r_x_data[21]), .C(n807), .D(w_mult_Z[21]), .Y(
        n888) );
  scg2d1_hd U40 ( .A(n536), .B(r_x_data[22]), .C(n807), .D(w_mult_Z[22]), .Y(
        n889) );
  scg2d1_hd U42 ( .A(n536), .B(r_x_data[23]), .C(n807), .D(w_mult_Z[23]), .Y(
        n890) );
  scg2d1_hd U43 ( .A(n536), .B(r_x_data[24]), .C(n807), .D(w_mult_Z[24]), .Y(
        n891) );
  scg2d1_hd U44 ( .A(n536), .B(r_x_data[25]), .C(n807), .D(w_mult_Z[25]), .Y(
        n892) );
  scg2d1_hd U45 ( .A(n536), .B(r_x_data[26]), .C(n807), .D(w_mult_Z[26]), .Y(
        n893) );
  scg2d1_hd U46 ( .A(n536), .B(r_x_data[27]), .C(n807), .D(w_mult_Z[27]), .Y(
        n894) );
  scg2d1_hd U47 ( .A(n536), .B(r_x_data[28]), .C(n807), .D(w_mult_Z[28]), .Y(
        n895) );
  scg2d1_hd U48 ( .A(n536), .B(r_x_data[29]), .C(n807), .D(w_mult_Z[29]), .Y(
        n896) );
  scg2d1_hd U49 ( .A(n536), .B(r_x_data[30]), .C(n807), .D(w_mult_Z[30]), .Y(
        n897) );
  scg2d1_hd U50 ( .A(n536), .B(r_x_data[31]), .C(n807), .D(w_mult_Z[31]), .Y(
        n898) );
  scg2d1_hd U51 ( .A(n536), .B(r_x_data[32]), .C(n807), .D(o_Y_DATA[0]), .Y(
        n899) );
  scg2d1_hd U52 ( .A(n536), .B(r_x_data[33]), .C(n807), .D(o_Y_DATA[1]), .Y(
        n900) );
  scg2d1_hd U53 ( .A(n536), .B(r_x_data[34]), .C(n807), .D(o_Y_DATA[2]), .Y(
        n901) );
  scg2d1_hd U54 ( .A(n536), .B(r_x_data[35]), .C(n807), .D(o_Y_DATA[3]), .Y(
        n902) );
  scg2d1_hd U55 ( .A(n536), .B(r_x_data[36]), .C(n807), .D(o_Y_DATA[4]), .Y(
        n903) );
  scg2d1_hd U56 ( .A(n536), .B(r_x_data[37]), .C(n807), .D(o_Y_DATA[5]), .Y(
        n904) );
  scg2d1_hd U57 ( .A(n536), .B(r_x_data[38]), .C(n807), .D(o_Y_DATA[6]), .Y(
        n905) );
  scg2d1_hd U58 ( .A(n536), .B(r_x_data[39]), .C(n807), .D(o_Y_DATA[7]), .Y(
        n906) );
  scg2d1_hd U59 ( .A(n536), .B(r_x_data[40]), .C(n807), .D(o_Y_DATA[8]), .Y(
        n907) );
  scg2d1_hd U60 ( .A(n536), .B(r_x_data[41]), .C(n807), .D(o_Y_DATA[9]), .Y(
        n908) );
  scg2d1_hd U61 ( .A(n536), .B(r_x_data[42]), .C(n807), .D(o_Y_DATA[10]), .Y(
        n909) );
  scg2d1_hd U62 ( .A(n536), .B(r_x_data[43]), .C(n807), .D(o_Y_DATA[11]), .Y(
        n910) );
  scg2d1_hd U63 ( .A(n536), .B(r_x_data[44]), .C(n807), .D(o_Y_DATA[12]), .Y(
        n911) );
  scg2d1_hd U64 ( .A(n536), .B(r_x_data[45]), .C(n807), .D(o_Y_DATA[13]), .Y(
        n912) );
  scg2d1_hd U65 ( .A(n536), .B(r_x_data[46]), .C(n807), .D(o_Y_DATA[14]), .Y(
        n913) );
  scg2d1_hd U66 ( .A(n536), .B(r_x_data[47]), .C(n807), .D(o_Y_DATA[15]), .Y(
        n914) );
  scg2d1_hd U67 ( .A(n536), .B(r_x_data[48]), .C(n807), .D(o_Y_DATA[16]), .Y(
        n915) );
  scg2d1_hd U68 ( .A(n536), .B(r_x_data[49]), .C(n807), .D(o_Y_DATA[17]), .Y(
        n916) );
  scg2d1_hd U69 ( .A(n536), .B(r_x_data[50]), .C(n807), .D(o_Y_DATA[18]), .Y(
        n917) );
  scg2d1_hd U70 ( .A(n536), .B(r_x_data[51]), .C(n807), .D(o_Y_DATA[19]), .Y(
        n918) );
  scg2d1_hd U71 ( .A(n536), .B(r_x_data[52]), .C(n807), .D(o_Y_DATA[20]), .Y(
        n919) );
  scg2d1_hd U72 ( .A(n536), .B(r_x_data[53]), .C(n807), .D(o_Y_DATA[21]), .Y(
        n920) );
  scg2d1_hd U73 ( .A(n536), .B(r_x_data[54]), .C(n807), .D(o_Y_DATA[22]), .Y(
        n921) );
  scg2d1_hd U74 ( .A(n536), .B(r_x_data[55]), .C(n807), .D(o_Y_DATA[23]), .Y(
        n922) );
  scg2d1_hd U75 ( .A(n536), .B(r_x_data[56]), .C(n807), .D(o_Y_DATA[24]), .Y(
        n923) );
  scg2d1_hd U76 ( .A(n536), .B(r_x_data[57]), .C(n807), .D(o_Y_DATA[25]), .Y(
        n924) );
  scg2d1_hd U77 ( .A(n536), .B(r_x_data[58]), .C(n807), .D(o_Y_DATA[26]), .Y(
        n925) );
  scg2d1_hd U78 ( .A(n536), .B(r_x_data[59]), .C(n807), .D(o_Y_DATA[27]), .Y(
        n926) );
  scg2d1_hd U79 ( .A(n536), .B(r_x_data[60]), .C(n807), .D(o_Y_DATA[28]), .Y(
        n927) );
  scg2d1_hd U80 ( .A(n536), .B(r_x_data[61]), .C(n807), .D(o_Y_DATA[29]), .Y(
        n928) );
  scg2d1_hd U81 ( .A(n536), .B(r_x_data[62]), .C(n807), .D(o_Y_DATA[30]), .Y(
        n929) );
  scg2d1_hd U82 ( .A(n536), .B(r_y_data[0]), .C(n807), .D(w_add_Z[0]), .Y(n830) );
  scg2d1_hd U83 ( .A(n536), .B(r_y_data[1]), .C(n807), .D(w_add_Z[1]), .Y(n831) );
  scg2d1_hd U84 ( .A(n536), .B(r_y_data[2]), .C(n807), .D(w_add_Z[2]), .Y(n832) );
  scg2d1_hd U85 ( .A(n536), .B(r_y_data[3]), .C(n807), .D(w_add_Z[3]), .Y(n833) );
  scg2d1_hd U86 ( .A(n536), .B(r_y_data[4]), .C(n807), .D(w_add_Z[4]), .Y(n834) );
  scg2d1_hd U87 ( .A(n536), .B(r_y_data[5]), .C(n807), .D(w_add_Z[5]), .Y(n835) );
  scg2d1_hd U88 ( .A(n536), .B(r_y_data[6]), .C(n807), .D(w_add_Z[6]), .Y(n836) );
  scg2d1_hd U89 ( .A(n536), .B(r_y_data[7]), .C(n807), .D(w_add_Z[7]), .Y(n837) );
  scg2d1_hd U90 ( .A(n536), .B(r_y_data[8]), .C(n807), .D(w_add_Z[8]), .Y(n838) );
  scg2d1_hd U91 ( .A(n536), .B(r_y_data[9]), .C(n807), .D(w_add_Z[9]), .Y(n839) );
  scg2d1_hd U92 ( .A(n536), .B(r_y_data[10]), .C(n807), .D(w_add_Z[10]), .Y(
        n840) );
  scg2d1_hd U93 ( .A(n536), .B(r_y_data[11]), .C(n807), .D(w_add_Z[11]), .Y(
        n841) );
  scg2d1_hd U94 ( .A(n536), .B(r_y_data[12]), .C(n807), .D(w_add_Z[12]), .Y(
        n842) );
  scg2d1_hd U95 ( .A(n536), .B(r_y_data[13]), .C(n807), .D(w_add_Z[13]), .Y(
        n843) );
  scg2d1_hd U96 ( .A(n536), .B(r_y_data[14]), .C(n807), .D(w_add_Z[14]), .Y(
        n844) );
  scg2d1_hd U97 ( .A(n536), .B(r_y_data[15]), .C(n807), .D(w_add_Z[15]), .Y(
        n845) );
  scg2d1_hd U98 ( .A(n536), .B(r_y_data[16]), .C(n807), .D(w_add_Z[16]), .Y(
        n846) );
  scg2d1_hd U99 ( .A(n536), .B(r_y_data[17]), .C(n807), .D(w_add_Z[17]), .Y(
        n847) );
  scg2d1_hd U100 ( .A(n536), .B(r_y_data[18]), .C(n807), .D(w_add_Z[18]), .Y(
        n848) );
  scg2d1_hd U103 ( .A(n536), .B(r_y_data[19]), .C(n807), .D(w_add_Z[19]), .Y(
        n849) );
  scg2d1_hd U104 ( .A(n536), .B(r_y_data[20]), .C(n807), .D(w_add_Z[20]), .Y(
        n850) );
  scg2d1_hd U105 ( .A(n536), .B(r_y_data[21]), .C(n807), .D(w_add_Z[21]), .Y(
        n851) );
  scg2d1_hd U106 ( .A(n536), .B(r_y_data[22]), .C(n807), .D(w_add_Z[22]), .Y(
        n852) );
  scg2d1_hd U107 ( .A(n536), .B(r_y_data[23]), .C(n807), .D(w_add_Z[23]), .Y(
        n853) );
  scg2d1_hd U108 ( .A(n536), .B(r_y_data[24]), .C(n807), .D(w_add_Z[24]), .Y(
        n854) );
  scg2d1_hd U109 ( .A(n536), .B(r_y_data[25]), .C(n807), .D(w_add_Z[25]), .Y(
        n855) );
  scg2d1_hd U110 ( .A(n536), .B(r_y_data[26]), .C(n807), .D(w_add_Z[26]), .Y(
        n856) );
  scg2d1_hd U111 ( .A(n536), .B(r_y_data[27]), .C(n807), .D(w_add_Z[27]), .Y(
        n857) );
  scg2d1_hd U112 ( .A(n536), .B(r_y_data[28]), .C(n807), .D(w_add_Z[28]), .Y(
        n858) );
  scg2d1_hd U113 ( .A(n536), .B(r_y_data[29]), .C(n807), .D(w_add_Z[29]), .Y(
        n859) );
  scg2d1_hd U114 ( .A(n536), .B(r_y_data[30]), .C(n807), .D(w_add_Z[30]), .Y(
        n860) );
  scg2d1_hd U117 ( .A(n536), .B(r_y_data[31]), .C(n807), .D(w_add_Z[31]), .Y(
        n861) );
  mx2d1_hd U118 ( .D0(r_add_AB_STB), .D1(N546), .S(N548), .Y(n814) );
  mx2d1_hd U119 ( .D0(r_mult_AB_STB), .D1(N511), .S(N548), .Y(n813) );
  mx2d1_hd U121 ( .D0(r_pstate[0]), .D1(n827), .S(n828), .Y(n815) );
  clknd2d1_hd U125 ( .A(n820), .B(n821), .Y(n827) );
  nr2d1_hd U126 ( .A(n536), .B(n807), .Y(n124) );
  or2d1_hd U127 ( .A(N25), .B(r_pstate[0]), .Y(n805) );
  nid1_hd U128 ( .A(w_rst), .Y(n806) );
  ivd6_hd U129 ( .A(n805), .Y(n807) );
  ivd6_hd U131 ( .A(n535), .Y(n536) );
  ivd1_hd U132 ( .A(n124), .Y(n863) );
  ivd1_hd U133 ( .A(n124), .Y(n862) );
  ivd1_hd U134 ( .A(r_pstate[0]), .Y(N26) );
  ad2d1_hd U136 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(n808) );
  ivd1_hd U137 ( .A(n101), .Y(N556) );
  ivd1_hd U138 ( .A(r_pstate[1]), .Y(N25) );
  oa211d1_hd U139 ( .A(n545), .B(N26), .C(r_pstate[1]), .D(n554), .Y(n821) );
  oa211d1_hd U140 ( .A(n539), .B(N26), .C(n808), .D(N25), .Y(n820) );
  scg10d1_hd U142 ( .A(r_pstate[1]), .B(n822), .C(n554), .D(n823), .Y(n828) );
  ao21d1_hd U145 ( .A(n123), .B(n124), .C(n101), .Y(n865) );
  ivd1_hd U146 ( .A(r_x_data[63]), .Y(n824) );
  oa21d1_hd U147 ( .A(N563), .B(n539), .C(n826), .Y(n825) );
  ao22d1_hd U148 ( .A(n536), .B(r_x_data[62]), .C(n807), .D(o_Y_DATA[30]), .Y(
        n826) );
endmodule


module converter_f2i_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62;

  had1_hd U2 ( .A(n33), .B(n2), .CO(n1), .S(DIFF[30]) );
  had1_hd U3 ( .A(n34), .B(n3), .CO(n2), .S(DIFF[29]) );
  had1_hd U4 ( .A(n35), .B(n4), .CO(n3), .S(DIFF[28]) );
  had1_hd U5 ( .A(n36), .B(n5), .CO(n4), .S(DIFF[27]) );
  had1_hd U6 ( .A(n37), .B(n6), .CO(n5), .S(DIFF[26]) );
  had1_hd U7 ( .A(n38), .B(n7), .CO(n6), .S(DIFF[25]) );
  had1_hd U8 ( .A(n39), .B(n8), .CO(n7), .S(DIFF[24]) );
  had1_hd U9 ( .A(n40), .B(n9), .CO(n8), .S(DIFF[23]) );
  had1_hd U10 ( .A(n41), .B(n10), .CO(n9), .S(DIFF[22]) );
  had1_hd U11 ( .A(n42), .B(n11), .CO(n10), .S(DIFF[21]) );
  had1_hd U12 ( .A(n43), .B(n12), .CO(n11), .S(DIFF[20]) );
  had1_hd U13 ( .A(n44), .B(n13), .CO(n12), .S(DIFF[19]) );
  had1_hd U14 ( .A(n45), .B(n14), .CO(n13), .S(DIFF[18]) );
  had1_hd U15 ( .A(n46), .B(n15), .CO(n14), .S(DIFF[17]) );
  had1_hd U16 ( .A(n47), .B(n16), .CO(n15), .S(DIFF[16]) );
  had1_hd U17 ( .A(n48), .B(n17), .CO(n16), .S(DIFF[15]) );
  had1_hd U18 ( .A(n49), .B(n18), .CO(n17), .S(DIFF[14]) );
  had1_hd U19 ( .A(n50), .B(n19), .CO(n18), .S(DIFF[13]) );
  had1_hd U20 ( .A(n51), .B(n20), .CO(n19), .S(DIFF[12]) );
  had1_hd U21 ( .A(n52), .B(n21), .CO(n20), .S(DIFF[11]) );
  had1_hd U22 ( .A(n53), .B(n22), .CO(n21), .S(DIFF[10]) );
  had1_hd U23 ( .A(n54), .B(n23), .CO(n22), .S(DIFF[9]) );
  had1_hd U24 ( .A(n55), .B(n24), .CO(n23), .S(DIFF[8]) );
  had1_hd U25 ( .A(n56), .B(n25), .CO(n24), .S(DIFF[7]) );
  had1_hd U26 ( .A(n57), .B(n26), .CO(n25), .S(DIFF[6]) );
  had1_hd U27 ( .A(n58), .B(n27), .CO(n26), .S(DIFF[5]) );
  had1_hd U28 ( .A(n59), .B(n28), .CO(n27), .S(DIFF[4]) );
  had1_hd U29 ( .A(n60), .B(n29), .CO(n28), .S(DIFF[3]) );
  had1_hd U30 ( .A(n61), .B(n30), .CO(n29), .S(DIFF[2]) );
  had1_hd U31 ( .A(n62), .B(n31), .CO(n30), .S(DIFF[1]) );
  nid1_hd U68 ( .A(B[0]), .Y(DIFF[0]) );
  ivd1_hd U69 ( .A(B[1]), .Y(n62) );
  ivd1_hd U70 ( .A(B[2]), .Y(n61) );
  ivd1_hd U71 ( .A(B[3]), .Y(n60) );
  ivd1_hd U72 ( .A(B[4]), .Y(n59) );
  ivd1_hd U73 ( .A(B[5]), .Y(n58) );
  ivd1_hd U74 ( .A(B[6]), .Y(n57) );
  ivd1_hd U75 ( .A(B[7]), .Y(n56) );
  ivd1_hd U76 ( .A(B[8]), .Y(n55) );
  ivd1_hd U77 ( .A(B[9]), .Y(n54) );
  ivd1_hd U78 ( .A(B[10]), .Y(n53) );
  ivd1_hd U79 ( .A(B[11]), .Y(n52) );
  ivd1_hd U80 ( .A(B[12]), .Y(n51) );
  ivd1_hd U81 ( .A(B[13]), .Y(n50) );
  ivd1_hd U82 ( .A(B[14]), .Y(n49) );
  ivd1_hd U83 ( .A(B[15]), .Y(n48) );
  ivd1_hd U84 ( .A(B[16]), .Y(n47) );
  ivd1_hd U85 ( .A(B[17]), .Y(n46) );
  ivd1_hd U86 ( .A(B[18]), .Y(n45) );
  ivd1_hd U87 ( .A(B[19]), .Y(n44) );
  ivd1_hd U88 ( .A(B[20]), .Y(n43) );
  ivd1_hd U89 ( .A(B[21]), .Y(n42) );
  ivd1_hd U90 ( .A(B[22]), .Y(n41) );
  ivd1_hd U91 ( .A(B[23]), .Y(n40) );
  ivd1_hd U92 ( .A(B[24]), .Y(n39) );
  ivd1_hd U93 ( .A(B[25]), .Y(n38) );
  ivd1_hd U94 ( .A(B[26]), .Y(n37) );
  ivd1_hd U95 ( .A(B[27]), .Y(n36) );
  ivd1_hd U96 ( .A(B[28]), .Y(n35) );
  ivd1_hd U97 ( .A(B[29]), .Y(n34) );
  ivd1_hd U98 ( .A(B[30]), .Y(n33) );
  ivd1_hd U99 ( .A(B[0]), .Y(n31) );
  xn2d1_hd U100 ( .A(n1), .B(B[31]), .Y(DIFF[31]) );
endmodule


module converter_f2i_DP_OP_15_125_5858_0 ( I1, O1, U170_Y, i_CLK, IN0 );
  input [7:0] I1;
  output [8:0] O1;
  input U170_Y, i_CLK, IN0;
  wire   n2, n3, n4, n5, n6, n7, n29, n30, n1, n8, n9, n10, n11, n12, n13, n14
;

  had1_hd U4 ( .A(n13), .B(n3), .CO(n2), .S(O1[6]) );
  had1_hd U5 ( .A(n12), .B(n4), .CO(n3), .S(O1[5]) );
  had1_hd U6 ( .A(n11), .B(n5), .CO(n4), .S(O1[4]) );
  had1_hd U7 ( .A(n10), .B(n6), .CO(n5), .S(O1[3]) );
  had1_hd U8 ( .A(n9), .B(n7), .CO(n6), .S(O1[2]) );
  had1_hd U9 ( .A(n8), .B(n1), .CO(n7), .S(O1[1]) );
  nr2d1_hd U13 ( .A(n14), .B(n2), .Y(O1[8]) );
  ao22d1_hd U14 ( .A(n14), .B(n29), .C(n2), .D(n30), .Y(O1[7]) );
  ivd1_hd U15 ( .A(n14), .Y(n30) );
  ivd1_hd U16 ( .A(n2), .Y(n29) );
  ivd1_hd U17 ( .A(n1), .Y(O1[0]) );
  fd1qd1_hd clk_r_REG66_S1 ( .D(I1[7]), .CK(IN0), .Q(n14) );
  fd1qd1_hd clk_r_REG111_S1 ( .D(I1[6]), .CK(IN0), .Q(n13) );
  fd1qd1_hd clk_r_REG112_S1 ( .D(I1[5]), .CK(IN0), .Q(n12) );
  fd1qd1_hd clk_r_REG113_S1 ( .D(I1[4]), .CK(IN0), .Q(n11) );
  fd1qd1_hd clk_r_REG114_S1 ( .D(I1[3]), .CK(IN0), .Q(n10) );
  fd1qd1_hd clk_r_REG115_S1 ( .D(I1[2]), .CK(IN0), .Q(n9) );
  fd1qd1_hd clk_r_REG116_S1 ( .D(I1[1]), .CK(IN0), .Q(n8) );
  fd1qd1_hd clk_r_REG117_S1 ( .D(I1[0]), .CK(IN0), .Q(n1) );
endmodule


module converter_f2i_DP_OP_16_126_6114_0 ( I1, O1 );
  input [8:0] I1;
  output [8:0] O1;
  wire   n1, n2, n3, n4, n5, n6, n7;

  had1_hd U2 ( .A(I1[7]), .B(n2), .CO(n1), .S(O1[7]) );
  had1_hd U3 ( .A(I1[6]), .B(n3), .CO(n2), .S(O1[6]) );
  had1_hd U4 ( .A(I1[5]), .B(n4), .CO(n3), .S(O1[5]) );
  had1_hd U5 ( .A(I1[4]), .B(n5), .CO(n4), .S(O1[4]) );
  had1_hd U6 ( .A(I1[3]), .B(n6), .CO(n5), .S(O1[3]) );
  had1_hd U7 ( .A(I1[2]), .B(n7), .CO(n6), .S(O1[2]) );
  had1_hd U8 ( .A(I1[1]), .B(I1[0]), .CO(n7), .S(O1[1]) );
  xo2d1_hd U12 ( .A(I1[8]), .B(n1), .Y(O1[8]) );
  ivd1_hd U13 ( .A(I1[0]), .Y(O1[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_f2i_3_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_f2i_2_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_f2i_1_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_converter_f2i_0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module converter_f2i ( i_A, i_A_STB, o_A_ACK, o_Z, o_Z_STB, i_Z_ACK, i_CLK, 
        i_RST );
  input [31:0] i_A;
  output [31:0] o_Z;
  input i_A_STB, i_Z_ACK, i_CLK, i_RST;
  output o_A_ACK, o_Z_STB;
  wire   n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n195,
         n228, N17, N29, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N135, N139, N171, N181, n1, n2, n3,
         n4, n5, C1_DATA1_8, C1_DATA1_7, C1_DATA1_6, C1_DATA1_5, C1_DATA1_4,
         C1_DATA1_3, C1_DATA1_2, C1_DATA1_1, C1_DATA1_0, C1_DATA2_8,
         C1_DATA2_7, C1_DATA2_6, C1_DATA2_5, C1_DATA2_4, C1_DATA2_3,
         C1_DATA2_2, C1_DATA2_1, C1_DATA2_0, n21, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86,
         n88, n90, n92, n94, n96, n98, n100, n102, n104, n106, n108, n110,
         n112, n114, n116, n118, n120, n122, n124, n126, n128, n130, n132,
         n134, n136, n138, n140, n142, n144, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n159, n160, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n336;
  wire   [2:0] state;
  wire   [8:0] a_e;
  wire   [30:0] a_m;

  ivd1_hd U3 ( .A(i_RST), .Y(n1) );
  ivd1_hd U4 ( .A(i_RST), .Y(n2) );
  ivd1_hd U5 ( .A(i_RST), .Y(n3) );
  ivd1_hd U6 ( .A(i_RST), .Y(n4) );
  ivd1_hd U7 ( .A(i_RST), .Y(n5) );
  clknd2d1_hd U94 ( .A(n31), .B(n189), .Y(n25) );
  clknd2d1_hd U95 ( .A(n160), .B(n47), .Y(n36) );
  clknd2d1_hd U96 ( .A(n27), .B(n38), .Y(n40) );
  clknd2d1_hd U97 ( .A(n24), .B(n25), .Y(n196) );
  scg2d1_hd U98 ( .A(n26), .B(N93), .C(n29), .D(n147), .Y(n197) );
  scg2d1_hd U99 ( .A(n26), .B(N92), .C(n29), .D(n11), .Y(n198) );
  scg2d1_hd U100 ( .A(n26), .B(N91), .C(n29), .D(n12), .Y(n199) );
  scg2d1_hd U101 ( .A(n26), .B(N90), .C(n29), .D(n13), .Y(n200) );
  scg2d1_hd U102 ( .A(n26), .B(N89), .C(n29), .D(n14), .Y(n201) );
  scg2d1_hd U103 ( .A(n26), .B(N88), .C(n29), .D(n15), .Y(n202) );
  scg2d1_hd U104 ( .A(n26), .B(N63), .C(n29), .D(n149), .Y(n227) );
  scg2d1_hd U105 ( .A(n26), .B(N64), .C(n29), .D(n150), .Y(n226) );
  scg2d1_hd U106 ( .A(n26), .B(N65), .C(n29), .D(n151), .Y(n225) );
  scg2d1_hd U107 ( .A(n26), .B(N66), .C(n29), .D(n152), .Y(n224) );
  scg2d1_hd U108 ( .A(n26), .B(N67), .C(n29), .D(n153), .Y(n223) );
  scg2d1_hd U109 ( .A(n26), .B(N68), .C(n29), .D(n154), .Y(n222) );
  scg2d1_hd U110 ( .A(n26), .B(N69), .C(n29), .D(n155), .Y(n221) );
  scg2d1_hd U111 ( .A(n26), .B(N70), .C(n29), .D(n156), .Y(n220) );
  scg2d1_hd U112 ( .A(n26), .B(N71), .C(n29), .D(n75), .Y(n219) );
  scg2d1_hd U113 ( .A(n26), .B(N72), .C(n29), .D(n74), .Y(n218) );
  scg2d1_hd U114 ( .A(n26), .B(N73), .C(n29), .D(n73), .Y(n217) );
  scg2d1_hd U115 ( .A(n26), .B(N74), .C(n29), .D(n72), .Y(n216) );
  scg2d1_hd U116 ( .A(n26), .B(N75), .C(n29), .D(n71), .Y(n215) );
  scg2d1_hd U117 ( .A(n26), .B(N76), .C(n29), .D(n70), .Y(n214) );
  scg2d1_hd U118 ( .A(n26), .B(N77), .C(n29), .D(n69), .Y(n213) );
  scg2d1_hd U119 ( .A(n26), .B(N78), .C(n29), .D(n68), .Y(n212) );
  scg2d1_hd U120 ( .A(n26), .B(N79), .C(n29), .D(n67), .Y(n211) );
  scg2d1_hd U121 ( .A(n26), .B(N80), .C(n29), .D(n66), .Y(n210) );
  scg2d1_hd U122 ( .A(n26), .B(N81), .C(n29), .D(n65), .Y(n209) );
  scg2d1_hd U123 ( .A(n26), .B(N82), .C(n29), .D(n64), .Y(n208) );
  scg2d1_hd U124 ( .A(n26), .B(N83), .C(n29), .D(n20), .Y(n207) );
  scg2d1_hd U125 ( .A(n26), .B(N84), .C(n29), .D(n19), .Y(n206) );
  scg2d1_hd U126 ( .A(n26), .B(N85), .C(n29), .D(n18), .Y(n205) );
  scg2d1_hd U127 ( .A(n26), .B(N86), .C(n29), .D(n17), .Y(n204) );
  scg2d1_hd U128 ( .A(n26), .B(N87), .C(n29), .D(n16), .Y(n203) );
  scg2d1_hd U129 ( .A(n31), .B(C1_DATA2_0), .C(n186), .D(C1_DATA1_0), .Y(
        a_e[0]) );
  scg2d1_hd U130 ( .A(n31), .B(C1_DATA2_1), .C(n186), .D(C1_DATA1_1), .Y(
        a_e[1]) );
  scg2d1_hd U131 ( .A(n31), .B(C1_DATA2_2), .C(n186), .D(C1_DATA1_2), .Y(
        a_e[2]) );
  scg2d1_hd U132 ( .A(n31), .B(C1_DATA2_3), .C(n186), .D(C1_DATA1_3), .Y(
        a_e[3]) );
  scg2d1_hd U133 ( .A(n31), .B(C1_DATA2_4), .C(n186), .D(C1_DATA1_4), .Y(
        a_e[4]) );
  scg2d1_hd U134 ( .A(n31), .B(C1_DATA2_5), .C(n186), .D(C1_DATA1_5), .Y(
        a_e[5]) );
  scg2d1_hd U135 ( .A(n31), .B(C1_DATA2_6), .C(n186), .D(C1_DATA1_6), .Y(
        a_e[6]) );
  scg2d1_hd U136 ( .A(n31), .B(C1_DATA2_7), .C(n186), .D(C1_DATA1_7), .Y(
        a_e[7]) );
  scg2d1_hd U137 ( .A(n31), .B(C1_DATA2_8), .C(n186), .D(C1_DATA1_8), .Y(
        a_e[8]) );
  clknd2d1_hd U160 ( .A(n39), .B(n40), .Y(state[1]) );
  clknd2d1_hd U161 ( .A(n37), .B(n33), .Y(state[2]) );
  clknd2d1_hd U162 ( .A(i_Z_ACK), .B(o_Z_STB), .Y(n228) );
  or2d1_hd U163 ( .A(n148), .B(n36), .Y(n21) );
  ad2bd2_hd U164 ( .B(n187), .AN(n30), .Y(n26) );
  nr2d4_hd U168 ( .A(n187), .B(n30), .Y(n29) );
  clknd2d1_hd U169 ( .A(n148), .B(n47), .Y(n63) );
  clknd2d1_hd U171 ( .A(i_A_STB), .B(o_A_ACK), .Y(n195) );
  clknd2d1_hd U173 ( .A(n62), .B(n34), .Y(n48) );
  ao22d1_hd U175 ( .A(n26), .B(N94), .C(n27), .D(n28), .Y(n24) );
  nd2bd1_hd U176 ( .AN(n189), .B(n31), .Y(n30) );
  scg14d1_hd U177 ( .A(n186), .B(n185), .C(n25), .Y(a_m[30]) );
  nr2bd1_hd U180 ( .AN(n155), .B(n37), .Y(a_m[5]) );
  nr2bd1_hd U181 ( .AN(n154), .B(n37), .Y(a_m[4]) );
  nr2bd1_hd U182 ( .AN(n153), .B(n37), .Y(a_m[3]) );
  nr2bd1_hd U183 ( .AN(n152), .B(n37), .Y(a_m[2]) );
  nr2bd1_hd U184 ( .AN(n151), .B(n37), .Y(a_m[1]) );
  nr2bd1_hd U185 ( .AN(n150), .B(n37), .Y(a_m[0]) );
  nd2bd1_hd U186 ( .AN(n38), .B(n27), .Y(n33) );
  nd2bd1_hd U187 ( .AN(n186), .B(n40), .Y(state[0]) );
  nr2bd1_hd U188 ( .AN(n41), .B(n28), .Y(n38) );
  ao21d1_hd U189 ( .A(n42), .B(n43), .C(n76), .Y(n28) );
  nd4d1_hd U190 ( .A(n42), .B(n84), .C(n44), .D(n45), .Y(n41) );
  nr4d1_hd U191 ( .A(n82), .B(n81), .C(n83), .D(n43), .Y(n44) );
  scg16d1_hd U192 ( .A(N29), .B(n228), .C(n46), .Y(N135) );
  nr4d1_hd U193 ( .A(n27), .B(n32), .C(N139), .D(n186), .Y(n46) );
  ivd1_hd U194 ( .A(N17), .Y(n39) );
  nr2d1_hd U195 ( .A(n159), .B(n48), .Y(N17) );
  nr2d1_hd U196 ( .A(n37), .B(n35), .Y(n32) );
  scg10d1_hd U197 ( .A(n49), .B(n50), .C(n51), .D(n76), .Y(n35) );
  ao211d1_hd U198 ( .A(n52), .B(n81), .C(n53), .D(n77), .Y(n51) );
  ivd1_hd U199 ( .A(n42), .Y(n53) );
  nr2d1_hd U200 ( .A(n79), .B(n78), .Y(n42) );
  ad4d1_hd U201 ( .A(n82), .B(n83), .C(n80), .D(n84), .Y(n52) );
  nd4d1_hd U202 ( .A(n54), .B(n55), .C(n56), .D(n57), .Y(n50) );
  nr4d1_hd U203 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(n57) );
  nr4d1_hd U204 ( .A(n64), .B(n65), .C(n66), .D(n67), .Y(n56) );
  nr4d1_hd U205 ( .A(n147), .B(n11), .C(n12), .D(n149), .Y(n55) );
  nr4d1_hd U206 ( .A(n13), .B(n14), .C(n15), .D(n16), .Y(n54) );
  nd4d1_hd U207 ( .A(n58), .B(n59), .C(n60), .D(n61), .Y(n49) );
  nr4d1_hd U208 ( .A(n156), .B(n155), .C(n154), .D(n153), .Y(n61) );
  nr4d1_hd U209 ( .A(n189), .B(n152), .C(n151), .D(n150), .Y(n60) );
  nr4d1_hd U210 ( .A(n68), .B(n69), .C(n70), .D(n71), .Y(n59) );
  nr4d1_hd U211 ( .A(n72), .B(n73), .C(n74), .D(n75), .Y(n58) );
  ivd1_hd U212 ( .A(n31), .Y(n37) );
  nr2d1_hd U213 ( .A(n160), .B(n63), .Y(n27) );
  ivd1_hd U214 ( .A(n148), .Y(n34) );
  ivd1_hd U215 ( .A(n160), .Y(n62) );
  ivd1_hd U216 ( .A(n159), .Y(n47) );
  ivd1_hd U1 ( .A(i_RST), .Y(n6) );
  ivd1_hd U2 ( .A(i_RST), .Y(n7) );
  ivd1_hd U8 ( .A(i_RST), .Y(n8) );
  ivd1_hd U9 ( .A(i_RST), .Y(n9) );
  ivd1_hd U10 ( .A(i_RST), .Y(n10) );
  ivd6_hd U14 ( .A(n5) );
  ivd6_hd U15 ( .A(n1) );
  ivd6_hd U16 ( .A(n4) );
  ivd6_hd U17 ( .A(n2) );
  ivd6_hd U18 ( .A(n3) );
  fds2eqd1_hd clk_r_REG107_S3 ( .CRN(n6), .D(state[0]), .E(N135), .CK(i_CLK), 
        .Q(n148) );
  fds2eqd1_hd clk_r_REG69_S3 ( .CRN(n9), .D(state[2]), .E(N135), .CK(i_CLK), 
        .Q(n159) );
  fds2eqd1_hd clk_r_REG68_S3 ( .CRN(n10), .D(state[1]), .E(N135), .CK(i_CLK), 
        .Q(n160) );
  fd1eqd1_hd clk_r_REG1_S2 ( .D(n188), .E(n186), .CK(n230), .Q(n187) );
  fd1eqd1_hd clk_r_REG109_S4 ( .D(a_e[1]), .E(N171), .CK(i_CLK), .Q(n83) );
  fd1eqd1_hd clk_r_REG108_S4 ( .D(a_e[0]), .E(N171), .CK(i_CLK), .Q(n84) );
  fd1eqd1_hd clk_r_REG72_S5 ( .D(a_e[4]), .E(N171), .CK(i_CLK), .Q(n80) );
  fd1eqd1_hd clk_r_REG71_S4 ( .D(a_e[3]), .E(N171), .CK(i_CLK), .Q(n81) );
  fd1eqd1_hd clk_r_REG70_S4 ( .D(a_e[2]), .E(N171), .CK(i_CLK), .Q(n82) );
  fd1eqd1_hd clk_r_REG75_S5 ( .D(a_e[7]), .E(N171), .CK(i_CLK), .Q(n77) );
  fd1eqd1_hd clk_r_REG67_S2 ( .D(a_e[8]), .E(N171), .CK(i_CLK), .Q(n76) );
  ivd1_hd U11 ( .A(n77), .Y(n43) );
  ivd1_hd U12 ( .A(n80), .Y(n45) );
  ivd2_hd U20 ( .A(n21), .Y(n186) );
  fd1qd1_hd clk_r_REG79_S7 ( .D(a_m[5]), .CK(n230), .Q(n154) );
  fd1qd1_hd clk_r_REG80_S8 ( .D(a_m[4]), .CK(n230), .Q(n153) );
  fd1qd1_hd clk_r_REG81_S9 ( .D(a_m[3]), .CK(n230), .Q(n152) );
  fd1qd1_hd clk_r_REG82_S10 ( .D(a_m[2]), .CK(n230), .Q(n151) );
  fd1qd1_hd clk_r_REG83_S11 ( .D(a_m[1]), .CK(n230), .Q(n150) );
  fd1qd1_hd clk_r_REG84_S12 ( .D(a_m[0]), .CK(n230), .Q(n149) );
  fd1qd1_hd clk_r_REG76_S4 ( .D(n332), .CK(n230), .Q(n75) );
  fd1qd1_hd clk_r_REG77_S5 ( .D(n331), .CK(n230), .Q(n156) );
  fd1qd1_hd clk_r_REG78_S6 ( .D(n330), .CK(n230), .Q(n155) );
  fd1qd1_hd clk_r_REG85_S4 ( .D(n329), .CK(n230), .Q(n72) );
  fd1qd1_hd clk_r_REG86_S5 ( .D(n328), .CK(n230), .Q(n73) );
  fd1qd1_hd clk_r_REG87_S6 ( .D(n327), .CK(n230), .Q(n74) );
  fd1qd1_hd clk_r_REG88_S4 ( .D(n326), .CK(n230), .Q(n69) );
  fd1qd1_hd clk_r_REG89_S5 ( .D(n325), .CK(n230), .Q(n70) );
  fd1qd1_hd clk_r_REG90_S6 ( .D(n324), .CK(n230), .Q(n71) );
  fd1qd1_hd clk_r_REG91_S4 ( .D(n323), .CK(n230), .Q(n66) );
  fd1qd1_hd clk_r_REG92_S5 ( .D(n322), .CK(n230), .Q(n67) );
  fd1qd1_hd clk_r_REG93_S6 ( .D(n321), .CK(n230), .Q(n68) );
  fd1qd1_hd clk_r_REG94_S4 ( .D(n320), .CK(n230), .Q(n20) );
  fd1qd1_hd clk_r_REG95_S5 ( .D(n319), .CK(n230), .Q(n64) );
  fd1qd1_hd clk_r_REG96_S6 ( .D(n318), .CK(n230), .Q(n65) );
  fd1qd1_hd clk_r_REG97_S4 ( .D(n317), .CK(n230), .Q(n17) );
  fd1qd1_hd clk_r_REG98_S5 ( .D(n316), .CK(n230), .Q(n18) );
  fd1qd1_hd clk_r_REG99_S6 ( .D(n315), .CK(n230), .Q(n19) );
  fd1qd1_hd clk_r_REG100_S4 ( .D(n314), .CK(n230), .Q(n14) );
  fd1qd1_hd clk_r_REG101_S5 ( .D(n313), .CK(n230), .Q(n15) );
  fd1qd1_hd clk_r_REG102_S6 ( .D(n312), .CK(n230), .Q(n16) );
  fd1qd1_hd clk_r_REG103_S4 ( .D(n311), .CK(n230), .Q(n11) );
  fd1qd1_hd clk_r_REG104_S5 ( .D(n310), .CK(n230), .Q(n12) );
  fd1qd1_hd clk_r_REG105_S6 ( .D(n309), .CK(n230), .Q(n13) );
  fd1qd1_hd clk_r_REG106_S4 ( .D(a_m[30]), .CK(n230), .Q(n147) );
  fd1qd1_hd clk_r_REG110_S4 ( .D(n34), .CK(n230), .Q(n189) );
  fd1qd1_hd clk_r_REG64_S3 ( .D(n196), .CK(n231), .Q(n162) );
  fd1qd1_hd clk_r_REG2_S3 ( .D(n197), .CK(n231), .Q(n146) );
  fd1qd1_hd clk_r_REG4_S3 ( .D(n198), .CK(n231), .Q(n144) );
  fd1qd1_hd clk_r_REG6_S3 ( .D(n199), .CK(n231), .Q(n142) );
  fd1qd1_hd clk_r_REG8_S3 ( .D(n200), .CK(n231), .Q(n140) );
  fd1qd1_hd clk_r_REG10_S3 ( .D(n201), .CK(n231), .Q(n138) );
  fd1qd1_hd clk_r_REG12_S3 ( .D(n202), .CK(n231), .Q(n136) );
  fd1qd1_hd clk_r_REG62_S3 ( .D(n203), .CK(n231), .Q(n86) );
  fd1qd1_hd clk_r_REG60_S3 ( .D(n204), .CK(n231), .Q(n88) );
  fd1qd1_hd clk_r_REG58_S3 ( .D(n205), .CK(n231), .Q(n90) );
  fd1qd1_hd clk_r_REG56_S3 ( .D(n206), .CK(n231), .Q(n92) );
  fd1qd1_hd clk_r_REG54_S3 ( .D(n207), .CK(n231), .Q(n94) );
  fd1qd1_hd clk_r_REG52_S3 ( .D(n208), .CK(n231), .Q(n96) );
  fd1qd1_hd clk_r_REG50_S3 ( .D(n209), .CK(n231), .Q(n98) );
  fd1qd1_hd clk_r_REG48_S3 ( .D(n210), .CK(n231), .Q(n100) );
  fd1qd1_hd clk_r_REG46_S3 ( .D(n211), .CK(n231), .Q(n102) );
  fd1qd1_hd clk_r_REG44_S3 ( .D(n212), .CK(n231), .Q(n104) );
  fd1qd1_hd clk_r_REG42_S3 ( .D(n213), .CK(n231), .Q(n106) );
  fd1qd1_hd clk_r_REG40_S3 ( .D(n214), .CK(n231), .Q(n108) );
  fd1qd1_hd clk_r_REG38_S3 ( .D(n215), .CK(n231), .Q(n110) );
  fd1qd1_hd clk_r_REG14_S3 ( .D(n227), .CK(n231), .Q(n134) );
  fd1qd1_hd clk_r_REG16_S3 ( .D(n226), .CK(n231), .Q(n132) );
  fd1qd1_hd clk_r_REG18_S3 ( .D(n225), .CK(n231), .Q(n130) );
  fd1qd1_hd clk_r_REG20_S3 ( .D(n224), .CK(n231), .Q(n128) );
  fd1qd1_hd clk_r_REG22_S3 ( .D(n223), .CK(n231), .Q(n126) );
  fd1qd1_hd clk_r_REG24_S3 ( .D(n222), .CK(n231), .Q(n124) );
  fd1qd1_hd clk_r_REG26_S3 ( .D(n221), .CK(n231), .Q(n122) );
  fd1qd1_hd clk_r_REG28_S3 ( .D(n220), .CK(n231), .Q(n120) );
  fd1qd1_hd clk_r_REG30_S3 ( .D(n219), .CK(n231), .Q(n118) );
  fd1qd1_hd clk_r_REG32_S3 ( .D(n218), .CK(n231), .Q(n116) );
  fd1qd1_hd clk_r_REG34_S3 ( .D(n217), .CK(n231), .Q(n114) );
  fd1qd1_hd clk_r_REG36_S3 ( .D(n216), .CK(n231), .Q(n112) );
  fd1qd1_hd clk_r_REG3_S4 ( .D(n146), .CK(n232), .Q(o_Z[30]) );
  fd1qd1_hd clk_r_REG5_S4 ( .D(n144), .CK(n232), .Q(o_Z[29]) );
  fd1qd1_hd clk_r_REG7_S4 ( .D(n142), .CK(n232), .Q(o_Z[28]) );
  fd1qd1_hd clk_r_REG9_S4 ( .D(n140), .CK(n232), .Q(o_Z[27]) );
  fd1qd1_hd clk_r_REG11_S4 ( .D(n138), .CK(n232), .Q(o_Z[26]) );
  fd1qd1_hd clk_r_REG13_S4 ( .D(n136), .CK(n232), .Q(o_Z[25]) );
  fd1qd1_hd clk_r_REG15_S4 ( .D(n134), .CK(n232), .Q(o_Z[0]) );
  fd1qd1_hd clk_r_REG17_S4 ( .D(n132), .CK(n232), .Q(o_Z[1]) );
  fd1qd1_hd clk_r_REG19_S4 ( .D(n130), .CK(n232), .Q(o_Z[2]) );
  fd1qd1_hd clk_r_REG21_S4 ( .D(n128), .CK(n232), .Q(o_Z[3]) );
  fd1qd1_hd clk_r_REG23_S4 ( .D(n126), .CK(n232), .Q(o_Z[4]) );
  fd1qd1_hd clk_r_REG25_S4 ( .D(n124), .CK(n232), .Q(o_Z[5]) );
  fd1qd1_hd clk_r_REG27_S4 ( .D(n122), .CK(n232), .Q(o_Z[6]) );
  fd1qd1_hd clk_r_REG29_S4 ( .D(n120), .CK(n232), .Q(o_Z[7]) );
  fd1qd1_hd clk_r_REG31_S4 ( .D(n118), .CK(n232), .Q(o_Z[8]) );
  fd1qd1_hd clk_r_REG33_S4 ( .D(n116), .CK(n232), .Q(o_Z[9]) );
  fd1qd1_hd clk_r_REG35_S4 ( .D(n114), .CK(n232), .Q(o_Z[10]) );
  fd1qd1_hd clk_r_REG37_S4 ( .D(n112), .CK(n232), .Q(o_Z[11]) );
  fd1qd1_hd clk_r_REG39_S4 ( .D(n110), .CK(n232), .Q(o_Z[12]) );
  fd1qd1_hd clk_r_REG41_S4 ( .D(n108), .CK(n232), .Q(o_Z[13]) );
  fd1qd1_hd clk_r_REG43_S4 ( .D(n106), .CK(n232), .Q(o_Z[14]) );
  fd1qd1_hd clk_r_REG45_S4 ( .D(n104), .CK(n232), .Q(o_Z[15]) );
  fd1qd1_hd clk_r_REG47_S4 ( .D(n102), .CK(n232), .Q(o_Z[16]) );
  fd1qd1_hd clk_r_REG49_S4 ( .D(n100), .CK(n232), .Q(o_Z[17]) );
  fd1qd1_hd clk_r_REG51_S4 ( .D(n98), .CK(n232), .Q(o_Z[18]) );
  fd1qd1_hd clk_r_REG53_S4 ( .D(n96), .CK(n232), .Q(o_Z[19]) );
  fd1qd1_hd clk_r_REG55_S4 ( .D(n94), .CK(n232), .Q(o_Z[20]) );
  fd1qd1_hd clk_r_REG57_S4 ( .D(n92), .CK(n232), .Q(o_Z[21]) );
  fd1qd1_hd clk_r_REG59_S4 ( .D(n90), .CK(n232), .Q(o_Z[22]) );
  fd1qd1_hd clk_r_REG61_S4 ( .D(n88), .CK(n232), .Q(o_Z[23]) );
  fd1qd1_hd clk_r_REG63_S4 ( .D(n86), .CK(n232), .Q(o_Z[24]) );
  fd1qd1_hd clk_r_REG65_S4 ( .D(n162), .CK(n232), .Q(o_Z[31]) );
  fd1qd1_hd clk_r_REG0_S1 ( .D(i_A[31]), .CK(n233), .Q(n188) );
  fd1qd1_hd clk_r_REG118_S1 ( .D(i_A[22]), .CK(n233), .Q(n185) );
  fd1qd1_hd clk_r_REG119_S1 ( .D(i_A[21]), .CK(n233), .Q(n184) );
  fd1qd1_hd clk_r_REG120_S1 ( .D(i_A[20]), .CK(n233), .Q(n183) );
  fd1qd1_hd clk_r_REG121_S1 ( .D(i_A[19]), .CK(n233), .Q(n182) );
  fd1qd1_hd clk_r_REG122_S1 ( .D(i_A[18]), .CK(n233), .Q(n181) );
  fd1qd1_hd clk_r_REG123_S1 ( .D(i_A[17]), .CK(n233), .Q(n180) );
  fd1qd1_hd clk_r_REG124_S1 ( .D(i_A[16]), .CK(n233), .Q(n179) );
  fd1qd1_hd clk_r_REG125_S1 ( .D(i_A[15]), .CK(n233), .Q(n178) );
  fd1qd1_hd clk_r_REG126_S1 ( .D(i_A[14]), .CK(n233), .Q(n177) );
  fd1qd1_hd clk_r_REG127_S1 ( .D(i_A[13]), .CK(n233), .Q(n176) );
  fd1qd1_hd clk_r_REG128_S1 ( .D(i_A[12]), .CK(n233), .Q(n175) );
  fd1qd1_hd clk_r_REG129_S1 ( .D(i_A[11]), .CK(n233), .Q(n174) );
  fd1qd1_hd clk_r_REG130_S1 ( .D(i_A[10]), .CK(n233), .Q(n173) );
  fd1qd1_hd clk_r_REG131_S1 ( .D(i_A[9]), .CK(n233), .Q(n172) );
  fd1qd1_hd clk_r_REG132_S1 ( .D(i_A[8]), .CK(n233), .Q(n171) );
  fd1qd1_hd clk_r_REG133_S1 ( .D(i_A[7]), .CK(n233), .Q(n170) );
  fd1qd1_hd clk_r_REG134_S1 ( .D(i_A[6]), .CK(n233), .Q(n169) );
  fd1qd1_hd clk_r_REG135_S1 ( .D(i_A[5]), .CK(n233), .Q(n168) );
  fd1qd1_hd clk_r_REG136_S1 ( .D(i_A[4]), .CK(n233), .Q(n167) );
  fd1qd1_hd clk_r_REG137_S1 ( .D(i_A[3]), .CK(n233), .Q(n166) );
  fd1qd1_hd clk_r_REG138_S1 ( .D(i_A[2]), .CK(n233), .Q(n165) );
  fd1qd1_hd clk_r_REG139_S1 ( .D(i_A[1]), .CK(n233), .Q(n164) );
  fd1qd1_hd clk_r_REG140_S1 ( .D(i_A[0]), .CK(n233), .Q(n163) );
  fd1eqd1_hd clk_r_REG141_S1 ( .D(n236), .E(n303), .CK(i_CLK), .Q(o_A_ACK) );
  fd1eqd1_hd clk_r_REG142_S1 ( .D(n234), .E(n305), .CK(i_CLK), .Q(o_Z_STB) );
  fd1eqd1_hd clk_r_REG74_S4 ( .D(a_e[6]), .E(N171), .CK(n230), .Q(n78) );
  fd1eqd1_hd clk_r_REG73_S4 ( .D(a_e[5]), .E(N171), .CK(n230), .Q(n79) );
  converter_f2i_DW01_sub_0 sub_x_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({n189, n147, n11, n12, n13, n14, n15, n16, n17, n18, 
        n19, n20, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
        n156, n155, n154, n153, n152, n151, n150, n149}), .CI(1'b0), .DIFF({
        N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, 
        N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        N66, N65, N64, N63}) );
  converter_f2i_DP_OP_15_125_5858_0 DP_OP_15_125_5858 ( .I1(i_A[30:23]), .O1({
        C1_DATA1_8, C1_DATA1_7, C1_DATA1_6, C1_DATA1_5, C1_DATA1_4, C1_DATA1_3, 
        C1_DATA1_2, C1_DATA1_1, C1_DATA1_0}), .U170_Y(1'b0), .i_CLK(i_CLK), 
        .IN0(n233) );
  converter_f2i_DP_OP_16_126_6114_0 DP_OP_16_126_6114 ( .I1({n76, n77, n78, 
        n79, n80, n81, n82, n83, n84}), .O1({C1_DATA2_8, C1_DATA2_7, 
        C1_DATA2_6, C1_DATA2_5, C1_DATA2_4, C1_DATA2_3, C1_DATA2_2, C1_DATA2_1, 
        C1_DATA2_0}) );
  SNPS_CLOCK_GATE_HIGH_converter_f2i_3_0 clk_gate_clk_r_REG66_S1 ( .CLK(i_CLK), 
        .EN(N139), .ENCLK(n233), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_f2i_2_0 clk_gate_clk_r_REG3_S4_0 ( .CLK(i_CLK), .EN(N29), .ENCLK(n232), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_f2i_1_0 clk_gate_clk_r_REG64_S3_0 ( .CLK(
        i_CLK), .EN(N181), .ENCLK(n231), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_converter_f2i_0_0 clk_gate_clk_r_REG73_S4_0 ( .CLK(
        i_CLK), .EN(n336), .ENCLK(n230), .TE(1'b0) );
  ad2bd1_hd U13 ( .B(n160), .AN(n63), .Y(n31) );
  nd2bd1_hd U19 ( .AN(n32), .B(n33), .Y(N181) );
  nr2d1_hd U21 ( .A(n47), .B(n48), .Y(N29) );
  nr2d1_hd U22 ( .A(n195), .B(n39), .Y(N139) );
  ivd1_hd U23 ( .A(n235), .Y(n234) );
  clknd2d1_hd U24 ( .A(n8), .B(n304), .Y(n235) );
  ivd1_hd U25 ( .A(n237), .Y(n236) );
  clknd2d1_hd U26 ( .A(n7), .B(n302), .Y(n237) );
  scg2d1_hd U27 ( .A(n186), .B(n163), .C(n74), .D(n334), .Y(n332) );
  scg20d2_hd U28 ( .A(n34), .B(n35), .C(n36), .Y(N171) );
  or2d2_hd U29 ( .A(n186), .B(n334), .Y(n333) );
  ivd2_hd U30 ( .A(n63), .Y(n334) );
  ad2d1_hd U32 ( .A(n195), .B(n7), .Y(n302) );
  nd2bd1_hd U33 ( .AN(N17), .B(n7), .Y(n303) );
  ad2d1_hd U34 ( .A(n228), .B(n8), .Y(n304) );
  nd2bd1_hd U35 ( .AN(N29), .B(n8), .Y(n305) );
  ao21d1_hd U36 ( .A(n182), .B(n238), .C(n239), .Y(n309) );
  ao21d1_hd U37 ( .A(n12), .B(n334), .C(n182), .Y(n239) );
  ao22d1_hd U38 ( .A(n12), .B(n333), .C(n186), .D(n240), .Y(n238) );
  ivd1_hd U39 ( .A(n12), .Y(n240) );
  ao21d1_hd U40 ( .A(n183), .B(n241), .C(n242), .Y(n310) );
  ao21d1_hd U41 ( .A(n11), .B(n334), .C(n183), .Y(n242) );
  ao22d1_hd U42 ( .A(n11), .B(n333), .C(n186), .D(n243), .Y(n241) );
  ivd1_hd U43 ( .A(n11), .Y(n243) );
  ao21d1_hd U44 ( .A(n184), .B(n244), .C(n245), .Y(n311) );
  ao21d1_hd U45 ( .A(n147), .B(n334), .C(n184), .Y(n245) );
  ao22d1_hd U46 ( .A(n147), .B(n333), .C(n186), .D(n246), .Y(n244) );
  ivd1_hd U47 ( .A(n147), .Y(n246) );
  ao21d1_hd U48 ( .A(n179), .B(n247), .C(n248), .Y(n312) );
  ao21d1_hd U49 ( .A(n15), .B(n334), .C(n179), .Y(n248) );
  ao22d1_hd U50 ( .A(n15), .B(n333), .C(n186), .D(n249), .Y(n247) );
  ivd1_hd U51 ( .A(n15), .Y(n249) );
  ao21d1_hd U52 ( .A(n180), .B(n250), .C(n251), .Y(n313) );
  ao21d1_hd U53 ( .A(n14), .B(n334), .C(n180), .Y(n251) );
  ao22d1_hd U54 ( .A(n14), .B(n333), .C(n186), .D(n252), .Y(n250) );
  ivd1_hd U55 ( .A(n14), .Y(n252) );
  ao21d1_hd U56 ( .A(n181), .B(n253), .C(n254), .Y(n314) );
  ao21d1_hd U57 ( .A(n13), .B(n334), .C(n181), .Y(n254) );
  ao22d1_hd U58 ( .A(n13), .B(n333), .C(n186), .D(n255), .Y(n253) );
  ivd1_hd U59 ( .A(n13), .Y(n255) );
  ao21d1_hd U60 ( .A(n176), .B(n256), .C(n257), .Y(n315) );
  ao21d1_hd U61 ( .A(n18), .B(n334), .C(n176), .Y(n257) );
  ao22d1_hd U62 ( .A(n18), .B(n333), .C(n186), .D(n258), .Y(n256) );
  ivd1_hd U63 ( .A(n18), .Y(n258) );
  ao21d1_hd U64 ( .A(n177), .B(n259), .C(n260), .Y(n316) );
  ao21d1_hd U65 ( .A(n17), .B(n334), .C(n177), .Y(n260) );
  ao22d1_hd U66 ( .A(n17), .B(n333), .C(n186), .D(n261), .Y(n259) );
  ivd1_hd U67 ( .A(n17), .Y(n261) );
  ao21d1_hd U68 ( .A(n178), .B(n262), .C(n263), .Y(n317) );
  ao21d1_hd U69 ( .A(n16), .B(n334), .C(n178), .Y(n263) );
  ao22d1_hd U70 ( .A(n16), .B(n333), .C(n186), .D(n264), .Y(n262) );
  ivd1_hd U71 ( .A(n16), .Y(n264) );
  ao21d1_hd U72 ( .A(n173), .B(n265), .C(n266), .Y(n318) );
  ao21d1_hd U73 ( .A(n64), .B(n334), .C(n173), .Y(n266) );
  ao22d1_hd U74 ( .A(n64), .B(n333), .C(n186), .D(n267), .Y(n265) );
  ivd1_hd U75 ( .A(n64), .Y(n267) );
  ao21d1_hd U76 ( .A(n174), .B(n268), .C(n269), .Y(n319) );
  ao21d1_hd U77 ( .A(n20), .B(n334), .C(n174), .Y(n269) );
  ao22d1_hd U78 ( .A(n20), .B(n333), .C(n186), .D(n270), .Y(n268) );
  ivd1_hd U79 ( .A(n20), .Y(n270) );
  ao21d1_hd U80 ( .A(n175), .B(n271), .C(n272), .Y(n320) );
  ao21d1_hd U81 ( .A(n19), .B(n334), .C(n175), .Y(n272) );
  ao22d1_hd U82 ( .A(n19), .B(n333), .C(n186), .D(n273), .Y(n271) );
  ivd1_hd U83 ( .A(n19), .Y(n273) );
  ao21d1_hd U84 ( .A(n170), .B(n274), .C(n275), .Y(n321) );
  ao21d1_hd U85 ( .A(n67), .B(n334), .C(n170), .Y(n275) );
  ao22d1_hd U86 ( .A(n67), .B(n333), .C(n186), .D(n276), .Y(n274) );
  ivd1_hd U87 ( .A(n67), .Y(n276) );
  ao21d1_hd U88 ( .A(n171), .B(n277), .C(n278), .Y(n322) );
  ao21d1_hd U89 ( .A(n66), .B(n334), .C(n171), .Y(n278) );
  ao22d1_hd U90 ( .A(n66), .B(n333), .C(n186), .D(n279), .Y(n277) );
  ivd1_hd U91 ( .A(n66), .Y(n279) );
  ao21d1_hd U92 ( .A(n172), .B(n280), .C(n281), .Y(n323) );
  ao21d1_hd U93 ( .A(n65), .B(n334), .C(n172), .Y(n281) );
  ao22d1_hd U138 ( .A(n65), .B(n333), .C(n186), .D(n282), .Y(n280) );
  ivd1_hd U139 ( .A(n65), .Y(n282) );
  ao21d1_hd U140 ( .A(n167), .B(n283), .C(n284), .Y(n324) );
  ao21d1_hd U141 ( .A(n70), .B(n334), .C(n167), .Y(n284) );
  ao22d1_hd U142 ( .A(n70), .B(n333), .C(n186), .D(n285), .Y(n283) );
  ivd1_hd U143 ( .A(n70), .Y(n285) );
  ao21d1_hd U144 ( .A(n168), .B(n286), .C(n287), .Y(n325) );
  ao21d1_hd U145 ( .A(n69), .B(n334), .C(n168), .Y(n287) );
  ao22d1_hd U146 ( .A(n69), .B(n333), .C(n186), .D(n288), .Y(n286) );
  ivd1_hd U147 ( .A(n69), .Y(n288) );
  ao21d1_hd U148 ( .A(n169), .B(n289), .C(n290), .Y(n326) );
  ao21d1_hd U149 ( .A(n68), .B(n334), .C(n169), .Y(n290) );
  ao22d1_hd U150 ( .A(n68), .B(n333), .C(n186), .D(n291), .Y(n289) );
  ivd1_hd U151 ( .A(n68), .Y(n291) );
  ao21d1_hd U152 ( .A(n164), .B(n292), .C(n293), .Y(n327) );
  ao21d1_hd U153 ( .A(n73), .B(n334), .C(n164), .Y(n293) );
  ao22d1_hd U154 ( .A(n73), .B(n333), .C(n186), .D(n294), .Y(n292) );
  ivd1_hd U155 ( .A(n73), .Y(n294) );
  ao21d1_hd U156 ( .A(n165), .B(n295), .C(n296), .Y(n328) );
  ao21d1_hd U157 ( .A(n72), .B(n334), .C(n165), .Y(n296) );
  ao22d1_hd U158 ( .A(n72), .B(n333), .C(n186), .D(n297), .Y(n295) );
  ivd1_hd U159 ( .A(n72), .Y(n297) );
  ao21d1_hd U165 ( .A(n166), .B(n298), .C(n299), .Y(n329) );
  ao21d1_hd U166 ( .A(n71), .B(n334), .C(n166), .Y(n299) );
  ao22d1_hd U167 ( .A(n71), .B(n333), .C(n186), .D(n300), .Y(n298) );
  ivd1_hd U170 ( .A(n71), .Y(n300) );
  ad2d1_hd U172 ( .A(n334), .B(n156), .Y(n330) );
  ad2d1_hd U174 ( .A(n334), .B(n75), .Y(n331) );
  nr2d1_hd U178 ( .A(n301), .B(n36), .Y(n336) );
  nr3d1_hd U179 ( .A(n51), .B(n34), .C(n76), .Y(n301) );
endmodule


module ads1292_filter_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;

  had1_hd U2 ( .A(A[6]), .B(n2), .CO(n1), .S(SUM[6]) );
  had1_hd U3 ( .A(A[5]), .B(n3), .CO(n2), .S(SUM[5]) );
  had1_hd U4 ( .A(A[4]), .B(n4), .CO(n3), .S(SUM[4]) );
  had1_hd U5 ( .A(A[3]), .B(n5), .CO(n4), .S(SUM[3]) );
  had1_hd U6 ( .A(A[2]), .B(n6), .CO(n5), .S(SUM[2]) );
  had1_hd U7 ( .A(A[1]), .B(A[0]), .CO(n6), .S(SUM[1]) );
  xo2d1_hd U11 ( .A(n1), .B(A[7]), .Y(SUM[7]) );
  ivd1_hd U12 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_filter_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module ads1292_filter ( i_ADS1292_DATA_OUT, i_ADS1292_DATA_VALID, 
        o_ADS1292_FILTERED_DATA, o_ADS1292_FILTERED_DATA_VALID, 
        i_ADS1292_FILTERED_DATA_ACK, i_CLK, i_RSTN );
  input [23:0] i_ADS1292_DATA_OUT;
  output [23:0] o_ADS1292_FILTERED_DATA;
  input i_ADS1292_DATA_VALID, i_ADS1292_FILTERED_DATA_ACK, i_CLK, i_RSTN;
  output o_ADS1292_FILTERED_DATA_VALID;
  wire   w_rstn, w_rst, r_converter_i2f_a_stb, w_converter_i2f_a_ack,
         w_converter_i2f_z_stb, r_converter_i2f_z_ack, r_iir_lpf_x_valid,
         w_iir_lpf_x_ready, w_iir_lpf_y_valid, r_iir_lpf_y_ack,
         r_iir_notch_x_valid, w_iir_notch_x_ready, w_iir_notch_y_valid,
         r_iir_notch_y_ack, r_iir_hpf_x_valid, w_iir_hpf_x_ready,
         w_iir_hpf_y_valid, r_iir_hpf_y_ack, r_converter_f2i_a_stb,
         w_converter_f2i_a_ack, w_converter_f2i_z_stb, r_converter_f2i_z_ack,
         N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N50, N53, N56, N59, N60, N61, N62, N63, N86, N87, N88, N91, N94, N97,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N111, N121,
         N131, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N200, N201, N209,
         N216, N217, N218, N219, N220, N221, N222, N223, alt140_n29,
         alt140_n30, alt140_n31, alt140_n32, alt140_n90, alt140_n113,
         alt140_n114, alt140_n115, n1, n2, n4, n5, n6, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n640, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8;
  wire   [31:8] r_converter_i2f_a;
  wire   [31:0] w_converter_i2f_z;
  wire   [31:0] r_iir_lpf_x;
  wire   [31:0] w_iir_lpf_y;
  wire   [31:0] r_iir_notch_x;
  wire   [31:0] w_iir_notch_y;
  wire   [31:0] r_iir_hpf_x;
  wire   [31:0] w_iir_hpf_y;
  wire   [31:0] r_converter_f2i_a;
  wire   [31:8] w_converter_f2i_z;
  wire   [1:0] r_pstate;
  wire   [7:0] r_counter;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  async_rst_synchronizer async_rst_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RST(w_rst) );
  converter_i2f converter_i2f ( .i_A({r_converter_i2f_a, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .i_A_STB(r_converter_i2f_a_stb), 
        .o_A_ACK(w_converter_i2f_a_ack), .o_Z(w_converter_i2f_z), .o_Z_STB(
        w_converter_i2f_z_stb), .i_Z_ACK(r_converter_i2f_z_ack), .i_CLK(i_CLK), 
        .i_RST(w_rst) );
  iir_lpf iir_lpf ( .i_X_DATA(r_iir_lpf_x), .i_X_DATA_VALID(r_iir_lpf_x_valid), 
        .o_X_DATA_READY(w_iir_lpf_x_ready), .o_Y_DATA(w_iir_lpf_y), 
        .o_Y_DATA_VALID(w_iir_lpf_y_valid), .i_Y_ACK(r_iir_lpf_y_ack), .i_CLK(
        i_CLK), .i_RSTN(n427) );
  iir_notch iir_notch ( .i_X_DATA(r_iir_notch_x), .i_X_DATA_VALID(
        r_iir_notch_x_valid), .o_X_DATA_READY(w_iir_notch_x_ready), .o_Y_DATA(
        w_iir_notch_y), .o_Y_DATA_VALID(w_iir_notch_y_valid), .i_Y_ACK(
        r_iir_notch_y_ack), .i_CLK(i_CLK), .i_RSTN(n427) );
  iir_hpf iir_hpf ( .i_X_DATA(r_iir_hpf_x), .i_X_DATA_VALID(r_iir_hpf_x_valid), 
        .o_X_DATA_READY(w_iir_hpf_x_ready), .o_Y_DATA(w_iir_hpf_y), 
        .o_Y_DATA_VALID(w_iir_hpf_y_valid), .i_Y_ACK(r_iir_hpf_y_ack), .i_CLK(
        i_CLK), .i_RSTN(n427) );
  converter_f2i converter_f2i ( .i_A(r_converter_f2i_a), .i_A_STB(
        r_converter_f2i_a_stb), .o_A_ACK(w_converter_f2i_a_ack), .o_Z({
        w_converter_f2i_z, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8}), .o_Z_STB(w_converter_f2i_z_stb), .i_Z_ACK(r_converter_f2i_z_ack), .i_CLK(
        i_CLK), .i_RST(n628) );
  scg22d1_hd U12 ( .A(N46), .B(w_converter_i2f_a_ack), .C(n2), .D(N39), .Y(
        N192) );
  scg22d1_hd U13 ( .A(n422), .B(w_converter_f2i_a_ack), .C(n2), .D(N39), .Y(
        N191) );
  oa21d1_hd U14 ( .A(n2), .B(n4), .C(N39), .Y(N190) );
  oa21d1_hd U15 ( .A(n2), .B(n5), .C(N39), .Y(N189) );
  oa21d1_hd U16 ( .A(n2), .B(n6), .C(N39), .Y(N188) );
  oa211d1_hd U17 ( .A(alt140_n90), .B(n416), .C(n1), .D(N37), .Y(N187) );
  or2d1_hd U18 ( .A(n8), .B(n9), .Y(n1) );
  oa21d1_hd U19 ( .A(n9), .B(n10), .C(N37), .Y(N186) );
  oa21d1_hd U20 ( .A(n9), .B(n11), .C(N37), .Y(N185) );
  oa21d1_hd U21 ( .A(n9), .B(n12), .C(N37), .Y(N184) );
  oa21d1_hd U22 ( .A(n9), .B(n13), .C(N37), .Y(N183) );
  scg17d1_hd U24 ( .A(n15), .B(n16), .C(N169), .D(n17), .Y(N181) );
  oa31d1_hd U25 ( .A(n18), .B(n421), .C(N209), .D(N40), .Y(n17) );
  scg4d1_hd U26 ( .A(n417), .B(N121), .C(N87), .D(N101), .E(N111), .F(n420), 
        .G(n415), .H(N131), .Y(n18) );
  nd4d1_hd U27 ( .A(n19), .B(n4), .C(n5), .D(n6), .Y(n16) );
  ao22d1_hd U31 ( .A(n422), .B(w_converter_f2i_a_ack), .C(N46), .D(
        w_converter_i2f_a_ack), .Y(n19) );
  ivd1_hd U32 ( .A(n2), .Y(n15) );
  oa211d1_hd U34 ( .A(n21), .B(N37), .C(n22), .D(n14), .Y(N180) );
  nr2d1_hd U36 ( .A(N169), .B(n23), .Y(n22) );
  ao21d1_hd U38 ( .A(n422), .B(N63), .C(n24), .Y(n21) );
  nd4d1_hd U39 ( .A(alt140_n29), .B(n25), .C(n26), .D(n20), .Y(n24) );
  ao22d1_hd U40 ( .A(n419), .B(N61), .C(n424), .D(N62), .Y(n26) );
  ao22d1_hd U41 ( .A(N46), .B(N59), .C(n423), .D(N60), .Y(n25) );
  ad2d1_hd U42 ( .A(n27), .B(N109), .Y(N179) );
  ad2d1_hd U43 ( .A(n27), .B(N108), .Y(N178) );
  ad2d1_hd U44 ( .A(n27), .B(N107), .Y(N177) );
  ad2d1_hd U45 ( .A(n27), .B(N106), .Y(N176) );
  ad2d1_hd U46 ( .A(n27), .B(N105), .Y(N175) );
  ad2d1_hd U47 ( .A(n27), .B(N104), .Y(N174) );
  ad2d1_hd U48 ( .A(n27), .B(N103), .Y(N173) );
  ad2d1_hd U49 ( .A(n27), .B(N102), .Y(N172) );
  nr4d1_hd U52 ( .A(n417), .B(n420), .C(N87), .D(n415), .Y(n28) );
  or2d1_hd U53 ( .A(N36), .B(n23), .Y(N171) );
  ao21d1_hd U54 ( .A(n29), .B(n11), .C(n9), .Y(n23) );
  ivd1_hd U56 ( .A(n421), .Y(n20) );
  ad4d1_hd U58 ( .A(n12), .B(n13), .C(n8), .D(n10), .Y(n29) );
  nr2bd1_hd U63 ( .AN(n416), .B(alt140_n90), .Y(N169) );
  clknd2d1_hd U259 ( .A(w_converter_f2i_z_stb), .B(n418), .Y(n8) );
  clknd2d1_hd U260 ( .A(w_iir_hpf_y_valid), .B(n415), .Y(n10) );
  clknd2d1_hd U261 ( .A(w_converter_i2f_z_stb), .B(N87), .Y(n13) );
  clknd2d1_hd U262 ( .A(w_iir_lpf_y_valid), .B(n420), .Y(n12) );
  clknd2d1_hd U263 ( .A(w_iir_notch_y_valid), .B(n417), .Y(n11) );
  clknd2d1_hd U264 ( .A(N40), .B(n20), .Y(n9) );
  or2d1_hd U265 ( .A(n424), .B(alt140_n31), .Y(alt140_n30) );
  or2d1_hd U266 ( .A(n419), .B(alt140_n32), .Y(alt140_n31) );
  or2d1_hd U267 ( .A(n423), .B(N46), .Y(alt140_n32) );
  ivd1_hd U268 ( .A(w_iir_hpf_x_ready), .Y(N62) );
  ivd1_hd U269 ( .A(w_iir_notch_x_ready), .Y(N61) );
  ivd1_hd U270 ( .A(w_iir_lpf_x_ready), .Y(N60) );
  ivd1_hd U271 ( .A(w_converter_i2f_a_ack), .Y(N59) );
  or2d1_hd U272 ( .A(n420), .B(N87), .Y(alt140_n115) );
  ad2d1_hd U273 ( .A(N86), .B(N44), .Y(N87) );
  ad2d1_hd U274 ( .A(N42), .B(N43), .Y(N86) );
  ivd1_hd U275 ( .A(w_iir_hpf_y_valid), .Y(N131) );
  clknd2d1_hd U277 ( .A(n14), .B(N37), .Y(N182) );
  ad2d1_hd U278 ( .A(N34), .B(N35), .Y(N36) );
  ad2d1_hd U279 ( .A(r_pstate[1]), .B(r_pstate[0]), .Y(N41) );
  ivd1_hd U280 ( .A(N41), .Y(alt140_n90) );
  clknd2d1_hd U286 ( .A(alt140_n90), .B(n1), .Y(N193) );
  ad2d1_hd U287 ( .A(N184), .B(N37), .Y(N197) );
  or2d1_hd U288 ( .A(N34), .B(r_pstate[0]), .Y(N39) );
  ad2d1_hd U289 ( .A(N45), .B(N44), .Y(N46) );
  ad2d1_hd U290 ( .A(N42), .B(N43), .Y(N45) );
  clknd2d1_hd U291 ( .A(N36), .B(i_ADS1292_DATA_VALID), .Y(n14) );
  or2d2_hd U292 ( .A(r_pstate[1]), .B(N35), .Y(N37) );
  or2d1_hd U293 ( .A(n422), .B(alt140_n30), .Y(alt140_n29) );
  ad2d1_hd U294 ( .A(N220), .B(N221), .Y(N222) );
  ad2d1_hd U295 ( .A(N218), .B(N219), .Y(N220) );
  ad2d1_hd U296 ( .A(N216), .B(N217), .Y(N218) );
  or2d1_hd U297 ( .A(n418), .B(n425), .Y(N209) );
  or2d1_hd U298 ( .A(n415), .B(alt140_n114), .Y(alt140_n113) );
  or2d1_hd U299 ( .A(n417), .B(alt140_n115), .Y(alt140_n114) );
  ivd1_hd U300 ( .A(w_converter_i2f_z_stb), .Y(N101) );
  ivd1_hd U301 ( .A(w_iir_lpf_y_valid), .Y(N111) );
  ivd1_hd U302 ( .A(w_iir_notch_y_valid), .Y(N121) );
  clknd2d1_hd U303 ( .A(n424), .B(w_iir_hpf_x_ready), .Y(n4) );
  clknd2d1_hd U304 ( .A(n419), .B(w_iir_notch_x_ready), .Y(n5) );
  clknd2d1_hd U305 ( .A(n423), .B(w_iir_lpf_x_ready), .Y(n6) );
  clknd2d1_hd U306 ( .A(n20), .B(N38), .Y(n2) );
  ivd1_hd U307 ( .A(N39), .Y(N40) );
  or2d1_hd U333 ( .A(N36), .B(N41), .Y(N170) );
  mx2d1_hd U487 ( .D0(r_iir_lpf_y_ack), .D1(N40), .S(N184), .Y(n208) );
  mx2d1_hd U488 ( .D0(r_iir_hpf_x_valid), .D1(N38), .S(N190), .Y(n213) );
  mx2d1_hd U489 ( .D0(r_iir_lpf_x_valid), .D1(N38), .S(N188), .Y(n211) );
  mx2d1_hd U490 ( .D0(r_iir_notch_x_valid), .D1(N38), .S(N189), .Y(n212) );
  mx2d1_hd U491 ( .D0(r_converter_f2i_a_stb), .D1(N38), .S(N191), .Y(n214) );
  mx2d1_hd U492 ( .D0(r_converter_i2f_a_stb), .D1(N38), .S(N192), .Y(n215) );
  mx2d1_hd U493 ( .D0(r_converter_i2f_z_ack), .D1(N40), .S(N183), .Y(n207) );
  nid6_hd U494 ( .A(w_rstn), .Y(n426) );
  mx2d1_hd U495 ( .D0(r_iir_hpf_y_ack), .D1(N40), .S(N186), .Y(n210) );
  mx2d1_hd U496 ( .D0(r_iir_notch_y_ack), .D1(N40), .S(N185), .Y(n209) );
  ivd1_hd U497 ( .A(w_converter_f2i_a_ack), .Y(N63) );
  nr2ad1_hd U504 ( .A(n28), .B(N39), .Y(n27) );
  or2d1_hd U506 ( .A(N42), .B(r_counter[1]), .Y(N56) );
  ivd1_hd U507 ( .A(r_counter[1]), .Y(N43) );
  or2d1_hd U508 ( .A(N42), .B(r_counter[1]), .Y(N97) );
  or2d1_hd U510 ( .A(r_counter[2]), .B(N43), .Y(N53) );
  or2d1_hd U511 ( .A(r_counter[2]), .B(N43), .Y(N50) );
  or2d1_hd U512 ( .A(r_counter[2]), .B(r_counter[1]), .Y(N47) );
  or2d1_hd U513 ( .A(r_counter[2]), .B(N43), .Y(N91) );
  or2d1_hd U514 ( .A(r_counter[2]), .B(r_counter[1]), .Y(N88) );
  or2d1_hd U515 ( .A(r_counter[2]), .B(N43), .Y(N94) );
  ivd1_hd U516 ( .A(r_counter[2]), .Y(N42) );
  ivd1_hd U517 ( .A(r_counter[7]), .Y(N216) );
  nid6_hd U708 ( .A(w_rstn), .Y(n427) );
  nr2d1_hd U709 ( .A(N94), .B(N44), .Y(n415) );
  clknd2d1_hd U710 ( .A(o_ADS1292_FILTERED_DATA_VALID), .B(
        i_ADS1292_FILTERED_DATA_ACK), .Y(n416) );
  nr2d1_hd U711 ( .A(N91), .B(r_counter[0]), .Y(n417) );
  nr2d1_hd U712 ( .A(N97), .B(r_counter[0]), .Y(n418) );
  nr2d1_hd U713 ( .A(N50), .B(r_counter[0]), .Y(n419) );
  nr2d1_hd U714 ( .A(N88), .B(N44), .Y(n420) );
  clknd2d1_hd U715 ( .A(N222), .B(N223), .Y(n421) );
  ivd1_hd U716 ( .A(N37), .Y(N38) );
  nr2d1_hd U717 ( .A(N56), .B(r_counter[0]), .Y(n422) );
  nr2d1_hd U718 ( .A(N47), .B(N44), .Y(n423) );
  nr2d1_hd U719 ( .A(N53), .B(N44), .Y(n424) );
  nr2d1_hd U720 ( .A(n418), .B(alt140_n113), .Y(n425) );
  ads1292_filter_DW01_inc_0 add_x_1 ( .A(r_counter), .SUM({N109, N108, N107, 
        N106, N105, N104, N103, N102}) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_10 clk_gate_r_iir_notch_y_ack_reg_0 ( 
        .CLK(i_CLK), .EN(n640), .ENCLK(n636), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_11 clk_gate_r_counter_reg_2__0 ( .CLK(
        i_CLK), .EN(N171), .ENCLK(n635), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_12 clk_gate_o_ADS1292_FILTERED_DATA_reg_23__0 ( 
        .CLK(i_CLK), .EN(N200), .ENCLK(n634), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_13 clk_gate_r_converter_i2f_a_reg_31__0 ( 
        .CLK(i_CLK), .EN(N201), .ENCLK(n633), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_14 clk_gate_r_converter_f2i_a_reg_31__0 ( 
        .CLK(i_CLK), .EN(N194), .ENCLK(n632), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_15 clk_gate_r_iir_hpf_x_reg_31__0 ( 
        .CLK(i_CLK), .EN(N196), .ENCLK(n631), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_16 clk_gate_r_iir_lpf_x_reg_31__0 ( 
        .CLK(i_CLK), .EN(N195), .ENCLK(n630), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_filter_17 clk_gate_r_iir_notch_x_reg_31__0 ( 
        .CLK(i_CLK), .EN(N197), .ENCLK(n629), .TE(1'b0) );
  fd2qd1_hd r_iir_notch_x_reg_28_ ( .D(w_iir_lpf_y[28]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[28]) );
  fd2qd1_hd r_iir_notch_x_reg_27_ ( .D(w_iir_lpf_y[27]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[27]) );
  fd2qd1_hd r_iir_notch_x_reg_26_ ( .D(w_iir_lpf_y[26]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[26]) );
  fd2qd1_hd r_iir_notch_x_reg_25_ ( .D(w_iir_lpf_y[25]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[25]) );
  fd2qd1_hd r_iir_notch_x_reg_24_ ( .D(w_iir_lpf_y[24]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[24]) );
  fd2qd1_hd r_iir_notch_x_reg_23_ ( .D(w_iir_lpf_y[23]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[23]) );
  fd2qd1_hd r_iir_notch_x_reg_22_ ( .D(w_iir_lpf_y[22]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[22]) );
  fd2qd1_hd r_iir_notch_x_reg_21_ ( .D(w_iir_lpf_y[21]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[21]) );
  fd2qd1_hd r_iir_notch_x_reg_20_ ( .D(w_iir_lpf_y[20]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[20]) );
  fd2qd1_hd r_iir_notch_x_reg_19_ ( .D(w_iir_lpf_y[19]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[19]) );
  fd2qd1_hd r_iir_notch_x_reg_18_ ( .D(w_iir_lpf_y[18]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[18]) );
  fd2qd1_hd r_iir_notch_x_reg_17_ ( .D(w_iir_lpf_y[17]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[17]) );
  fd2qd1_hd r_iir_notch_x_reg_16_ ( .D(w_iir_lpf_y[16]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[16]) );
  fd2qd1_hd r_iir_notch_x_reg_15_ ( .D(w_iir_lpf_y[15]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[15]) );
  fd2qd1_hd r_iir_notch_x_reg_14_ ( .D(w_iir_lpf_y[14]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[14]) );
  fd2qd1_hd r_iir_notch_x_reg_13_ ( .D(w_iir_lpf_y[13]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[13]) );
  fd2qd1_hd r_iir_notch_x_reg_12_ ( .D(w_iir_lpf_y[12]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[12]) );
  fd2qd1_hd r_iir_notch_x_reg_11_ ( .D(w_iir_lpf_y[11]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[11]) );
  fd2qd1_hd r_iir_notch_x_reg_10_ ( .D(w_iir_lpf_y[10]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[10]) );
  fd2qd1_hd r_iir_notch_x_reg_9_ ( .D(w_iir_lpf_y[9]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[9]) );
  fd2qd1_hd r_iir_notch_x_reg_8_ ( .D(w_iir_lpf_y[8]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[8]) );
  fd2qd1_hd r_iir_notch_x_reg_7_ ( .D(w_iir_lpf_y[7]), .CK(n629), .RN(n427), 
        .Q(r_iir_notch_x[7]) );
  fd2qd1_hd r_iir_hpf_x_reg_31_ ( .D(w_iir_notch_y[31]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[31]) );
  fd2qd1_hd r_iir_hpf_x_reg_30_ ( .D(w_iir_notch_y[30]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[30]) );
  fd2qd1_hd r_iir_hpf_x_reg_29_ ( .D(w_iir_notch_y[29]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[29]) );
  fd2qd1_hd r_iir_hpf_x_reg_28_ ( .D(w_iir_notch_y[28]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[28]) );
  fd2qd1_hd r_iir_hpf_x_reg_27_ ( .D(w_iir_notch_y[27]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[27]) );
  fd2qd1_hd r_iir_hpf_x_reg_26_ ( .D(w_iir_notch_y[26]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[26]) );
  fd2qd1_hd r_iir_hpf_x_reg_25_ ( .D(w_iir_notch_y[25]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[25]) );
  fd2qd1_hd r_iir_hpf_x_reg_24_ ( .D(w_iir_notch_y[24]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[24]) );
  fd2qd1_hd r_iir_hpf_x_reg_23_ ( .D(w_iir_notch_y[23]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[23]) );
  fd2qd1_hd r_iir_hpf_x_reg_22_ ( .D(w_iir_notch_y[22]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[22]) );
  fd2qd1_hd r_iir_hpf_x_reg_21_ ( .D(w_iir_notch_y[21]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[21]) );
  fd2qd1_hd r_iir_hpf_x_reg_20_ ( .D(w_iir_notch_y[20]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[20]) );
  fd2qd1_hd r_iir_hpf_x_reg_19_ ( .D(w_iir_notch_y[19]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[19]) );
  fd2qd1_hd r_iir_hpf_x_reg_18_ ( .D(w_iir_notch_y[18]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[18]) );
  fd2qd1_hd r_iir_hpf_x_reg_17_ ( .D(w_iir_notch_y[17]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[17]) );
  fd2qd1_hd r_iir_hpf_x_reg_16_ ( .D(w_iir_notch_y[16]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[16]) );
  fd2qd1_hd r_iir_hpf_x_reg_15_ ( .D(w_iir_notch_y[15]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[15]) );
  fd2qd1_hd r_iir_hpf_x_reg_14_ ( .D(w_iir_notch_y[14]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[14]) );
  fd2qd1_hd r_iir_hpf_x_reg_13_ ( .D(w_iir_notch_y[13]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[13]) );
  fd2qd1_hd r_iir_hpf_x_reg_12_ ( .D(w_iir_notch_y[12]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[12]) );
  fd2qd1_hd r_iir_hpf_x_reg_11_ ( .D(w_iir_notch_y[11]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[11]) );
  fd2qd1_hd r_iir_hpf_x_reg_10_ ( .D(w_iir_notch_y[10]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[10]) );
  fd2qd1_hd r_iir_hpf_x_reg_9_ ( .D(w_iir_notch_y[9]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[9]) );
  fd2qd1_hd r_iir_hpf_x_reg_7_ ( .D(w_iir_notch_y[7]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[7]) );
  fd2qd1_hd r_iir_hpf_x_reg_6_ ( .D(w_iir_notch_y[6]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[6]) );
  fd2qd1_hd r_iir_hpf_x_reg_5_ ( .D(w_iir_notch_y[5]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[5]) );
  fd2qd1_hd r_iir_hpf_x_reg_4_ ( .D(w_iir_notch_y[4]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[4]) );
  fd2qd1_hd r_iir_hpf_x_reg_3_ ( .D(w_iir_notch_y[3]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[3]) );
  fd2qd1_hd r_iir_hpf_x_reg_2_ ( .D(w_iir_notch_y[2]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[2]) );
  fd2qd1_hd r_iir_hpf_x_reg_1_ ( .D(w_iir_notch_y[1]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[1]) );
  fd2qd1_hd r_iir_hpf_x_reg_0_ ( .D(w_iir_notch_y[0]), .CK(n631), .RN(n427), 
        .Q(r_iir_hpf_x[0]) );
  fd2qd1_hd r_converter_f2i_a_reg_31_ ( .D(w_iir_hpf_y[31]), .CK(n632), .RN(
        n427), .Q(r_converter_f2i_a[31]) );
  fd2qd1_hd r_converter_f2i_a_reg_30_ ( .D(w_iir_hpf_y[30]), .CK(n632), .RN(
        n427), .Q(r_converter_f2i_a[30]) );
  fd2qd1_hd r_converter_f2i_a_reg_29_ ( .D(w_iir_hpf_y[29]), .CK(n632), .RN(
        n427), .Q(r_converter_f2i_a[29]) );
  fd2qd1_hd r_converter_f2i_a_reg_28_ ( .D(w_iir_hpf_y[28]), .CK(n632), .RN(
        n427), .Q(r_converter_f2i_a[28]) );
  fd2qd1_hd r_converter_f2i_a_reg_27_ ( .D(w_iir_hpf_y[27]), .CK(n632), .RN(
        n427), .Q(r_converter_f2i_a[27]) );
  fd2qd1_hd r_converter_f2i_a_reg_26_ ( .D(w_iir_hpf_y[26]), .CK(n632), .RN(
        n427), .Q(r_converter_f2i_a[26]) );
  fd2qd1_hd r_converter_f2i_a_reg_25_ ( .D(w_iir_hpf_y[25]), .CK(n632), .RN(
        n427), .Q(r_converter_f2i_a[25]) );
  fd2qd1_hd r_converter_f2i_a_reg_0_ ( .D(w_iir_hpf_y[0]), .CK(n632), .RN(n427), .Q(r_converter_f2i_a[0]) );
  fd2qd1_hd r_iir_notch_x_reg_31_ ( .D(w_iir_lpf_y[31]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[31]) );
  fd2qd1_hd r_iir_notch_x_reg_30_ ( .D(w_iir_lpf_y[30]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[30]) );
  fd2qd1_hd r_iir_notch_x_reg_29_ ( .D(w_iir_lpf_y[29]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[29]) );
  fd2qd1_hd r_iir_notch_x_reg_6_ ( .D(w_iir_lpf_y[6]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[6]) );
  fd2qd1_hd r_iir_notch_x_reg_5_ ( .D(w_iir_lpf_y[5]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[5]) );
  fd2qd1_hd r_iir_notch_x_reg_4_ ( .D(w_iir_lpf_y[4]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[4]) );
  fd2qd1_hd r_iir_notch_x_reg_3_ ( .D(w_iir_lpf_y[3]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[3]) );
  fd2qd1_hd r_iir_notch_x_reg_2_ ( .D(w_iir_lpf_y[2]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[2]) );
  fd2qd1_hd r_iir_notch_x_reg_1_ ( .D(w_iir_lpf_y[1]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[1]) );
  fd2qd1_hd r_iir_notch_x_reg_0_ ( .D(w_iir_lpf_y[0]), .CK(n629), .RN(n426), 
        .Q(r_iir_notch_x[0]) );
  fd2qd1_hd r_iir_lpf_x_reg_31_ ( .D(w_converter_i2f_z[31]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[31]) );
  fd2qd1_hd r_iir_lpf_x_reg_30_ ( .D(w_converter_i2f_z[30]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[30]) );
  fd2qd1_hd r_iir_lpf_x_reg_29_ ( .D(w_converter_i2f_z[29]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[29]) );
  fd2qd1_hd r_iir_lpf_x_reg_28_ ( .D(w_converter_i2f_z[28]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[28]) );
  fd2qd1_hd r_iir_lpf_x_reg_27_ ( .D(w_converter_i2f_z[27]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[27]) );
  fd2qd1_hd r_iir_lpf_x_reg_26_ ( .D(w_converter_i2f_z[26]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[26]) );
  fd2qd1_hd r_iir_lpf_x_reg_25_ ( .D(w_converter_i2f_z[25]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[25]) );
  fd2qd1_hd r_iir_lpf_x_reg_24_ ( .D(w_converter_i2f_z[24]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[24]) );
  fd2qd1_hd r_iir_lpf_x_reg_23_ ( .D(w_converter_i2f_z[23]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[23]) );
  fd2qd1_hd r_iir_lpf_x_reg_22_ ( .D(w_converter_i2f_z[22]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[22]) );
  fd2qd1_hd r_iir_lpf_x_reg_21_ ( .D(w_converter_i2f_z[21]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[21]) );
  fd2qd1_hd r_iir_lpf_x_reg_20_ ( .D(w_converter_i2f_z[20]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[20]) );
  fd2qd1_hd r_iir_lpf_x_reg_19_ ( .D(w_converter_i2f_z[19]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[19]) );
  fd2qd1_hd r_iir_lpf_x_reg_18_ ( .D(w_converter_i2f_z[18]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[18]) );
  fd2qd1_hd r_iir_lpf_x_reg_17_ ( .D(w_converter_i2f_z[17]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[17]) );
  fd2qd1_hd r_iir_lpf_x_reg_16_ ( .D(w_converter_i2f_z[16]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[16]) );
  fd2qd1_hd r_iir_lpf_x_reg_15_ ( .D(w_converter_i2f_z[15]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[15]) );
  fd2qd1_hd r_iir_lpf_x_reg_14_ ( .D(w_converter_i2f_z[14]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[14]) );
  fd2qd1_hd r_iir_lpf_x_reg_13_ ( .D(w_converter_i2f_z[13]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[13]) );
  fd2qd1_hd r_iir_lpf_x_reg_12_ ( .D(w_converter_i2f_z[12]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[12]) );
  fd2qd1_hd r_iir_lpf_x_reg_11_ ( .D(w_converter_i2f_z[11]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[11]) );
  fd2qd1_hd r_iir_lpf_x_reg_10_ ( .D(w_converter_i2f_z[10]), .CK(n630), .RN(
        n426), .Q(r_iir_lpf_x[10]) );
  fd2qd1_hd r_iir_lpf_x_reg_9_ ( .D(w_converter_i2f_z[9]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[9]) );
  fd2qd1_hd r_iir_lpf_x_reg_8_ ( .D(w_converter_i2f_z[8]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[8]) );
  fd2qd1_hd r_iir_lpf_x_reg_7_ ( .D(w_converter_i2f_z[7]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[7]) );
  fd2qd1_hd r_iir_lpf_x_reg_6_ ( .D(w_converter_i2f_z[6]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[6]) );
  fd2qd1_hd r_iir_lpf_x_reg_5_ ( .D(w_converter_i2f_z[5]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[5]) );
  fd2qd1_hd r_iir_lpf_x_reg_4_ ( .D(w_converter_i2f_z[4]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[4]) );
  fd2qd1_hd r_iir_lpf_x_reg_3_ ( .D(w_converter_i2f_z[3]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[3]) );
  fd2qd1_hd r_iir_lpf_x_reg_2_ ( .D(w_converter_i2f_z[2]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[2]) );
  fd2qd1_hd r_iir_lpf_x_reg_1_ ( .D(w_converter_i2f_z[1]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[1]) );
  fd2qd1_hd r_iir_lpf_x_reg_0_ ( .D(w_converter_i2f_z[0]), .CK(n630), .RN(n426), .Q(r_iir_lpf_x[0]) );
  fd2qd1_hd r_iir_hpf_x_reg_8_ ( .D(w_iir_notch_y[8]), .CK(n631), .RN(n426), 
        .Q(r_iir_hpf_x[8]) );
  fd2qd1_hd r_converter_f2i_a_reg_24_ ( .D(w_iir_hpf_y[24]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[24]) );
  fd2qd1_hd r_converter_f2i_a_reg_23_ ( .D(w_iir_hpf_y[23]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[23]) );
  fd2qd1_hd r_converter_f2i_a_reg_22_ ( .D(w_iir_hpf_y[22]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[22]) );
  fd2qd1_hd r_converter_f2i_a_reg_21_ ( .D(w_iir_hpf_y[21]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[21]) );
  fd2qd1_hd r_converter_f2i_a_reg_20_ ( .D(w_iir_hpf_y[20]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[20]) );
  fd2qd1_hd r_converter_f2i_a_reg_19_ ( .D(w_iir_hpf_y[19]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[19]) );
  fd2qd1_hd r_converter_f2i_a_reg_18_ ( .D(w_iir_hpf_y[18]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[18]) );
  fd2qd1_hd r_converter_f2i_a_reg_17_ ( .D(w_iir_hpf_y[17]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[17]) );
  fd2qd1_hd r_converter_f2i_a_reg_16_ ( .D(w_iir_hpf_y[16]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[16]) );
  fd2qd1_hd r_converter_f2i_a_reg_15_ ( .D(w_iir_hpf_y[15]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[15]) );
  fd2qd1_hd r_converter_f2i_a_reg_14_ ( .D(w_iir_hpf_y[14]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[14]) );
  fd2qd1_hd r_converter_f2i_a_reg_13_ ( .D(w_iir_hpf_y[13]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[13]) );
  fd2qd1_hd r_converter_f2i_a_reg_12_ ( .D(w_iir_hpf_y[12]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[12]) );
  fd2qd1_hd r_converter_f2i_a_reg_11_ ( .D(w_iir_hpf_y[11]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[11]) );
  fd2qd1_hd r_converter_f2i_a_reg_10_ ( .D(w_iir_hpf_y[10]), .CK(n632), .RN(
        n426), .Q(r_converter_f2i_a[10]) );
  fd2qd1_hd r_converter_f2i_a_reg_9_ ( .D(w_iir_hpf_y[9]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[9]) );
  fd2qd1_hd r_converter_f2i_a_reg_8_ ( .D(w_iir_hpf_y[8]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[8]) );
  fd2qd1_hd r_converter_f2i_a_reg_7_ ( .D(w_iir_hpf_y[7]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[7]) );
  fd2qd1_hd r_converter_f2i_a_reg_6_ ( .D(w_iir_hpf_y[6]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[6]) );
  fd2qd1_hd r_converter_f2i_a_reg_5_ ( .D(w_iir_hpf_y[5]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[5]) );
  fd2qd1_hd r_converter_f2i_a_reg_4_ ( .D(w_iir_hpf_y[4]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[4]) );
  fd2qd1_hd r_converter_f2i_a_reg_3_ ( .D(w_iir_hpf_y[3]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[3]) );
  fd2qd1_hd r_converter_f2i_a_reg_2_ ( .D(w_iir_hpf_y[2]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[2]) );
  fd2qd1_hd r_converter_f2i_a_reg_1_ ( .D(w_iir_hpf_y[1]), .CK(n632), .RN(n426), .Q(r_converter_f2i_a[1]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_23_ ( .D(w_converter_f2i_z[31]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[23]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_22_ ( .D(w_converter_f2i_z[30]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[22]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_21_ ( .D(w_converter_f2i_z[29]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[21]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_20_ ( .D(w_converter_f2i_z[28]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[20]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_19_ ( .D(w_converter_f2i_z[27]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[19]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_18_ ( .D(w_converter_f2i_z[26]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[18]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_17_ ( .D(w_converter_f2i_z[25]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[17]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_16_ ( .D(w_converter_f2i_z[24]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[16]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_15_ ( .D(w_converter_f2i_z[23]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[15]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_14_ ( .D(w_converter_f2i_z[22]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[14]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_13_ ( .D(w_converter_f2i_z[21]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[13]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_12_ ( .D(w_converter_f2i_z[20]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[12]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_11_ ( .D(w_converter_f2i_z[19]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[11]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_10_ ( .D(w_converter_f2i_z[18]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[10]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_9_ ( .D(w_converter_f2i_z[17]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[9]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_8_ ( .D(w_converter_f2i_z[16]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[8]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_7_ ( .D(w_converter_f2i_z[15]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[7]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_6_ ( .D(w_converter_f2i_z[14]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[6]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_5_ ( .D(w_converter_f2i_z[13]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[5]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_4_ ( .D(w_converter_f2i_z[12]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[4]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_3_ ( .D(w_converter_f2i_z[11]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[3]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_2_ ( .D(w_converter_f2i_z[10]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[2]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_1_ ( .D(w_converter_f2i_z[9]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[1]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_0_ ( .D(w_converter_f2i_z[8]), .CK(
        n634), .RN(n426), .Q(o_ADS1292_FILTERED_DATA[0]) );
  fd2qd1_hd r_counter_reg_7_ ( .D(N179), .CK(n635), .RN(n427), .Q(r_counter[7]) );
  fd2qd1_hd r_counter_reg_2_ ( .D(N174), .CK(n635), .RN(n426), .Q(r_counter[2]) );
  fd2qd1_hd r_counter_reg_1_ ( .D(N173), .CK(n635), .RN(n426), .Q(r_counter[1]) );
  fd2qd1_hd r_converter_i2f_a_stb_reg ( .D(n215), .CK(n636), .RN(n426), .Q(
        r_converter_i2f_a_stb) );
  fd2qd1_hd r_converter_f2i_a_stb_reg ( .D(n214), .CK(n636), .RN(n426), .Q(
        r_converter_f2i_a_stb) );
  fd2qd1_hd r_iir_notch_x_valid_reg ( .D(n212), .CK(n636), .RN(n426), .Q(
        r_iir_notch_x_valid) );
  fd2qd1_hd r_iir_lpf_x_valid_reg ( .D(n211), .CK(n636), .RN(n426), .Q(
        r_iir_lpf_x_valid) );
  fd2qd1_hd r_iir_hpf_x_valid_reg ( .D(n213), .CK(n636), .RN(n426), .Q(
        r_iir_hpf_x_valid) );
  fd2qd1_hd r_iir_lpf_y_ack_reg ( .D(n208), .CK(n636), .RN(n427), .Q(
        r_iir_lpf_y_ack) );
  fd2qd1_hd r_iir_notch_y_ack_reg ( .D(n209), .CK(n636), .RN(n427), .Q(
        r_iir_notch_y_ack) );
  fd2qd1_hd r_iir_hpf_y_ack_reg ( .D(n210), .CK(n636), .RN(n426), .Q(
        r_iir_hpf_y_ack) );
  fd2qd1_hd r_converter_i2f_z_ack_reg ( .D(n207), .CK(n636), .RN(n426), .Q(
        r_converter_i2f_z_ack) );
  fd2qd1_hd r_converter_i2f_a_reg_31_ ( .D(i_ADS1292_DATA_OUT[23]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[31]) );
  fd2qd1_hd r_converter_i2f_a_reg_30_ ( .D(i_ADS1292_DATA_OUT[22]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[30]) );
  fd2qd1_hd r_converter_i2f_a_reg_29_ ( .D(i_ADS1292_DATA_OUT[21]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[29]) );
  fd2qd1_hd r_converter_i2f_a_reg_28_ ( .D(i_ADS1292_DATA_OUT[20]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[28]) );
  fd2qd1_hd r_converter_i2f_a_reg_27_ ( .D(i_ADS1292_DATA_OUT[19]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[27]) );
  fd2qd1_hd r_converter_i2f_a_reg_26_ ( .D(i_ADS1292_DATA_OUT[18]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[26]) );
  fd2qd1_hd r_converter_i2f_a_reg_25_ ( .D(i_ADS1292_DATA_OUT[17]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[25]) );
  fd2qd1_hd r_converter_i2f_a_reg_24_ ( .D(i_ADS1292_DATA_OUT[16]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[24]) );
  fd2qd1_hd r_converter_i2f_a_reg_23_ ( .D(i_ADS1292_DATA_OUT[15]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[23]) );
  fd2qd1_hd r_converter_i2f_a_reg_22_ ( .D(i_ADS1292_DATA_OUT[14]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[22]) );
  fd2qd1_hd r_converter_i2f_a_reg_21_ ( .D(i_ADS1292_DATA_OUT[13]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[21]) );
  fd2qd1_hd r_converter_i2f_a_reg_20_ ( .D(i_ADS1292_DATA_OUT[12]), .CK(n633), 
        .RN(n426), .Q(r_converter_i2f_a[20]) );
  fd2qd1_hd r_converter_i2f_a_reg_19_ ( .D(i_ADS1292_DATA_OUT[11]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[19]) );
  fd2qd1_hd r_converter_i2f_a_reg_18_ ( .D(i_ADS1292_DATA_OUT[10]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[18]) );
  fd2qd1_hd r_converter_i2f_a_reg_17_ ( .D(i_ADS1292_DATA_OUT[9]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[17]) );
  fd2qd1_hd r_converter_i2f_a_reg_16_ ( .D(i_ADS1292_DATA_OUT[8]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[16]) );
  fd2qd1_hd r_converter_i2f_a_reg_15_ ( .D(i_ADS1292_DATA_OUT[7]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[15]) );
  fd2qd1_hd r_converter_i2f_a_reg_14_ ( .D(i_ADS1292_DATA_OUT[6]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[14]) );
  fd2qd1_hd r_converter_i2f_a_reg_13_ ( .D(i_ADS1292_DATA_OUT[5]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[13]) );
  fd2qd1_hd r_converter_i2f_a_reg_12_ ( .D(i_ADS1292_DATA_OUT[4]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[12]) );
  fd2qd1_hd r_converter_i2f_a_reg_11_ ( .D(i_ADS1292_DATA_OUT[3]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[11]) );
  fd2qd1_hd r_converter_i2f_a_reg_10_ ( .D(i_ADS1292_DATA_OUT[2]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[10]) );
  fd2qd1_hd r_converter_i2f_a_reg_9_ ( .D(i_ADS1292_DATA_OUT[1]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[9]) );
  fd2qd1_hd r_converter_i2f_a_reg_8_ ( .D(i_ADS1292_DATA_OUT[0]), .CK(n633), 
        .RN(n427), .Q(r_converter_i2f_a[8]) );
  fd2qd1_hd r_converter_f2i_z_ack_reg ( .D(n637), .CK(i_CLK), .RN(n426), .Q(
        r_converter_f2i_z_ack) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_VALID_reg ( .D(n638), .CK(i_CLK), .RN(n427), .Q(o_ADS1292_FILTERED_DATA_VALID) );
  fd2qd1_hd r_counter_reg_6_ ( .D(N178), .CK(n635), .RN(n427), .Q(r_counter[6]) );
  fd2qd1_hd r_counter_reg_5_ ( .D(N177), .CK(n635), .RN(n427), .Q(r_counter[5]) );
  fd2qd1_hd r_counter_reg_4_ ( .D(N176), .CK(n635), .RN(n427), .Q(r_counter[4]) );
  fd2qd1_hd r_counter_reg_3_ ( .D(N175), .CK(n635), .RN(n427), .Q(r_counter[3]) );
  fd2qd1_hd r_counter_reg_0_ ( .D(N172), .CK(n635), .RN(n427), .Q(r_counter[0]) );
  fd2qd1_hd r_pstate_reg_1_ ( .D(N181), .CK(i_CLK), .RN(n427), .Q(r_pstate[1])
         );
  fd2qd1_hd r_pstate_reg_0_ ( .D(N180), .CK(i_CLK), .RN(n427), .Q(r_pstate[0])
         );
  ivd1_hd U1 ( .A(r_counter[5]), .Y(N219) );
  ivd1_hd U2 ( .A(r_counter[6]), .Y(N217) );
  ivd1_hd U3 ( .A(r_pstate[0]), .Y(N35) );
  ivd1_hd U4 ( .A(r_counter[0]), .Y(N44) );
  ivd1_hd U5 ( .A(r_pstate[1]), .Y(N34) );
  ivd1_hd U6 ( .A(r_counter[3]), .Y(N223) );
  ivd1_hd U7 ( .A(r_counter[4]), .Y(N221) );
  ad2d1_hd U8 ( .A(N183), .B(N37), .Y(N195) );
  ad2d1_hd U9 ( .A(N185), .B(N37), .Y(N196) );
  ad2d1_hd U10 ( .A(N186), .B(N37), .Y(N194) );
  ad2d1_hd U11 ( .A(N182), .B(N37), .Y(N201) );
  ad2d1_hd U23 ( .A(N193), .B(alt140_n90), .Y(N200) );
  mx2d1_hd U28 ( .D0(r_pstate[1]), .D1(N34), .S(r_pstate[0]), .Y(n640) );
  mx2d1_hd U29 ( .D0(o_ADS1292_FILTERED_DATA_VALID), .D1(N169), .S(N170), .Y(
        n638) );
  mx2d1_hd U30 ( .D0(r_converter_f2i_z_ack), .D1(N40), .S(N187), .Y(n637) );
  nid1_hd U33 ( .A(w_rst), .Y(n628) );
endmodule


module spi_master_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  had1_hd U2 ( .A(A[12]), .B(n2), .CO(n1), .S(SUM[12]) );
  had1_hd U3 ( .A(A[11]), .B(n3), .CO(n2), .S(SUM[11]) );
  had1_hd U4 ( .A(A[10]), .B(n4), .CO(n3), .S(SUM[10]) );
  had1_hd U5 ( .A(A[9]), .B(n5), .CO(n4), .S(SUM[9]) );
  had1_hd U6 ( .A(A[8]), .B(n6), .CO(n5), .S(SUM[8]) );
  had1_hd U7 ( .A(A[7]), .B(n7), .CO(n6), .S(SUM[7]) );
  had1_hd U8 ( .A(A[6]), .B(n8), .CO(n7), .S(SUM[6]) );
  had1_hd U9 ( .A(A[5]), .B(n9), .CO(n8), .S(SUM[5]) );
  had1_hd U10 ( .A(A[4]), .B(n10), .CO(n9), .S(SUM[4]) );
  had1_hd U11 ( .A(A[3]), .B(n11), .CO(n10), .S(SUM[3]) );
  had1_hd U12 ( .A(A[2]), .B(n12), .CO(n11), .S(SUM[2]) );
  had1_hd U13 ( .A(A[1]), .B(A[0]), .CO(n12), .S(SUM[1]) );
  xo2d1_hd U17 ( .A(n1), .B(A[13]), .Y(SUM[13]) );
  ivd1_hd U18 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_spi_master_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_spi_master_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_spi_master_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module spi_master ( i_RSTN, i_CLK, i_TX_Byte, i_TX_DV, o_TX_Ready, o_RX_DV, 
        o_RX_Byte, o_SPI_Clk, i_SPI_MISO, o_SPI_MOSI );
  input [7:0] i_TX_Byte;
  output [7:0] o_RX_Byte;
  input i_RSTN, i_CLK, i_TX_DV, i_SPI_MISO;
  output o_TX_Ready, o_RX_DV, o_SPI_Clk, o_SPI_MOSI;
  wire   n90, n91, n92, n93, n94, n95, n96, n97, n89, n98, N0, N1, N11, w_rstn,
         r_SPI_Clk, N23, N26, N31, N32, N33, N34, N35, N36, N37, N38, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N75, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N110, N116, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N134, N139, N140,
         N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
         N152, N154, N155, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, alt9_n41, sub_x_13_n1,
         sub_x_11_n1, n1, n2, n3, n27, n30, n31, n32, n60, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n53, n54, n55, n56, n57, n58,
         n59, n61, n84, n86, n87, n88, n99, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n144, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158;
  wire   [7:0] r_SPI_Clk_Edges;
  wire   [3:0] r_SPI_Clk_Count;
  wire   [2:0] r_TX_Bit_Count;
  wire   [2:0] r_RX_Bit_Count;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  ivd1_hd U26 ( .A(N188), .Y(N189) );
  ivd1_hd U28 ( .A(n3), .Y(N110) );
  ivd1_hd U30 ( .A(i_TX_DV), .Y(n1) );
  or2d1_hd U34 ( .A(n86), .B(n60), .Y(N99) );
  ad2d1_hd U35 ( .A(n62), .B(N154), .Y(n89) );
  ad2d1_hd U36 ( .A(N194), .B(N154), .Y(N152) );
  ad2d1_hd U37 ( .A(N196), .B(N154), .Y(N151) );
  ad2d1_hd U38 ( .A(N198), .B(N154), .Y(N150) );
  ad2d1_hd U39 ( .A(N200), .B(N154), .Y(N149) );
  ad2d1_hd U40 ( .A(N202), .B(N154), .Y(N148) );
  ad2d1_hd U41 ( .A(N204), .B(N154), .Y(N147) );
  ad2d1_hd U42 ( .A(N206), .B(N154), .Y(N146) );
  ad2d1_hd U43 ( .A(N208), .B(N154), .Y(N145) );
  scg6d1_hd U44 ( .A(N154), .B(N140), .C(o_TX_Ready), .Y(N143) );
  scg6d1_hd U45 ( .A(N154), .B(N139), .C(o_TX_Ready), .Y(N142) );
  scg16d1_hd U46 ( .A(N154), .B(n40), .C(alt9_n41), .Y(N141) );
  ad2d1_hd U47 ( .A(N121), .B(N126), .Y(N127) );
  scg6d1_hd U48 ( .A(N126), .B(N120), .C(o_TX_Ready), .Y(N124) );
  scg6d1_hd U49 ( .A(N126), .B(N119), .C(o_TX_Ready), .Y(N123) );
  scg16d1_hd U50 ( .A(N126), .B(n37), .C(alt9_n41), .Y(N122) );
  ivd1_hd U54 ( .A(n30), .Y(N134) );
  ivd1_hd U55 ( .A(n31), .Y(N116) );
  ad2d1_hd U56 ( .A(N38), .B(n32), .Y(N107) );
  ad2d1_hd U57 ( .A(N37), .B(n32), .Y(N106) );
  ad2d1_hd U58 ( .A(N36), .B(n32), .Y(N105) );
  scg6d1_hd U59 ( .A(N35), .B(n32), .C(n86), .Y(N104) );
  ad2d1_hd U60 ( .A(N34), .B(n32), .Y(N103) );
  ad2d1_hd U61 ( .A(N33), .B(n32), .Y(N102) );
  ad2d1_hd U62 ( .A(N32), .B(n32), .Y(N101) );
  ad2d1_hd U63 ( .A(N31), .B(n32), .Y(N100) );
  clknd2d1_hd U93 ( .A(n30), .B(n31), .Y(n32) );
  or2d1_hd U94 ( .A(n28), .B(N177), .Y(N178) );
  or2d1_hd U95 ( .A(n26), .B(N176), .Y(N177) );
  or2d1_hd U96 ( .A(n25), .B(n12), .Y(N176) );
  or2d1_hd U97 ( .A(n26), .B(N160), .Y(N161) );
  or2d1_hd U98 ( .A(n25), .B(n12), .Y(N160) );
  or2d1_hd U99 ( .A(n35), .B(N181), .Y(N182) );
  or2d1_hd U100 ( .A(n34), .B(N180), .Y(N181) );
  or2d1_hd U101 ( .A(n33), .B(N179), .Y(N180) );
  or2d1_hd U102 ( .A(n29), .B(N178), .Y(N179) );
  or2d1_hd U103 ( .A(n34), .B(N164), .Y(N165) );
  or2d1_hd U104 ( .A(n33), .B(N163), .Y(N164) );
  or2d1_hd U105 ( .A(n29), .B(N162), .Y(N163) );
  or2d1_hd U106 ( .A(n28), .B(N161), .Y(N162) );
  or2d1_hd U107 ( .A(N174), .B(N184), .Y(N185) );
  ivd1_hd U108 ( .A(n9), .Y(N174) );
  or2d1_hd U109 ( .A(n7), .B(N183), .Y(N184) );
  or2d1_hd U110 ( .A(n36), .B(N182), .Y(N183) );
  or2d1_hd U111 ( .A(n8), .B(N168), .Y(N169) );
  or2d1_hd U112 ( .A(n7), .B(N167), .Y(N168) );
  or2d1_hd U113 ( .A(n36), .B(N166), .Y(N167) );
  or2d1_hd U114 ( .A(n35), .B(N165), .Y(N166) );
  ivd1_hd U115 ( .A(n11), .Y(N158) );
  or2d1_hd U116 ( .A(N175), .B(N187), .Y(N188) );
  ivd1_hd U117 ( .A(n16), .Y(N175) );
  or2d1_hd U118 ( .A(n13), .B(N186), .Y(N187) );
  or2d1_hd U119 ( .A(N158), .B(N185), .Y(N186) );
  or2d1_hd U120 ( .A(N159), .B(N170), .Y(N171) );
  ivd1_hd U121 ( .A(n14), .Y(N159) );
  or2d1_hd U122 ( .A(N158), .B(N169), .Y(N170) );
  clknd2d1_hd U123 ( .A(n63), .B(N31), .Y(n66) );
  clknd2d1_hd U124 ( .A(n69), .B(n68), .Y(n72) );
  clknd2d1_hd U125 ( .A(n75), .B(n74), .Y(n78) );
  or2d1_hd U126 ( .A(N189), .B(N173), .Y(N75) );
  clknd2d1_hd U127 ( .A(N110), .B(N173), .Y(n31) );
  clknd2d1_hd U128 ( .A(N110), .B(N189), .Y(n30) );
  clknd2d1_hd U129 ( .A(n83), .B(n82), .Y(N26) );
  ad2d1_hd U130 ( .A(N134), .B(alt9_n41), .Y(N154) );
  or2d1_hd U131 ( .A(o_TX_Ready), .B(N154), .Y(N144) );
  ad2d1_hd U132 ( .A(N116), .B(alt9_n41), .Y(N126) );
  clknd2d1_hd U133 ( .A(alt9_n41), .B(n27), .Y(N125) );
  ivd1_hd U134 ( .A(N126), .Y(n27) );
  mx2d1_hd U135 ( .D0(n84), .D1(N100), .S(N99), .Y(r_SPI_Clk_Edges[0]) );
  mx2d1_hd U136 ( .D0(n61), .D1(N101), .S(N99), .Y(r_SPI_Clk_Edges[1]) );
  mx2d1_hd U137 ( .D0(n59), .D1(N102), .S(N99), .Y(r_SPI_Clk_Edges[2]) );
  mx2d1_hd U138 ( .D0(n58), .D1(N103), .S(N99), .Y(r_SPI_Clk_Edges[3]) );
  mx2d1_hd U139 ( .D0(n57), .D1(N104), .S(N99), .Y(r_SPI_Clk_Edges[4]) );
  mx2d1_hd U140 ( .D0(n56), .D1(N105), .S(N99), .Y(r_SPI_Clk_Edges[5]) );
  mx2d1_hd U141 ( .D0(n55), .D1(N106), .S(N99), .Y(r_SPI_Clk_Edges[6]) );
  mx2d1_hd U142 ( .D0(n54), .D1(N107), .S(N99), .Y(r_SPI_Clk_Edges[7]) );
  xo2d1_hd U143 ( .A(n54), .B(n79), .Y(N38) );
  mx2d1_hd U152 ( .D0(o_SPI_Clk), .D1(N23), .S(n60), .Y(r_SPI_Clk) );
  ivd1_hd U153 ( .A(o_SPI_Clk), .Y(N23) );
  mx2d1_hd U162 ( .D0(o_RX_Byte[0]), .D1(i_SPI_MISO), .S(N145), .Y(n97) );
  ad2d1_hd U163 ( .A(N207), .B(N11), .Y(N208) );
  ad2d1_hd U164 ( .A(N0), .B(N1), .Y(N207) );
  mx2d1_hd U165 ( .D0(o_RX_Byte[1]), .D1(i_SPI_MISO), .S(N146), .Y(n96) );
  ad2d1_hd U166 ( .A(N205), .B(N11), .Y(N206) );
  ad2d1_hd U167 ( .A(n40), .B(N1), .Y(N205) );
  mx2d1_hd U168 ( .D0(o_RX_Byte[2]), .D1(i_SPI_MISO), .S(N147), .Y(n95) );
  ad2d1_hd U169 ( .A(N203), .B(N11), .Y(N204) );
  ad2d1_hd U170 ( .A(N0), .B(n41), .Y(N203) );
  mx2d1_hd U171 ( .D0(o_RX_Byte[3]), .D1(i_SPI_MISO), .S(N148), .Y(n94) );
  ad2d1_hd U172 ( .A(N201), .B(N11), .Y(N202) );
  ad2d1_hd U173 ( .A(n40), .B(n41), .Y(N201) );
  mx2d1_hd U174 ( .D0(o_RX_Byte[4]), .D1(i_SPI_MISO), .S(N149), .Y(n93) );
  ad2d1_hd U175 ( .A(N199), .B(n42), .Y(N200) );
  ad2d1_hd U176 ( .A(N0), .B(N1), .Y(N199) );
  mx2d1_hd U177 ( .D0(o_RX_Byte[5]), .D1(i_SPI_MISO), .S(N150), .Y(n92) );
  ad2d1_hd U178 ( .A(N197), .B(n42), .Y(N198) );
  ad2d1_hd U179 ( .A(n40), .B(N1), .Y(N197) );
  mx2d1_hd U180 ( .D0(o_RX_Byte[6]), .D1(i_SPI_MISO), .S(N151), .Y(n91) );
  ad2d1_hd U181 ( .A(N195), .B(n42), .Y(N196) );
  ad2d1_hd U182 ( .A(N0), .B(n41), .Y(N195) );
  mx2d1_hd U183 ( .D0(o_RX_Byte[7]), .D1(i_SPI_MISO), .S(N152), .Y(n90) );
  ad2d1_hd U184 ( .A(N193), .B(n42), .Y(N194) );
  ad2d1_hd U185 ( .A(n40), .B(n41), .Y(N193) );
  or2d1_hd U186 ( .A(n41), .B(n42), .Y(N155) );
  mx2d1_hd U187 ( .D0(o_SPI_MOSI), .D1(N127), .S(N126), .Y(n98) );
  mx2d1_hd U188 ( .D0(n80), .D1(n81), .S(n39), .Y(N121) );
  mx2d1_hd U189 ( .D0(n42), .D1(N143), .S(N144), .Y(r_RX_Bit_Count[2]) );
  xn2d1_hd U190 ( .A(sub_x_13_n1), .B(n42), .Y(N140) );
  or2d1_hd U191 ( .A(n40), .B(n41), .Y(sub_x_13_n1) );
  mx2d1_hd U192 ( .D0(n41), .D1(N142), .S(N144), .Y(r_RX_Bit_Count[1]) );
  xn2d1_hd U193 ( .A(n40), .B(n41), .Y(N139) );
  mx2d1_hd U194 ( .D0(n40), .D1(N141), .S(N144), .Y(r_RX_Bit_Count[0]) );
  mx2d1_hd U195 ( .D0(n39), .D1(N124), .S(N125), .Y(r_TX_Bit_Count[2]) );
  xn2d1_hd U196 ( .A(sub_x_11_n1), .B(n39), .Y(N120) );
  or2d1_hd U197 ( .A(n37), .B(n38), .Y(sub_x_11_n1) );
  mx2d1_hd U198 ( .D0(n38), .D1(N123), .S(N125), .Y(r_TX_Bit_Count[1]) );
  xn2d1_hd U199 ( .A(n37), .B(n38), .Y(N119) );
  mx2d1_hd U200 ( .D0(n37), .D1(N122), .S(N125), .Y(r_TX_Bit_Count[0]) );
  scg2d1_hd U202 ( .A(N47), .B(n2), .C(n15), .D(n3), .Y(r_SPI_Clk_Count[0]) );
  scg2d1_hd U203 ( .A(N48), .B(n2), .C(n13), .D(n3), .Y(r_SPI_Clk_Count[1]) );
  scg2d1_hd U205 ( .A(N49), .B(n2), .C(n10), .D(n3), .Y(r_SPI_Clk_Count[2]) );
  scg2d1_hd U206 ( .A(N50), .B(n2), .C(n8), .D(n3), .Y(r_SPI_Clk_Count[3]) );
  ad2d1_hd U209 ( .A(N75), .B(N110), .Y(n60) );
  nr2d1_hd U210 ( .A(N26), .B(n86), .Y(o_TX_Ready) );
  ivd1_hd U212 ( .A(n40), .Y(N0) );
  nr2d1_hd U214 ( .A(n40), .B(N155), .Y(n62) );
  ivd1_hd U215 ( .A(o_TX_Ready), .Y(alt9_n41) );
  ivd1_hd U216 ( .A(n84), .Y(N31) );
  ivd1_hd U217 ( .A(n61), .Y(n63) );
  ao22d1_hd U218 ( .A(n61), .B(N31), .C(n84), .D(n63), .Y(N32) );
  ivd1_hd U219 ( .A(n66), .Y(n65) );
  ivd1_hd U220 ( .A(n59), .Y(n64) );
  ao22d1_hd U221 ( .A(n59), .B(n65), .C(n66), .D(n64), .Y(N33) );
  nr2d1_hd U222 ( .A(n59), .B(n66), .Y(n69) );
  ivd1_hd U223 ( .A(n69), .Y(n67) );
  ivd1_hd U224 ( .A(n58), .Y(n68) );
  ao22d1_hd U225 ( .A(n58), .B(n69), .C(n67), .D(n68), .Y(N34) );
  ivd1_hd U226 ( .A(n72), .Y(n71) );
  ivd1_hd U227 ( .A(n57), .Y(n70) );
  ao22d1_hd U228 ( .A(n57), .B(n71), .C(n72), .D(n70), .Y(N35) );
  nr2d1_hd U229 ( .A(n57), .B(n72), .Y(n75) );
  ivd1_hd U230 ( .A(n75), .Y(n73) );
  ivd1_hd U231 ( .A(n56), .Y(n74) );
  ao22d1_hd U232 ( .A(n56), .B(n75), .C(n73), .D(n74), .Y(N36) );
  ivd1_hd U233 ( .A(n78), .Y(n77) );
  ivd1_hd U234 ( .A(n55), .Y(n76) );
  ao22d1_hd U235 ( .A(n55), .B(n77), .C(n78), .D(n76), .Y(N37) );
  nr2d1_hd U236 ( .A(n55), .B(n78), .Y(n79) );
  mx4d1_hd U237 ( .D0(n24), .D1(n23), .D2(n22), .D3(n21), .S0(n37), .S1(n38), 
        .Y(n80) );
  mx4d1_hd U238 ( .D0(n20), .D1(n19), .D2(n18), .D3(n17), .S0(n37), .S1(n38), 
        .Y(n81) );
  nr4d1_hd U239 ( .A(n58), .B(n59), .C(n61), .D(n84), .Y(n83) );
  nr4d1_hd U240 ( .A(n53), .B(n55), .C(n56), .D(n57), .Y(n82) );
  fd3qd1_hd clk_r_REG10_S1 ( .D(n1), .CK(i_CLK), .SN(n6), .Q(n88) );
  fd3qd1_hd clk_r_REG14_S2 ( .D(r_SPI_Clk_Edges[7]), .CK(i_CLK), .SN(n6), .Q(
        n53) );
  fd3qd1_hd clk_r_REG27_S3 ( .D(r_RX_Bit_Count[0]), .CK(n134), .SN(n99), .Q(
        n40) );
  fd3qd1_hd clk_r_REG11_S2 ( .D(r_TX_Bit_Count[2]), .CK(n134), .SN(n99), .Q(
        n39) );
  fd3qd1_hd clk_r_REG12_S2 ( .D(r_TX_Bit_Count[1]), .CK(n134), .SN(n99), .Q(
        n38) );
  fd3qd1_hd clk_r_REG13_S2 ( .D(r_TX_Bit_Count[0]), .CK(n134), .SN(n99), .Q(
        n37) );
  fd3qd1_hd clk_r_REG36_S2 ( .D(n146), .CK(n132), .SN(n6), .Q(n36) );
  fd3qd1_hd clk_r_REG37_S2 ( .D(n147), .CK(n132), .SN(n6), .Q(n35) );
  fd3qd1_hd clk_r_REG38_S2 ( .D(n148), .CK(n132), .SN(n6), .Q(n34) );
  fd3qd1_hd clk_r_REG39_S2 ( .D(n149), .CK(n132), .SN(n6), .Q(n33) );
  fd3qd1_hd clk_r_REG40_S2 ( .D(n150), .CK(n132), .SN(n6), .Q(n29) );
  fd3qd1_hd clk_r_REG41_S2 ( .D(n151), .CK(n132), .SN(n6), .Q(n28) );
  fd3qd1_hd clk_r_REG42_S2 ( .D(n152), .CK(n132), .SN(n6), .Q(n26) );
  fd3qd1_hd clk_r_REG43_S2 ( .D(n153), .CK(n132), .SN(n6), .Q(n25) );
  fd3qd1_hd clk_r_REG45_S2 ( .D(n154), .CK(n132), .SN(n6), .Q(n15) );
  fd3qd1_hd clk_r_REG47_S2 ( .D(r_SPI_Clk_Count[1]), .CK(n132), .SN(n6), .Q(
        n13) );
  fd3qd1_hd clk_r_REG44_S2 ( .D(n155), .CK(n132), .SN(n6), .Q(n12) );
  fd3qd1_hd clk_r_REG49_S2 ( .D(n156), .CK(n132), .SN(n6), .Q(n10) );
  fd3qd1_hd clk_r_REG51_S2 ( .D(n157), .CK(n132), .SN(n6), .Q(n8) );
  fd3qd1_hd clk_r_REG53_S2 ( .D(n158), .CK(n132), .SN(n6), .Q(n7) );
  fd3d1_hd clk_r_REG26_S3 ( .D(r_RX_Bit_Count[1]), .CK(n134), .SN(n99), .Q(n41), .QN(N1) );
  fd3d1_hd clk_r_REG16_S3 ( .D(r_RX_Bit_Count[2]), .CK(n134), .SN(n99), .Q(n42), .QN(N11) );
  clknd2d1_hd U1 ( .A(N26), .B(n88), .Y(n3) );
  ivd1_hd U2 ( .A(n87), .Y(n99) );
  ivd2_hd U3 ( .A(n87), .Y(n6) );
  ivd1_hd U4 ( .A(w_rstn), .Y(n87) );
  spi_master_DW01_inc_0 add_x_3 ( .A({n12, n25, n26, n28, n29, n33, n34, n35, 
        n36, n7, n8, n10, n13, n15}), .SUM({N60, N59, N58, N57, N56, N55, N54, 
        N53, N52, N51, N50, N49, N48, N47}) );
  SNPS_CLOCK_GATE_HIGH_spi_master_3 clk_gate_clk_r_REG34_S2_0 ( .CLK(i_CLK), 
        .EN(n144), .ENCLK(n134), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_spi_master_4 clk_gate_clk_r_REG0_S1_0 ( .CLK(i_CLK), 
        .EN(i_TX_DV), .ENCLK(n133), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_spi_master_5 clk_gate_clk_r_REG53_S2_0 ( .CLK(i_CLK), 
        .EN(N110), .ENCLK(n132), .TE(1'b0) );
  fd4qd1_hd clk_r_REG8_S1 ( .D(i_TX_Byte[0]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n24) );
  fd4qd1_hd clk_r_REG7_S1 ( .D(i_TX_Byte[1]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n23) );
  fd4qd1_hd clk_r_REG6_S1 ( .D(i_TX_Byte[2]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n22) );
  fd4qd1_hd clk_r_REG5_S1 ( .D(i_TX_Byte[3]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n21) );
  fd4qd1_hd clk_r_REG4_S1 ( .D(i_TX_Byte[4]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n20) );
  fd4qd1_hd clk_r_REG3_S1 ( .D(i_TX_Byte[5]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n19) );
  fd4qd1_hd clk_r_REG2_S1 ( .D(i_TX_Byte[6]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n18) );
  fd4qd1_hd clk_r_REG0_S1 ( .D(i_TX_Byte[7]), .CK(n133), .SN(1'b1), .RN(w_rstn), .Q(n17) );
  fd4qd1_hd clk_r_REG9_S1 ( .D(i_TX_DV), .CK(i_CLK), .SN(1'b1), .RN(n6), .Q(
        n86) );
  fd4qd1_hd clk_r_REG52_S2 ( .D(r_SPI_Clk_Count[3]), .CK(i_CLK), .SN(1'b1), 
        .RN(n6), .Q(n9) );
  fd4qd1_hd clk_r_REG50_S2 ( .D(r_SPI_Clk_Count[2]), .CK(i_CLK), .SN(1'b1), 
        .RN(n6), .Q(n11) );
  fd4qd1_hd clk_r_REG46_S2 ( .D(r_SPI_Clk_Count[0]), .CK(i_CLK), .SN(1'b1), 
        .RN(n6), .Q(n16) );
  fd4qd1_hd clk_r_REG48_S2 ( .D(r_SPI_Clk_Count[1]), .CK(i_CLK), .SN(1'b1), 
        .RN(n6), .Q(n14) );
  fd4qd1_hd clk_r_REG35_S2 ( .D(r_SPI_Clk), .CK(n132), .SN(1'b1), .RN(n6), .Q(
        o_SPI_Clk) );
  fd4qd1_hd clk_r_REG21_S4 ( .D(n89), .CK(i_CLK), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_DV) );
  fd4qd1_hd clk_r_REG25_S4 ( .D(n94), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[3]) );
  fd4qd1_hd clk_r_REG24_S4 ( .D(n95), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[2]) );
  fd4qd1_hd clk_r_REG23_S4 ( .D(n96), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[1]) );
  fd4qd1_hd clk_r_REG22_S4 ( .D(n97), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[0]) );
  fd4qd1_hd clk_r_REG20_S4 ( .D(n90), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[7]) );
  fd4qd1_hd clk_r_REG19_S4 ( .D(n91), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[6]) );
  fd4qd1_hd clk_r_REG18_S4 ( .D(n92), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[5]) );
  fd4qd1_hd clk_r_REG17_S4 ( .D(n93), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_RX_Byte[4]) );
  fd4qd1_hd clk_r_REG1_S2 ( .D(n98), .CK(n132), .SN(1'b1), .RN(w_rstn), .Q(
        o_SPI_MOSI) );
  fd4qd1_hd clk_r_REG34_S2 ( .D(r_SPI_Clk_Edges[0]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n84) );
  fd4qd1_hd clk_r_REG33_S2 ( .D(r_SPI_Clk_Edges[1]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n61) );
  fd4qd1_hd clk_r_REG32_S2 ( .D(r_SPI_Clk_Edges[2]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n59) );
  fd4qd1_hd clk_r_REG31_S2 ( .D(r_SPI_Clk_Edges[3]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n58) );
  fd4qd1_hd clk_r_REG30_S2 ( .D(r_SPI_Clk_Edges[4]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n57) );
  fd4qd1_hd clk_r_REG29_S2 ( .D(r_SPI_Clk_Edges[5]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n56) );
  fd4qd1_hd clk_r_REG28_S2 ( .D(r_SPI_Clk_Edges[6]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n55) );
  fd4qd1_hd clk_r_REG15_S2 ( .D(r_SPI_Clk_Edges[7]), .CK(n134), .SN(1'b1), 
        .RN(n6), .Q(n54) );
  scg20d1_hd U5 ( .A(N173), .B(N188), .C(n3), .Y(n2) );
  nr2ad1_hd U6 ( .A(n15), .B(N171), .Y(N173) );
  scg17d1_hd U69 ( .A(n135), .B(n136), .C(n86), .D(n137), .Y(n144) );
  nd3d1_hd U70 ( .A(n138), .B(n139), .C(n140), .Y(n137) );
  nr4d1_hd U71 ( .A(n35), .B(n7), .C(N158), .D(n141), .Y(n140) );
  ivd1_hd U72 ( .A(n88), .Y(n141) );
  nr4d1_hd U73 ( .A(n28), .B(n29), .C(n36), .D(n34), .Y(n139) );
  nr4d1_hd U74 ( .A(n26), .B(n12), .C(n25), .D(n33), .Y(n138) );
  nr4d1_hd U75 ( .A(n57), .B(n56), .C(n55), .D(n53), .Y(n136) );
  nr4d1_hd U76 ( .A(n84), .B(n61), .C(n59), .D(n58), .Y(n135) );
  scg9d1_hd U77 ( .A(N173), .B(N188), .C(N52), .Y(n146) );
  scg9d1_hd U78 ( .A(N173), .B(N188), .C(N53), .Y(n147) );
  scg9d1_hd U79 ( .A(N173), .B(N188), .C(N54), .Y(n148) );
  scg9d1_hd U80 ( .A(N173), .B(N188), .C(N55), .Y(n149) );
  scg9d1_hd U81 ( .A(N173), .B(N188), .C(N56), .Y(n150) );
  scg9d1_hd U82 ( .A(N173), .B(N188), .C(N57), .Y(n151) );
  scg9d1_hd U83 ( .A(N173), .B(N188), .C(N58), .Y(n152) );
  scg9d1_hd U84 ( .A(N173), .B(N188), .C(N59), .Y(n153) );
  scg9d1_hd U85 ( .A(n142), .B(N188), .C(N47), .Y(n154) );
  nr2d1_hd U86 ( .A(n15), .B(N171), .Y(n142) );
  scg9d1_hd U87 ( .A(N173), .B(N188), .C(N60), .Y(n155) );
  scg9d1_hd U88 ( .A(N173), .B(N188), .C(N49), .Y(n156) );
  scg9d1_hd U89 ( .A(N173), .B(N188), .C(N50), .Y(n157) );
  scg9d1_hd U90 ( .A(N173), .B(N188), .C(N51), .Y(n158) );
endmodule


module ads1292_controller_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  had1_hd U2 ( .A(A[30]), .B(n2), .CO(n1), .S(SUM[30]) );
  had1_hd U3 ( .A(A[29]), .B(n3), .CO(n2), .S(SUM[29]) );
  had1_hd U4 ( .A(A[28]), .B(n4), .CO(n3), .S(SUM[28]) );
  had1_hd U5 ( .A(A[27]), .B(n5), .CO(n4), .S(SUM[27]) );
  had1_hd U6 ( .A(A[26]), .B(n6), .CO(n5), .S(SUM[26]) );
  had1_hd U7 ( .A(A[25]), .B(n7), .CO(n6), .S(SUM[25]) );
  had1_hd U8 ( .A(A[24]), .B(n8), .CO(n7), .S(SUM[24]) );
  had1_hd U9 ( .A(A[23]), .B(n9), .CO(n8), .S(SUM[23]) );
  had1_hd U10 ( .A(A[22]), .B(n10), .CO(n9), .S(SUM[22]) );
  had1_hd U11 ( .A(A[21]), .B(n11), .CO(n10), .S(SUM[21]) );
  had1_hd U12 ( .A(A[20]), .B(n12), .CO(n11), .S(SUM[20]) );
  had1_hd U13 ( .A(A[19]), .B(n13), .CO(n12), .S(SUM[19]) );
  had1_hd U14 ( .A(A[18]), .B(n14), .CO(n13), .S(SUM[18]) );
  had1_hd U15 ( .A(A[17]), .B(n15), .CO(n14), .S(SUM[17]) );
  had1_hd U16 ( .A(A[16]), .B(n16), .CO(n15), .S(SUM[16]) );
  had1_hd U17 ( .A(A[15]), .B(n17), .CO(n16), .S(SUM[15]) );
  had1_hd U18 ( .A(A[14]), .B(n18), .CO(n17), .S(SUM[14]) );
  had1_hd U19 ( .A(A[13]), .B(n19), .CO(n18), .S(SUM[13]) );
  had1_hd U20 ( .A(A[12]), .B(n20), .CO(n19), .S(SUM[12]) );
  had1_hd U21 ( .A(A[11]), .B(n21), .CO(n20), .S(SUM[11]) );
  had1_hd U22 ( .A(A[10]), .B(n22), .CO(n21), .S(SUM[10]) );
  had1_hd U23 ( .A(A[9]), .B(n23), .CO(n22), .S(SUM[9]) );
  had1_hd U24 ( .A(A[8]), .B(n24), .CO(n23), .S(SUM[8]) );
  had1_hd U25 ( .A(A[7]), .B(n25), .CO(n24), .S(SUM[7]) );
  had1_hd U26 ( .A(A[6]), .B(n26), .CO(n25), .S(SUM[6]) );
  had1_hd U27 ( .A(A[5]), .B(n27), .CO(n26), .S(SUM[5]) );
  had1_hd U28 ( .A(A[4]), .B(n28), .CO(n27), .S(SUM[4]) );
  had1_hd U29 ( .A(A[3]), .B(n29), .CO(n28), .S(SUM[3]) );
  had1_hd U30 ( .A(A[2]), .B(n30), .CO(n29), .S(SUM[2]) );
  had1_hd U31 ( .A(A[1]), .B(A[0]), .CO(n30), .S(SUM[1]) );
  xo2d1_hd U35 ( .A(n1), .B(A[31]), .Y(SUM[31]) );
  ivd1_hd U36 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ads1292_controller_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  cglpd1_hd latch ( .EN(EN), .CK(CLK), .TE(TE), .GCK(ENCLK) );
endmodule


module ads1292_controller ( o_ADS1292_DATA_OUT, i_ADS1292_CONTROL, 
        i_ADS1292_REG_ADDR, i_ADS1292_DATA_IN, o_ADS1292_REG_DATA_OUT, 
        o_ADS1292_INIT_SET, o_ADS1292_DATA_VALID, o_ADS1292_BUSY, o_SPI_CLK, 
        i_SPI_MISO, o_SPI_MOSI, i_ADS1292_DRDY, o_ADS1292_RESET, 
        o_ADS1292_START, o_SPI_CSN, i_CLK, i_RSTN );
  output [23:0] o_ADS1292_DATA_OUT;
  input [2:0] i_ADS1292_CONTROL;
  input [7:0] i_ADS1292_REG_ADDR;
  input [7:0] i_ADS1292_DATA_IN;
  output [7:0] o_ADS1292_REG_DATA_OUT;
  input i_SPI_MISO, i_ADS1292_DRDY, i_CLK, i_RSTN;
  output o_ADS1292_INIT_SET, o_ADS1292_DATA_VALID, o_ADS1292_BUSY, o_SPI_CLK,
         o_SPI_MOSI, o_ADS1292_RESET, o_ADS1292_START, o_SPI_CSN;
  wire   n161, n162, n163, n164, n165, n166, w_rstn, r_spi_data_in_valid,
         w_spi_data_in_ready, w_spi_data_out_valid, N331, N332, N333, N334,
         N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345,
         N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N942, N983, N984, N985, N1171,
         n248, n253, n261, n262, n263, n265, n266, n267, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n322, n325, n326, n327, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, r_drdy_edge_counter_1_, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n24, n25, n26, n27, n28, n29, n30, n32,
         n33, n34, n35, n36, n37, n39, n41, n43, n45, n48, n50, n52, n54, n56,
         n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n82, n84,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n149, n150, n159, n160, n167, n168, n170,
         n171, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n588, n590, n591, n592, n593, n594, n595, n596,
         n597, n599, n600;
  wire   [7:0] w_spi_data_out;
  wire   [6:0] r_pstate;
  wire   [31:0] r_clk_counter;
  wire   [4:0] r_lstate;
  wire   [3:0] r_data_counter;

  async_rstn_synchronizer async_rstn_synchronizer ( .i_CLK(i_CLK), .i_RSTN(
        i_RSTN), .o_RSTN(w_rstn) );
  spi_master spi_master ( .i_RSTN(w_rstn), .i_CLK(i_CLK), .i_TX_Byte({n25, n87, 
        n88, n89, n90, n91, n92, n93}), .i_TX_DV(n24), .o_TX_Ready(
        w_spi_data_in_ready), .o_RX_DV(w_spi_data_out_valid), .o_RX_Byte(
        w_spi_data_out), .o_SPI_Clk(o_SPI_CLK), .i_SPI_MISO(i_SPI_MISO), 
        .o_SPI_MOSI(o_SPI_MOSI) );
  clknd2d1_hd U322 ( .A(n454), .B(n361), .Y(n333) );
  clknd2d1_hd U323 ( .A(n552), .B(n551), .Y(n547) );
  clknd2d1_hd U324 ( .A(n552), .B(n545), .Y(n394) );
  clknd2d1_hd U325 ( .A(n487), .B(n518), .Y(n273) );
  clknd2d1_hd U326 ( .A(n504), .B(n505), .Y(n272) );
  clknd2d1_hd U327 ( .A(n109), .B(n110), .Y(n508) );
  clknd2d1_hd U328 ( .A(n469), .B(n470), .Y(n457) );
  clknd2d1_hd U329 ( .A(n32), .B(n104), .Y(n296) );
  clknd2d1_hd U330 ( .A(n149), .B(n410), .Y(n546) );
  clknd2d1_hd U331 ( .A(n519), .B(n483), .Y(n285) );
  clknd2d1_hd U332 ( .A(n360), .B(n483), .Y(n358) );
  clknd2d1_hd U333 ( .A(n358), .B(n319), .Y(n366) );
  clknd2d1_hd U334 ( .A(n363), .B(n451), .Y(n368) );
  clknd2d1_hd U335 ( .A(n16), .B(n449), .Y(n455) );
  clknd2d1_hd U336 ( .A(n20), .B(n363), .Y(n499) );
  clknd2d1_hd U337 ( .A(n394), .B(n332), .Y(n407) );
  clknd2d1_hd U338 ( .A(n20), .B(n558), .Y(n500) );
  clknd2d1_hd U339 ( .A(n558), .B(n518), .Y(n340) );
  clknd2d1_hd U340 ( .A(n20), .B(n555), .Y(n541) );
  clknd2d1_hd U341 ( .A(n19), .B(n544), .Y(n542) );
  clknd2d1_hd U342 ( .A(n403), .B(n518), .Y(n478) );
  clknd2d1_hd U343 ( .A(n29), .B(n315), .Y(n307) );
  clknd2d1_hd U344 ( .A(n317), .B(n310), .Y(n311) );
  clknd2d1_hd U345 ( .A(n281), .B(n335), .Y(n334) );
  clknd2d1_hd U346 ( .A(n20), .B(n519), .Y(n423) );
  clknd2d1_hd U347 ( .A(n300), .B(n457), .Y(n419) );
  clknd2d1_hd U348 ( .A(n461), .B(n414), .Y(n424) );
  clknd2d1_hd U349 ( .A(n18), .B(n454), .Y(n322) );
  clknd2d1_hd U350 ( .A(n448), .B(n360), .Y(n447) );
  clknd2d1_hd U352 ( .A(n448), .B(n451), .Y(n486) );
  clknd2d1_hd U354 ( .A(n267), .B(i_ADS1292_REG_ADDR[3]), .Y(n269) );
  clknd2d1_hd U355 ( .A(n428), .B(n160), .Y(n383) );
  ivd1_hd U356 ( .A(n267), .Y(n265) );
  clknd2d1_hd U358 ( .A(n308), .B(n368), .Y(n465) );
  clknd2d1_hd U359 ( .A(n15), .B(n360), .Y(n434) );
  clknd2d1_hd U360 ( .A(n296), .B(n294), .Y(n291) );
  clknd2d1_hd U362 ( .A(n363), .B(n536), .Y(n319) );
  clknd2d1_hd U363 ( .A(n536), .B(n448), .Y(n406) );
  clknd2d1_hd U364 ( .A(n15), .B(n519), .Y(n556) );
  clknd2d1_hd U365 ( .A(n373), .B(n557), .Y(n498) );
  clknd2d1_hd U366 ( .A(n19), .B(n518), .Y(n540) );
  clknd2d1_hd U367 ( .A(n286), .B(n131), .Y(n320) );
  clknd2d1_hd U368 ( .A(n536), .B(n361), .Y(n350) );
  clknd2d1_hd U369 ( .A(n265), .B(n478), .Y(n304) );
  scg2d1_hd U370 ( .A(n141), .B(n270), .C(N362), .D(n271), .Y(
        r_clk_counter[31]) );
  scg2d1_hd U371 ( .A(n140), .B(n270), .C(N361), .D(n271), .Y(
        r_clk_counter[30]) );
  scg2d1_hd U372 ( .A(n139), .B(n270), .C(N360), .D(n271), .Y(
        r_clk_counter[29]) );
  scg2d1_hd U373 ( .A(n138), .B(n270), .C(N359), .D(n271), .Y(
        r_clk_counter[28]) );
  scg2d1_hd U374 ( .A(n137), .B(n270), .C(N358), .D(n271), .Y(
        r_clk_counter[27]) );
  scg2d1_hd U375 ( .A(n136), .B(n270), .C(N357), .D(n271), .Y(
        r_clk_counter[26]) );
  scg2d1_hd U376 ( .A(n135), .B(n270), .C(N356), .D(n271), .Y(
        r_clk_counter[25]) );
  scg2d1_hd U377 ( .A(n134), .B(n270), .C(N355), .D(n271), .Y(
        r_clk_counter[24]) );
  scg2d1_hd U378 ( .A(n133), .B(n270), .C(N354), .D(n271), .Y(
        r_clk_counter[23]) );
  scg2d1_hd U379 ( .A(n132), .B(n270), .C(N353), .D(n271), .Y(
        r_clk_counter[22]) );
  scg2d1_hd U380 ( .A(n131), .B(n305), .C(n306), .D(n28), .Y(r_data_counter[3]) );
  scg2d1_hd U381 ( .A(n130), .B(n270), .C(N352), .D(n271), .Y(
        r_clk_counter[21]) );
  scg2d1_hd U382 ( .A(n129), .B(n270), .C(N351), .D(n271), .Y(
        r_clk_counter[20]) );
  scg2d1_hd U383 ( .A(n128), .B(n270), .C(N331), .D(n271), .Y(r_clk_counter[0]) );
  scg2d1_hd U384 ( .A(n127), .B(n270), .C(N332), .D(n271), .Y(r_clk_counter[1]) );
  scg2d1_hd U385 ( .A(n126), .B(n270), .C(N333), .D(n271), .Y(r_clk_counter[2]) );
  scg2d1_hd U386 ( .A(n125), .B(n270), .C(N334), .D(n271), .Y(r_clk_counter[3]) );
  scg2d1_hd U387 ( .A(n124), .B(n270), .C(N335), .D(n271), .Y(r_clk_counter[4]) );
  scg2d1_hd U388 ( .A(n123), .B(n270), .C(N336), .D(n271), .Y(r_clk_counter[5]) );
  scg2d1_hd U389 ( .A(n122), .B(n270), .C(N337), .D(n271), .Y(r_clk_counter[6]) );
  scg2d1_hd U390 ( .A(n121), .B(n270), .C(N338), .D(n271), .Y(r_clk_counter[7]) );
  scg2d1_hd U391 ( .A(n120), .B(n270), .C(N339), .D(n271), .Y(r_clk_counter[8]) );
  scg2d1_hd U392 ( .A(n119), .B(n270), .C(N340), .D(n271), .Y(r_clk_counter[9]) );
  scg2d1_hd U393 ( .A(n118), .B(n270), .C(N341), .D(n271), .Y(
        r_clk_counter[10]) );
  scg2d1_hd U394 ( .A(n117), .B(n270), .C(N342), .D(n271), .Y(
        r_clk_counter[11]) );
  scg2d1_hd U395 ( .A(n116), .B(n270), .C(N343), .D(n271), .Y(
        r_clk_counter[12]) );
  scg2d1_hd U396 ( .A(n115), .B(n270), .C(N344), .D(n271), .Y(
        r_clk_counter[13]) );
  scg2d1_hd U397 ( .A(n114), .B(n270), .C(N345), .D(n271), .Y(
        r_clk_counter[14]) );
  scg2d1_hd U398 ( .A(n113), .B(n270), .C(N346), .D(n271), .Y(
        r_clk_counter[15]) );
  scg2d1_hd U399 ( .A(n112), .B(n270), .C(N347), .D(n271), .Y(
        r_clk_counter[16]) );
  scg2d1_hd U400 ( .A(n111), .B(n270), .C(N348), .D(n271), .Y(
        r_clk_counter[17]) );
  scg2d1_hd U401 ( .A(n110), .B(n270), .C(N349), .D(n271), .Y(
        r_clk_counter[18]) );
  scg2d1_hd U402 ( .A(n109), .B(n270), .C(N350), .D(n271), .Y(
        r_clk_counter[19]) );
  scg2d1_hd U408 ( .A(n32), .B(n289), .C(n104), .D(n290), .Y(
        r_drdy_edge_counter_1_) );
  clknd2d1_hd U409 ( .A(n291), .B(n288), .Y(n290) );
  clknd2d1_hd U410 ( .A(o_ADS1292_START), .B(n319), .Y(n388) );
  clknd2d1_hd U421 ( .A(n382), .B(o_ADS1292_BUSY), .Y(n381) );
  clknd2d1_hd U452 ( .A(n369), .B(n371), .Y(n370) );
  scg2d1_hd U453 ( .A(n395), .B(n396), .C(o_ADS1292_INIT_SET), .D(n319), .Y(
        n161) );
  clknd2d1_hd U454 ( .A(n422), .B(n556), .Y(r_lstate[1]) );
  clknd2d1_hd U455 ( .A(n553), .B(n329), .Y(N1171) );
  mx2d1_hd U457 ( .D0(n282), .D1(o_ADS1292_RESET), .S(n336), .Y(n164) );
  clknd2d1_hd U458 ( .A(n297), .B(o_SPI_CSN), .Y(n299) );
  clknd2d1_hd U465 ( .A(n267), .B(n160), .Y(n433) );
  clknd2d1_hd U466 ( .A(n267), .B(i_ADS1292_REG_ADDR[0]), .Y(n266) );
  oa211d4_hd U468 ( .A(n272), .B(n273), .C(n274), .D(n275), .Y(n271) );
  nr4d6_hd U469 ( .A(n280), .B(n281), .C(n282), .D(n283), .Y(n270) );
  clknd2d1_hd U470 ( .A(n284), .B(n285), .Y(n283) );
  ivd1_hd U509 ( .A(n35), .Y(n248) );
  ivd1_hd U522 ( .A(i_ADS1292_CONTROL[1]), .Y(n262) );
  ivd1_hd U523 ( .A(i_ADS1292_CONTROL[2]), .Y(n261) );
  ivd1_hd U525 ( .A(i_ADS1292_CONTROL[0]), .Y(n253) );
  ao211d1_hd U529 ( .A(n276), .B(n277), .C(n278), .D(n279), .Y(n275) );
  nr2d1_hd U531 ( .A(n292), .B(n291), .Y(n289) );
  ivd1_hd U532 ( .A(n292), .Y(n288) );
  ao21d1_hd U533 ( .A(n293), .B(n294), .C(n295), .Y(n292) );
  scg16d1_hd U534 ( .A(n159), .B(i_ADS1292_DRDY), .C(n296), .Y(n293) );
  oa211d1_hd U535 ( .A(n297), .B(n284), .C(n298), .D(n299), .Y(n166) );
  nr2d1_hd U536 ( .A(n300), .B(n301), .Y(n284) );
  ao211d1_hd U537 ( .A(n301), .B(n302), .C(n303), .D(n304), .Y(n297) );
  nr2d1_hd U538 ( .A(n131), .B(n307), .Y(n306) );
  oa21d1_hd U539 ( .A(n308), .B(n28), .C(n309), .Y(n305) );
  ao22d1_hd U540 ( .A(n30), .B(n310), .C(n311), .D(n312), .Y(r_data_counter[0]) );
  scg10d1_hd U541 ( .A(n313), .B(n314), .C(n315), .D(n29), .Y(
        r_data_counter[1]) );
  ao22d1_hd U542 ( .A(n28), .B(n309), .C(n307), .D(n316), .Y(r_data_counter[2]) );
  nr2d1_hd U544 ( .A(n312), .B(n311), .Y(n315) );
  ivd1_hd U545 ( .A(n30), .Y(n312) );
  ao21d1_hd U546 ( .A(n317), .B(n313), .C(n314), .Y(n309) );
  oa21d1_hd U547 ( .A(n308), .B(n30), .C(n310), .Y(n314) );
  oa211d1_hd U548 ( .A(n308), .B(n318), .C(n319), .D(n320), .Y(n310) );
  ivd1_hd U550 ( .A(n308), .Y(n317) );
  oa211d1_hd U558 ( .A(n332), .B(n333), .C(n265), .D(n334), .Y(n331) );
  scg21d1_hd U559 ( .A(n337), .B(n338), .C(n339), .D(n295), .Y(n336) );
  nr2d1_hd U560 ( .A(n18), .B(n340), .Y(n282) );
  scg14d1_hd U561 ( .A(n27), .B(n344), .C(n345), .Y(n341) );
  ao22d1_hd U562 ( .A(n346), .B(n103), .C(n147), .D(n347), .Y(n345) );
  oa21d1_hd U563 ( .A(n349), .B(n350), .C(n351), .Y(n348) );
  ao22d1_hd U564 ( .A(n346), .B(n102), .C(n95), .D(n347), .Y(n351) );
  oa21d1_hd U565 ( .A(n325), .B(n350), .C(n353), .Y(n352) );
  ao22d1_hd U566 ( .A(n346), .B(n101), .C(n146), .D(n347), .Y(n353) );
  oa21d1_hd U567 ( .A(n326), .B(n350), .C(n355), .Y(n354) );
  ao22d1_hd U568 ( .A(n346), .B(n100), .C(n145), .D(n347), .Y(n355) );
  oa21d1_hd U569 ( .A(n327), .B(n350), .C(n357), .Y(n356) );
  ao22d1_hd U570 ( .A(n346), .B(n99), .C(n94), .D(n347), .Y(n357) );
  ivd1_hd U571 ( .A(n358), .Y(n347) );
  ivd1_hd U572 ( .A(n26), .Y(n327) );
  scg5d1_hd U573 ( .A(n346), .B(n98), .C(n107), .D(n344), .E(n360), .F(n361), 
        .Y(n359) );
  scg5d1_hd U574 ( .A(n346), .B(n97), .C(n106), .D(n344), .E(n363), .F(n360), 
        .Y(n362) );
  scg13d1_hd U578 ( .A(n365), .B(n366), .C(n367), .Y(n342) );
  ivd1_hd U579 ( .A(n368), .Y(n346) );
  scg10d1_hd U580 ( .A(n24), .B(n369), .C(n344), .D(n370), .Y(
        r_spi_data_in_valid) );
  ao211d1_hd U581 ( .A(n372), .B(n373), .C(n365), .D(n374), .Y(n371) );
  nd3d1_hd U582 ( .A(n375), .B(n367), .C(n376), .Y(n369) );
  nr4d1_hd U583 ( .A(n295), .B(n377), .C(n360), .D(n378), .Y(n376) );
  ivd1_hd U584 ( .A(n319), .Y(n295) );
  ao21d1_hd U585 ( .A(n280), .B(n302), .C(n379), .Y(n367) );
  ao22d1_hd U586 ( .A(n267), .B(n380), .C(n381), .D(n265), .Y(n163) );
  nr2d1_hd U587 ( .A(n36), .B(n383), .Y(n380) );
  scg17d1_hd U588 ( .A(n384), .B(n349), .C(n385), .D(n386), .Y(n165) );
  nr4d1_hd U589 ( .A(n387), .B(n388), .C(n384), .D(n267), .Y(n385) );
  ivd1_hd U590 ( .A(n108), .Y(n349) );
  oa22ad1_hd U591 ( .A(n389), .B(n390), .C(n390), .D(o_ADS1292_DATA_VALID), 
        .Y(n162) );
  nr4d1_hd U592 ( .A(n391), .B(n330), .C(n387), .D(n392), .Y(n390) );
  nr2d1_hd U593 ( .A(n393), .B(n394), .Y(n387) );
  nr2d1_hd U594 ( .A(n397), .B(n168), .Y(N985) );
  ao211d1_hd U595 ( .A(n281), .B(n335), .C(n399), .D(n400), .Y(n397) );
  oa211d1_hd U596 ( .A(n401), .B(n350), .C(n402), .D(n320), .Y(n400) );
  nr4d1_hd U597 ( .A(N942), .B(n403), .C(n267), .D(n404), .Y(n402) );
  nr4d1_hd U598 ( .A(n405), .B(n318), .C(n406), .D(n407), .Y(n404) );
  ao21d1_hd U599 ( .A(n13), .B(n149), .C(n408), .Y(n401) );
  oa211d1_hd U600 ( .A(n149), .B(n409), .C(n410), .D(n411), .Y(n408) );
  ao22d1_hd U601 ( .A(n14), .B(n412), .C(n142), .D(n413), .Y(n411) );
  ad2d1_hd U603 ( .A(n415), .B(w_rstn), .Y(N983) );
  nd4d1_hd U604 ( .A(n416), .B(n417), .C(n418), .D(n419), .Y(r_pstate[6]) );
  nr4d1_hd U605 ( .A(n280), .B(n420), .C(n377), .D(n421), .Y(n418) );
  oa21d1_hd U606 ( .A(n318), .B(n422), .C(n423), .Y(n421) );
  ao211d1_hd U607 ( .A(n396), .B(n424), .C(n425), .D(n426), .Y(n417) );
  nd3d1_hd U608 ( .A(n308), .B(n427), .C(n386), .Y(n426) );
  scg13d1_hd U609 ( .A(n383), .B(n265), .C(n36), .Y(n386) );
  scg15d1_hd U610 ( .A(n429), .B(n303), .C(n416), .D(n430), .Y(r_pstate[5]) );
  nr4d1_hd U611 ( .A(n391), .B(n431), .C(n374), .D(n432), .Y(n430) );
  oa211d1_hd U612 ( .A(n428), .B(n433), .C(n434), .D(n422), .Y(n432) );
  oa21d1_hd U613 ( .A(n15), .B(n435), .C(n368), .Y(n374) );
  ivd1_hd U614 ( .A(n375), .Y(n431) );
  ivd1_hd U615 ( .A(n320), .Y(n391) );
  nr4d1_hd U616 ( .A(n278), .B(n436), .C(n384), .D(n437), .Y(n416) );
  scg20d1_hd U617 ( .A(n438), .B(n439), .C(n393), .Y(n437) );
  nr2d1_hd U618 ( .A(n350), .B(n440), .Y(n384) );
  nr2d1_hd U619 ( .A(n318), .B(n406), .Y(n436) );
  nr2bd1_hd U620 ( .AN(n301), .B(n302), .Y(n278) );
  ivd1_hd U621 ( .A(n419), .Y(n303) );
  oa211d1_hd U622 ( .A(n441), .B(n248), .C(n442), .D(n443), .Y(r_pstate[4]) );
  ao211d1_hd U623 ( .A(n444), .B(n318), .C(n378), .D(n445), .Y(n443) );
  oa211d1_hd U624 ( .A(n160), .B(n265), .C(n446), .D(n447), .Y(n445) );
  ao211d1_hd U625 ( .A(n449), .B(n361), .C(n399), .D(n450), .Y(n442) );
  scg18d1_hd U626 ( .A(n18), .B(n451), .C(n452), .D(n453), .E(n322), .Y(n450)
         );
  nd3d1_hd U627 ( .A(n267), .B(n263), .C(n37), .Y(n453) );
  ivd1_hd U628 ( .A(n33), .Y(n263) );
  nr2d1_hd U629 ( .A(n455), .B(n456), .Y(n452) );
  oa21d1_hd U630 ( .A(n429), .B(n419), .C(n329), .Y(n399) );
  nd4d1_hd U631 ( .A(n375), .B(n382), .C(n458), .D(n459), .Y(r_pstate[2]) );
  ao211d1_hd U632 ( .A(n460), .B(n461), .C(n462), .D(n463), .Y(n459) );
  nr4d1_hd U633 ( .A(n464), .B(n339), .C(n279), .D(n465), .Y(n458) );
  oa22d1_hd U634 ( .A(n457), .B(n466), .C(n302), .D(n467), .Y(n279) );
  ivd1_hd U635 ( .A(n300), .Y(n466) );
  nr2d1_hd U636 ( .A(n15), .B(n468), .Y(n300) );
  oa211d1_hd U637 ( .A(n471), .B(n120), .C(n119), .D(n118), .Y(n470) );
  ao211d1_hd U638 ( .A(n472), .B(n473), .C(n474), .D(n475), .Y(n471) );
  nd4d1_hd U639 ( .A(n128), .B(n127), .C(n126), .D(n476), .Y(n472) );
  oa21d1_hd U640 ( .A(n477), .B(n350), .C(n478), .Y(n339) );
  nr2d1_hd U641 ( .A(n35), .B(n467), .Y(n464) );
  ivd1_hd U642 ( .A(n280), .Y(n467) );
  ao22d1_hd U643 ( .A(n429), .B(n396), .C(n301), .D(n302), .Y(n382) );
  nr2d1_hd U644 ( .A(n479), .B(n480), .Y(n375) );
  oa22d1_hd U645 ( .A(n481), .B(n482), .C(n483), .D(n455), .Y(n480) );
  oa211d1_hd U646 ( .A(n337), .B(n338), .C(n484), .D(n485), .Y(r_pstate[1]) );
  ao211d1_hd U647 ( .A(n405), .B(n460), .C(n415), .D(n462), .Y(n485) );
  oa22d1_hd U648 ( .A(n131), .B(n287), .C(w_spi_data_in_ready), .D(n422), .Y(
        n462) );
  nr2bd1_hd U649 ( .AN(w_spi_data_out_valid), .B(n486), .Y(n415) );
  nr2d1_hd U650 ( .A(i_ADS1292_DRDY), .B(n427), .Y(n460) );
  ivd1_hd U651 ( .A(n392), .Y(n427) );
  nr4d1_hd U652 ( .A(n487), .B(n479), .C(n488), .D(n489), .Y(n484) );
  oa211d1_hd U653 ( .A(w_spi_data_in_ready), .B(n308), .C(n434), .D(n291), .Y(
        n489) );
  nr2d1_hd U654 ( .A(n490), .B(n482), .Y(n479) );
  ivd1_hd U655 ( .A(n451), .Y(n482) );
  ivd1_hd U656 ( .A(n491), .Y(n338) );
  or4d1_hd U657 ( .A(n463), .B(n492), .C(n493), .D(n494), .Y(r_pstate[0]) );
  oa22d1_hd U658 ( .A(n35), .B(n441), .C(w_spi_data_out_valid), .D(n486), .Y(
        n494) );
  ao22d1_hd U659 ( .A(i_ADS1292_DRDY), .B(n392), .C(n280), .D(n302), .Y(n441)
         );
  nd2bd1_hd U660 ( .AN(n495), .B(n496), .Y(n302) );
  oa211d1_hd U661 ( .A(n125), .B(n497), .C(n120), .D(n121), .Y(n496) );
  nr2d1_hd U662 ( .A(n498), .B(n499), .Y(n280) );
  nr2d1_hd U663 ( .A(n490), .B(n500), .Y(n392) );
  oa211d1_hd U664 ( .A(n276), .B(n501), .C(n274), .D(n502), .Y(n493) );
  ao22d1_hd U665 ( .A(n425), .B(i_ADS1292_DRDY), .C(n503), .D(n272), .Y(n502)
         );
  oa21d1_hd U666 ( .A(n132), .B(n133), .C(n506), .Y(n505) );
  oa21d1_hd U667 ( .A(n507), .B(n508), .C(n509), .Y(n506) );
  ao211d1_hd U668 ( .A(n510), .B(n511), .C(n112), .D(n111), .Y(n507) );
  scg22d1_hd U669 ( .A(n117), .B(n512), .C(n513), .D(n514), .Y(n510) );
  ao21d1_hd U670 ( .A(n119), .B(n120), .C(n118), .Y(n513) );
  oa211d1_hd U671 ( .A(n515), .B(n475), .C(n474), .D(n516), .Y(n512) );
  ivd1_hd U672 ( .A(n121), .Y(n474) );
  nr4d1_hd U673 ( .A(n125), .B(n126), .C(n123), .D(n517), .Y(n515) );
  ivd1_hd U674 ( .A(n273), .Y(n503) );
  ivd1_hd U675 ( .A(n285), .Y(n487) );
  nr2d1_hd U676 ( .A(n395), .B(n333), .Y(n425) );
  ivd1_hd U677 ( .A(n500), .Y(n454) );
  ivd1_hd U678 ( .A(n332), .Y(n395) );
  ao21d1_hd U679 ( .A(n491), .B(n337), .C(n420), .Y(n274) );
  nr2d1_hd U680 ( .A(n335), .B(n520), .Y(n420) );
  oa21d1_hd U681 ( .A(n521), .B(n522), .C(n523), .Y(n335) );
  ao211d1_hd U682 ( .A(n476), .B(n524), .C(n123), .D(n525), .Y(n521) );
  scg6d1_hd U683 ( .A(n128), .B(n127), .C(n126), .Y(n524) );
  ad2d1_hd U684 ( .A(n125), .B(n124), .Y(n476) );
  nr4d1_hd U685 ( .A(n121), .B(n120), .C(n497), .D(n495), .Y(n337) );
  nd3bd1_hd U686 ( .AN(n119), .B(n469), .C(n516), .Y(n495) );
  ivd1_hd U687 ( .A(n118), .Y(n516) );
  nr2bd1_hd U688 ( .AN(n523), .B(n117), .Y(n469) );
  scg12d1_hd U689 ( .A(n526), .B(n514), .C(n114), .Y(n523) );
  nr3d1_hd U690 ( .A(n113), .B(n116), .C(n115), .Y(n514) );
  nr4d1_hd U691 ( .A(n110), .B(n109), .C(n527), .D(n528), .Y(n526) );
  scg13d1_hd U692 ( .A(n124), .B(n123), .C(n475), .Y(n497) );
  nr2d1_hd U693 ( .A(n490), .B(n340), .Y(n491) );
  ivd1_hd U694 ( .A(n277), .Y(n501) );
  nr2d1_hd U695 ( .A(n15), .B(n423), .Y(n277) );
  scg20d1_hd U696 ( .A(n529), .B(n508), .C(n528), .Y(n276) );
  nd3bd1_hd U697 ( .AN(n132), .B(n509), .C(n504), .Y(n528) );
  nr2d1_hd U698 ( .A(n530), .B(n531), .Y(n504) );
  or4d1_hd U699 ( .A(n140), .B(n137), .C(n138), .D(n134), .Y(n531) );
  or4d1_hd U700 ( .A(n136), .B(n135), .C(n141), .D(n139), .Y(n530) );
  nr3d1_hd U701 ( .A(n133), .B(n129), .C(n130), .Y(n509) );
  scg21d1_hd U702 ( .A(n522), .B(n532), .C(n511), .D(n527), .Y(n529) );
  or2d1_hd U703 ( .A(n112), .B(n111), .Y(n527) );
  or2d1_hd U704 ( .A(n114), .B(n113), .Y(n511) );
  oa211d1_hd U705 ( .A(n533), .B(n525), .C(n116), .D(n115), .Y(n532) );
  scg13d1_hd U706 ( .A(n121), .B(n120), .C(n475), .Y(n525) );
  scg11d1_hd U708 ( .A(n126), .B(n517), .C(n125), .D(n124), .E(n473), .Y(n533)
         );
  or3d1_hd U710 ( .A(n128), .B(n127), .C(n124), .Y(n517) );
  nd3d1_hd U711 ( .A(n118), .B(n119), .C(n117), .Y(n522) );
  oa211d1_hd U712 ( .A(n438), .B(n393), .C(n534), .D(n535), .Y(n492) );
  nr4d1_hd U713 ( .A(n301), .B(n294), .C(n379), .D(n366), .Y(n535) );
  nr2d1_hd U714 ( .A(n16), .B(n435), .Y(n360) );
  ivd1_hd U715 ( .A(n449), .Y(n435) );
  oa21d1_hd U716 ( .A(n318), .B(n537), .C(n446), .Y(n379) );
  nd3d1_hd U717 ( .A(n344), .B(n477), .C(n440), .Y(n446) );
  nd3d1_hd U718 ( .A(n143), .B(n538), .C(n325), .Y(n440) );
  ivd1_hd U719 ( .A(n144), .Y(n325) );
  nd4d1_hd U720 ( .A(n144), .B(n108), .C(n538), .D(n326), .Y(n477) );
  nr2d1_hd U722 ( .A(n26), .B(n539), .Y(n538) );
  or4d1_hd U723 ( .A(n107), .B(n106), .C(n27), .D(n105), .Y(n539) );
  ivd1_hd U724 ( .A(n350), .Y(n344) );
  nr2d1_hd U725 ( .A(n488), .B(n465), .Y(n537) );
  nd3d1_hd U726 ( .A(n373), .B(n16), .C(n372), .Y(n308) );
  ivd1_hd U727 ( .A(n499), .Y(n372) );
  nr2d1_hd U728 ( .A(n15), .B(n455), .Y(n488) );
  nr2d1_hd U729 ( .A(n17), .B(n540), .Y(n449) );
  ivd1_hd U730 ( .A(w_spi_data_in_ready), .Y(n318) );
  nr2d1_hd U731 ( .A(n541), .B(n542), .Y(n301) );
  nr2d1_hd U732 ( .A(n365), .B(n378), .Y(n534) );
  nr2d1_hd U733 ( .A(w_spi_data_in_ready), .B(n406), .Y(n378) );
  ad3d1_hd U734 ( .A(n451), .B(n361), .C(w_spi_data_in_ready), .Y(n365) );
  nr2d1_hd U735 ( .A(n15), .B(n481), .Y(n361) );
  nr3d1_hd U736 ( .A(n540), .B(n543), .C(n16), .Y(n451) );
  ivd1_hd U737 ( .A(n396), .Y(n393) );
  nr2d1_hd U738 ( .A(n499), .B(n542), .Y(n396) );
  nr3d1_hd U739 ( .A(n429), .B(n439), .C(n424), .Y(n438) );
  nd3d1_hd U740 ( .A(n13), .B(n545), .C(n413), .Y(n414) );
  ivd1_hd U741 ( .A(n405), .Y(n461) );
  nr4d1_hd U742 ( .A(n14), .B(n13), .C(n142), .D(n546), .Y(n405) );
  oa211d1_hd U743 ( .A(n547), .B(n412), .C(n548), .D(n549), .Y(n439) );
  nd4d1_hd U744 ( .A(n150), .B(n12), .C(n409), .D(n550), .Y(n549) );
  ad2d1_hd U745 ( .A(n13), .B(n412), .Y(n409) );
  ivd1_hd U746 ( .A(n407), .Y(n548) );
  nd4d1_hd U747 ( .A(n13), .B(n551), .C(n413), .D(n412), .Y(n332) );
  nr2d1_hd U748 ( .A(n412), .B(n546), .Y(n545) );
  ivd1_hd U749 ( .A(n142), .Y(n412) );
  nr2d1_hd U750 ( .A(n142), .B(n547), .Y(n429) );
  ad2d1_hd U751 ( .A(n410), .B(n550), .Y(n551) );
  ivd1_hd U752 ( .A(n149), .Y(n550) );
  nr2d1_hd U753 ( .A(n150), .B(n12), .Y(n410) );
  nr2d1_hd U754 ( .A(n13), .B(n413), .Y(n552) );
  ivd1_hd U755 ( .A(n14), .Y(n413) );
  oa22d1_hd U756 ( .A(w_spi_data_out_valid), .B(n389), .C(n34), .D(n298), .Y(
        n463) );
  scg13d1_hd U757 ( .A(n36), .B(n433), .C(n428), .Y(n298) );
  nr2d1_hd U758 ( .A(n37), .B(n33), .Y(n428) );
  ivd1_hd U760 ( .A(n377), .Y(n389) );
  ivd1_hd U761 ( .A(n330), .Y(n329) );
  nr2d1_hd U762 ( .A(n499), .B(n554), .Y(n330) );
  nr2d1_hd U763 ( .A(n18), .B(n15), .Y(n363) );
  scg17d1_hd U764 ( .A(n536), .B(n18), .C(n444), .D(n520), .Y(r_lstate[4]) );
  ivd1_hd U765 ( .A(n281), .Y(n520) );
  nr2d1_hd U766 ( .A(n481), .B(n422), .Y(n444) );
  oa211d1_hd U767 ( .A(n498), .B(n490), .C(n468), .D(n422), .Y(r_lstate[2]) );
  ivd1_hd U768 ( .A(n555), .Y(n490) );
  ivd1_hd U769 ( .A(N942), .Y(n422) );
  nr4d1_hd U770 ( .A(n15), .B(n557), .C(n543), .D(n540), .Y(N942) );
  nd3bd1_hd U771 ( .AN(n304), .B(n553), .C(n406), .Y(r_lstate[0]) );
  ivd1_hd U772 ( .A(n340), .Y(n536) );
  nr3d1_hd U773 ( .A(n281), .B(n377), .C(n294), .Y(n553) );
  nr2d1_hd U774 ( .A(n483), .B(n423), .Y(n294) );
  nr2d1_hd U775 ( .A(n498), .B(n541), .Y(n377) );
  nr2d1_hd U776 ( .A(n18), .B(n483), .Y(n555) );
  nr2d1_hd U777 ( .A(n500), .B(n456), .Y(n281) );
  ivd1_hd U778 ( .A(n448), .Y(n456) );
  nr2d1_hd U779 ( .A(n481), .B(n483), .Y(n448) );
  ivd1_hd U780 ( .A(n554), .Y(n558) );
  nd2bd1_hd U781 ( .AN(n19), .B(n544), .Y(n554) );
  nr2d1_hd U782 ( .A(n17), .B(n16), .Y(n544) );
  ivd1_hd U783 ( .A(n556), .Y(n403) );
  nr4d1_hd U784 ( .A(n19), .B(n17), .C(n18), .D(n557), .Y(n519) );
  nd3bd1_hd U786 ( .AN(n498), .B(n518), .C(n481), .Y(n468) );
  nr2d1_hd U790 ( .A(n19), .B(n543), .Y(n373) );
  fd3qd1_hd clk_r_REG15_S5 ( .D(n164), .CK(n572), .SN(n167), .Q(
        o_ADS1292_RESET) );
  fd3qd1_hd clk_r_REG21_S6 ( .D(n166), .CK(n572), .SN(n167), .Q(o_SPI_CSN) );
  ivd1_hd clk_r_REG98_S6_U5 ( .A(n289), .Y(n171) );
  mx2id1_hd u_cell_7677 ( .D0(n171), .D1(n288), .S(n32), .YN(n170) );
  fd4qd1_hd clk_r_REG98_S6 ( .D(n170), .CK(i_CLK), .SN(1'b1), .RN(n167), .Q(
        n32) );
  fd1eqd1_hd clk_r_REG99_S8 ( .D(r_lstate[2]), .E(N985), .CK(n572), .Q(n13) );
  fd1eqd1_hd clk_r_REG96_S3 ( .D(r_lstate[0]), .E(N985), .CK(n572), .Q(n142)
         );
  fd1eqd1_hd clk_r_REG92_S3 ( .D(N1171), .E(N985), .CK(n572), .Q(n149) );
  fd2d1_hd clk_r_REG103_S8 ( .D(n597), .CK(n570), .RN(n167), .Q(n143), .QN(
        n326) );
  fd2d1_hd clk_r_REG128_S3 ( .D(r_clk_counter[5]), .CK(n572), .RN(n167), .Q(
        n123), .QN(n473) );
  fd2d1_hd clk_r_REG90_S13 ( .D(r_data_counter[1]), .CK(n572), .RN(n167), .Q(
        n29), .QN(n313) );
  fd2d1_hd clk_r_REG89_S13 ( .D(r_data_counter[2]), .CK(n572), .RN(n167), .Q(
        n28), .QN(n316) );
  fd2d1_hd clk_r_REG17_S6 ( .D(r_pstate[4]), .CK(i_CLK), .RN(n167), .Q(n18), 
        .QN(n481) );
  fd2d1_hd clk_r_REG16_S5 ( .D(r_pstate[2]), .CK(i_CLK), .RN(n167), .Q(n17), 
        .QN(n543) );
  fd2d1_hd clk_r_REG23_S7 ( .D(r_pstate[1]), .CK(i_CLK), .RN(n167), .Q(n16), 
        .QN(n557) );
  fd2d1_hd clk_r_REG22_S6 ( .D(r_pstate[0]), .CK(i_CLK), .RN(n167), .Q(n15), 
        .QN(n483) );
  nid4_hd U1 ( .A(w_rstn), .Y(n167) );
  ivd1_hd U2 ( .A(w_rstn), .Y(n168) );
  ivd1_hd U3 ( .A(n122), .Y(n475) );
  fd1qd1_hd clk_r_REG33_S14 ( .D(n86), .CK(n565), .Q(o_ADS1292_DATA_OUT[0]) );
  fd1qd1_hd clk_r_REG35_S15 ( .D(n70), .CK(n565), .Q(o_ADS1292_DATA_OUT[8]) );
  fd1qd1_hd clk_r_REG37_S16 ( .D(n54), .CK(n565), .Q(o_ADS1292_DATA_OUT[16])
         );
  fd1qd1_hd clk_r_REG40_S14 ( .D(n84), .CK(n565), .Q(o_ADS1292_DATA_OUT[1]) );
  fd1qd1_hd clk_r_REG42_S15 ( .D(n68), .CK(n565), .Q(o_ADS1292_DATA_OUT[9]) );
  fd1qd1_hd clk_r_REG44_S16 ( .D(n52), .CK(n565), .Q(o_ADS1292_DATA_OUT[17])
         );
  fd1qd1_hd clk_r_REG47_S14 ( .D(n82), .CK(n565), .Q(o_ADS1292_DATA_OUT[2]) );
  fd1qd1_hd clk_r_REG49_S15 ( .D(n66), .CK(n565), .Q(o_ADS1292_DATA_OUT[10])
         );
  fd1qd1_hd clk_r_REG51_S16 ( .D(n50), .CK(n565), .Q(o_ADS1292_DATA_OUT[18])
         );
  fd1qd1_hd clk_r_REG54_S14 ( .D(n80), .CK(n565), .Q(o_ADS1292_DATA_OUT[3]) );
  fd1qd1_hd clk_r_REG56_S15 ( .D(n64), .CK(n565), .Q(o_ADS1292_DATA_OUT[11])
         );
  fd1qd1_hd clk_r_REG58_S16 ( .D(n48), .CK(n565), .Q(o_ADS1292_DATA_OUT[19])
         );
  fd1qd1_hd clk_r_REG61_S14 ( .D(n78), .CK(n565), .Q(o_ADS1292_DATA_OUT[4]) );
  fd1qd1_hd clk_r_REG63_S15 ( .D(n62), .CK(n565), .Q(o_ADS1292_DATA_OUT[12])
         );
  fd1qd1_hd clk_r_REG65_S16 ( .D(n39), .CK(n565), .Q(o_ADS1292_DATA_OUT[20])
         );
  fd1qd1_hd clk_r_REG68_S14 ( .D(n76), .CK(n565), .Q(o_ADS1292_DATA_OUT[5]) );
  fd1qd1_hd clk_r_REG70_S15 ( .D(n60), .CK(n565), .Q(o_ADS1292_DATA_OUT[13])
         );
  fd1qd1_hd clk_r_REG72_S16 ( .D(n41), .CK(n565), .Q(o_ADS1292_DATA_OUT[21])
         );
  fd1qd1_hd clk_r_REG75_S14 ( .D(n74), .CK(n565), .Q(o_ADS1292_DATA_OUT[6]) );
  fd1qd1_hd clk_r_REG77_S15 ( .D(n58), .CK(n565), .Q(o_ADS1292_DATA_OUT[14])
         );
  fd1qd1_hd clk_r_REG79_S16 ( .D(n43), .CK(n565), .Q(o_ADS1292_DATA_OUT[22])
         );
  fd1qd1_hd clk_r_REG82_S14 ( .D(n72), .CK(n565), .Q(o_ADS1292_DATA_OUT[7]) );
  fd1qd1_hd clk_r_REG84_S15 ( .D(n56), .CK(n565), .Q(o_ADS1292_DATA_OUT[15])
         );
  fd1qd1_hd clk_r_REG86_S16 ( .D(n45), .CK(n565), .Q(o_ADS1292_DATA_OUT[23])
         );
  fd1qd1_hd clk_r_REG31_S13 ( .D(w_spi_data_out[0]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[0]) );
  fd1qd1_hd clk_r_REG38_S13 ( .D(w_spi_data_out[1]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[1]) );
  fd1qd1_hd clk_r_REG45_S13 ( .D(w_spi_data_out[2]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[2]) );
  fd1qd1_hd clk_r_REG52_S13 ( .D(w_spi_data_out[3]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[3]) );
  fd1qd1_hd clk_r_REG59_S13 ( .D(w_spi_data_out[4]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[4]) );
  fd1qd1_hd clk_r_REG66_S13 ( .D(w_spi_data_out[5]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[5]) );
  fd1qd1_hd clk_r_REG73_S13 ( .D(w_spi_data_out[6]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[6]) );
  fd1qd1_hd clk_r_REG80_S13 ( .D(w_spi_data_out[7]), .CK(n568), .Q(
        o_ADS1292_REG_DATA_OUT[7]) );
  fd1qd1_hd clk_r_REG95_S7 ( .D(r_lstate[4]), .CK(n571), .Q(n14) );
  fd1qd1_hd clk_r_REG118_S7 ( .D(N942), .CK(n571), .Q(n12) );
  fd1qd1_hd clk_r_REG119_S7 ( .D(r_lstate[1]), .CK(n571), .Q(n150) );
  fd3qd1_hd clk_r_REG146_S1 ( .D(n574), .CK(i_CLK), .SN(n167), .Q(n160) );
  ads1292_controller_DW01_inc_0 add_x_2 ( .A({n141, n140, n139, n138, n137, 
        n136, n135, n134, n133, n132, n130, n129, n109, n110, n111, n112, n113, 
        n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
        n126, n127, n128}), .SUM({N362, N361, N360, N359, N358, N357, N356, 
        N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, 
        N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, 
        N331}) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_14 clk_gate_clk_r_REG9_S3_0 ( .CLK(
        i_CLK), .EN(n588), .ENCLK(n572), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_15 clk_gate_clk_r_REG95_S7_0 ( .CLK(
        i_CLK), .EN(N985), .ENCLK(n571), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_16 clk_gate_clk_r_REG103_S8_0 ( 
        .CLK(i_CLK), .EN(n599), .ENCLK(n570), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_17 clk_gate_clk_r_REG14_S5_0 ( .CLK(
        i_CLK), .EN(n342), .ENCLK(n569), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_18 clk_gate_clk_r_REG31_S13_0 ( 
        .CLK(i_CLK), .EN(N983), .ENCLK(n568), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_19 clk_gate_clk_r_REG114_S8_0 ( 
        .CLK(i_CLK), .EN(n267), .ENCLK(n567), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_20 clk_gate_clk_r_REG32_S13_0 ( 
        .CLK(i_CLK), .EN(n286), .ENCLK(n566), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ads1292_controller_21 clk_gate_clk_r_REG33_S14_0 ( 
        .CLK(i_CLK), .EN(N984), .ENCLK(n565), .TE(1'b0) );
  fd4qd1_hd clk_r_REG3_S2 ( .D(r_pstate[6]), .CK(i_CLK), .SN(1'b1), .RN(n167), 
        .Q(n20) );
  fd4qd1_hd clk_r_REG85_S15 ( .D(n56), .CK(n566), .SN(1'b1), .RN(n167), .Q(n45) );
  fd4qd1_hd clk_r_REG83_S14 ( .D(n72), .CK(n566), .SN(1'b1), .RN(n167), .Q(n56) );
  fd4qd1_hd clk_r_REG81_S13 ( .D(w_spi_data_out[7]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n72) );
  fd4qd1_hd clk_r_REG78_S15 ( .D(n58), .CK(n566), .SN(1'b1), .RN(n167), .Q(n43) );
  fd4qd1_hd clk_r_REG76_S14 ( .D(n74), .CK(n566), .SN(1'b1), .RN(n167), .Q(n58) );
  fd4qd1_hd clk_r_REG74_S13 ( .D(w_spi_data_out[6]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n74) );
  fd4qd1_hd clk_r_REG71_S15 ( .D(n60), .CK(n566), .SN(1'b1), .RN(n167), .Q(n41) );
  fd4qd1_hd clk_r_REG69_S14 ( .D(n76), .CK(n566), .SN(1'b1), .RN(n167), .Q(n60) );
  fd4qd1_hd clk_r_REG67_S13 ( .D(w_spi_data_out[5]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n76) );
  fd4qd1_hd clk_r_REG64_S15 ( .D(n62), .CK(n566), .SN(1'b1), .RN(n167), .Q(n39) );
  fd4qd1_hd clk_r_REG62_S14 ( .D(n78), .CK(n566), .SN(1'b1), .RN(n167), .Q(n62) );
  fd4qd1_hd clk_r_REG60_S13 ( .D(w_spi_data_out[4]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n78) );
  fd4qd1_hd clk_r_REG57_S15 ( .D(n64), .CK(n566), .SN(1'b1), .RN(n167), .Q(n48) );
  fd4qd1_hd clk_r_REG55_S14 ( .D(n80), .CK(n566), .SN(1'b1), .RN(n167), .Q(n64) );
  fd4qd1_hd clk_r_REG53_S13 ( .D(w_spi_data_out[3]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n80) );
  fd4qd1_hd clk_r_REG50_S15 ( .D(n66), .CK(n566), .SN(1'b1), .RN(n167), .Q(n50) );
  fd4qd1_hd clk_r_REG48_S14 ( .D(n82), .CK(n566), .SN(1'b1), .RN(n167), .Q(n66) );
  fd4qd1_hd clk_r_REG46_S13 ( .D(w_spi_data_out[2]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n82) );
  fd4qd1_hd clk_r_REG43_S15 ( .D(n68), .CK(n566), .SN(1'b1), .RN(n167), .Q(n52) );
  fd4qd1_hd clk_r_REG41_S14 ( .D(n84), .CK(n566), .SN(1'b1), .RN(n167), .Q(n68) );
  fd4qd1_hd clk_r_REG39_S13 ( .D(w_spi_data_out[1]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n84) );
  fd4qd1_hd clk_r_REG36_S15 ( .D(n70), .CK(n566), .SN(1'b1), .RN(n167), .Q(n54) );
  fd4qd1_hd clk_r_REG34_S14 ( .D(n86), .CK(n566), .SN(1'b1), .RN(n167), .Q(n70) );
  fd4qd1_hd clk_r_REG32_S13 ( .D(w_spi_data_out[0]), .CK(n566), .SN(1'b1), 
        .RN(n167), .Q(n86) );
  fd4qd1_hd clk_r_REG93_S4 ( .D(n161), .CK(n572), .SN(1'b1), .RN(n167), .Q(
        o_ADS1292_INIT_SET) );
  fd4qd1_hd clk_r_REG29_S8 ( .D(n600), .CK(n569), .SN(1'b1), .RN(n167), .Q(n25) );
  fd4qd1_hd clk_r_REG26_S8 ( .D(n356), .CK(n569), .SN(1'b1), .RN(n167), .Q(n89) );
  fd4qd1_hd clk_r_REG25_S8 ( .D(n354), .CK(n569), .SN(1'b1), .RN(n167), .Q(n90) );
  fd4qd1_hd clk_r_REG24_S8 ( .D(n352), .CK(n569), .SN(1'b1), .RN(n167), .Q(n91) );
  fd4qd1_hd clk_r_REG14_S5 ( .D(n348), .CK(n569), .SN(1'b1), .RN(n167), .Q(n92) );
  fd4qd1_hd clk_r_REG19_S5 ( .D(n341), .CK(n569), .SN(1'b1), .RN(n167), .Q(n93) );
  fd4qd1_hd clk_r_REG28_S8 ( .D(n362), .CK(n569), .SN(1'b1), .RN(n167), .Q(n87) );
  fd4qd1_hd clk_r_REG27_S8 ( .D(n359), .CK(n569), .SN(1'b1), .RN(n167), .Q(n88) );
  fd4qd1_hd clk_r_REG91_S13 ( .D(n162), .CK(n572), .SN(1'b1), .RN(n167), .Q(
        o_ADS1292_DATA_VALID) );
  fd4qd1_hd clk_r_REG2_S2 ( .D(n165), .CK(n572), .SN(1'b1), .RN(n167), .Q(
        o_ADS1292_START) );
  fd4qd1_hd clk_r_REG87_S13 ( .D(r_data_counter[0]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n30) );
  fd4qd1_hd clk_r_REG20_S5 ( .D(r_pstate[5]), .CK(i_CLK), .SN(1'b1), .RN(n167), 
        .Q(n19) );
  fd4qd1_hd clk_r_REG1_S2 ( .D(n163), .CK(n572), .SN(1'b1), .RN(n167), .Q(
        o_ADS1292_BUSY) );
  fd4qd1_hd clk_r_REG148_S1 ( .D(i_ADS1292_DRDY), .CK(i_CLK), .SN(1'b1), .RN(
        n167), .Q(n159) );
  fd4qd1_hd clk_r_REG111_S8 ( .D(i_ADS1292_DATA_IN[7]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n96) );
  fd4qd1_hd clk_r_REG110_S8 ( .D(i_ADS1292_DATA_IN[6]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n97) );
  fd4qd1_hd clk_r_REG109_S8 ( .D(i_ADS1292_DATA_IN[5]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n98) );
  fd4qd1_hd clk_r_REG108_S8 ( .D(i_ADS1292_DATA_IN[4]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n99) );
  fd4qd1_hd clk_r_REG107_S8 ( .D(i_ADS1292_DATA_IN[3]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n100) );
  fd4qd1_hd clk_r_REG106_S8 ( .D(i_ADS1292_DATA_IN[2]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n101) );
  fd4qd1_hd clk_r_REG105_S8 ( .D(i_ADS1292_DATA_IN[1]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n102) );
  fd4qd1_hd clk_r_REG104_S8 ( .D(i_ADS1292_DATA_IN[0]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n103) );
  fd4qd1_hd clk_r_REG112_S8 ( .D(i_ADS1292_REG_ADDR[1]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n95) );
  fd4qd1_hd clk_r_REG100_S8 ( .D(i_ADS1292_REG_ADDR[2]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n146) );
  fd4qd1_hd clk_r_REG114_S8 ( .D(i_ADS1292_REG_ADDR[0]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n147) );
  fd4qd1_hd clk_r_REG113_S8 ( .D(i_ADS1292_REG_ADDR[4]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n94) );
  fd4qd1_hd clk_r_REG102_S8 ( .D(i_ADS1292_REG_ADDR[3]), .CK(n567), .SN(1'b1), 
        .RN(n167), .Q(n145) );
  fd4qd1_hd clk_r_REG88_S13 ( .D(r_data_counter[3]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n131) );
  fd4qd1_hd clk_r_REG135_S3 ( .D(r_clk_counter[12]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n116) );
  fd4qd1_hd clk_r_REG134_S3 ( .D(r_clk_counter[11]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n117) );
  fd4qd1_hd clk_r_REG133_S3 ( .D(r_clk_counter[10]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n118) );
  fd4qd1_hd clk_r_REG132_S3 ( .D(r_clk_counter[9]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n119) );
  fd4qd1_hd clk_r_REG131_S3 ( .D(r_clk_counter[8]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n120) );
  fd4qd1_hd clk_r_REG130_S3 ( .D(r_clk_counter[7]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n121) );
  fd4qd1_hd clk_r_REG129_S3 ( .D(r_clk_counter[6]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n122) );
  fd4qd1_hd clk_r_REG127_S3 ( .D(r_clk_counter[4]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n124) );
  fd4qd1_hd clk_r_REG126_S3 ( .D(r_clk_counter[3]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n125) );
  fd4qd1_hd clk_r_REG125_S3 ( .D(r_clk_counter[2]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n126) );
  fd4qd1_hd clk_r_REG124_S3 ( .D(r_clk_counter[1]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n127) );
  fd4qd1_hd clk_r_REG123_S3 ( .D(r_clk_counter[0]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n128) );
  fd4qd1_hd clk_r_REG136_S3 ( .D(r_clk_counter[13]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n115) );
  fd4qd1_hd clk_r_REG116_S4 ( .D(n590), .CK(n570), .SN(1'b1), .RN(n167), .Q(
        n106) );
  fd4qd1_hd clk_r_REG117_S4 ( .D(n591), .CK(n570), .SN(1'b1), .RN(n167), .Q(
        n105) );
  fd4qd1_hd clk_r_REG115_S4 ( .D(n592), .CK(n570), .SN(1'b1), .RN(n167), .Q(
        n107) );
  fd4qd1_hd clk_r_REG30_S8 ( .D(r_spi_data_in_valid), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n24) );
  fd4qd1_hd clk_r_REG101_S8 ( .D(n563), .CK(n570), .SN(1'b1), .RN(n167), .Q(
        n144) );
  fd4qd1_hd clk_r_REG13_S4 ( .D(n593), .CK(n570), .SN(1'b1), .RN(n167), .Q(
        n108) );
  fd4qd1_hd clk_r_REG94_S4 ( .D(n595), .CK(n570), .SN(1'b1), .RN(n167), .Q(n26) );
  fd4qd1_hd clk_r_REG137_S3 ( .D(r_clk_counter[14]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n114) );
  fd4qd1_hd clk_r_REG18_S4 ( .D(n594), .CK(n570), .SN(1'b1), .RN(n167), .Q(n27) );
  fd4qd1_hd clk_r_REG138_S3 ( .D(r_clk_counter[15]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n113) );
  fd4qd1_hd clk_r_REG97_S6 ( .D(r_drdy_edge_counter_1_), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n104) );
  fd4qd1_hd clk_r_REG139_S3 ( .D(r_clk_counter[16]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n112) );
  fd4qd1_hd clk_r_REG140_S3 ( .D(r_clk_counter[17]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n111) );
  fd4qd1_hd clk_r_REG141_S3 ( .D(r_clk_counter[18]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n110) );
  fd4qd1_hd clk_r_REG142_S3 ( .D(r_clk_counter[19]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n109) );
  fd4qd1_hd clk_r_REG147_S1 ( .D(n573), .CK(i_CLK), .SN(1'b1), .RN(n167), .Q(
        n33) );
  fd4qd1_hd clk_r_REG144_S1 ( .D(n576), .CK(i_CLK), .SN(1'b1), .RN(n167), .Q(
        n37) );
  fd4qd1_hd clk_r_REG143_S1 ( .D(n577), .CK(i_CLK), .SN(1'b1), .RN(n167), .Q(
        n35) );
  fd4qd1_hd clk_r_REG0_S1 ( .D(n578), .CK(i_CLK), .SN(1'b1), .RN(n167), .Q(n36) );
  fd4qd1_hd clk_r_REG122_S3 ( .D(r_clk_counter[20]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n129) );
  fd4qd1_hd clk_r_REG121_S3 ( .D(r_clk_counter[21]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n130) );
  fd4qd1_hd clk_r_REG120_S3 ( .D(r_clk_counter[22]), .CK(n572), .SN(1'b1), 
        .RN(n167), .Q(n132) );
  fd4qd1_hd clk_r_REG12_S3 ( .D(r_clk_counter[23]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n133) );
  fd4qd1_hd clk_r_REG145_S1 ( .D(n575), .CK(i_CLK), .SN(1'b1), .RN(n167), .Q(
        n34) );
  fd4qd1_hd clk_r_REG11_S3 ( .D(r_clk_counter[24]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n134) );
  fd4qd1_hd clk_r_REG10_S3 ( .D(r_clk_counter[25]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n135) );
  fd4qd1_hd clk_r_REG9_S3 ( .D(r_clk_counter[26]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n136) );
  fd4qd1_hd clk_r_REG8_S3 ( .D(r_clk_counter[27]), .CK(n572), .SN(1'b1), .RN(
        n167), .Q(n137) );
  fd4qd1_hd clk_r_REG7_S3 ( .D(r_clk_counter[28]), .CK(n572), .SN(1'b1), .RN(
        w_rstn), .Q(n138) );
  fd4qd1_hd clk_r_REG6_S3 ( .D(r_clk_counter[29]), .CK(n572), .SN(1'b1), .RN(
        w_rstn), .Q(n139) );
  fd4qd1_hd clk_r_REG5_S3 ( .D(r_clk_counter[30]), .CK(n572), .SN(1'b1), .RN(
        w_rstn), .Q(n140) );
  fd4qd1_hd clk_r_REG4_S3 ( .D(r_clk_counter[31]), .CK(n572), .SN(1'b1), .RN(
        w_rstn), .Q(n141) );
  clknd2d1_hd U5 ( .A(n377), .B(w_spi_data_out_valid), .Y(n287) );
  nr3d1_hd U6 ( .A(n393), .B(n168), .C(n414), .Y(N984) );
  ivd1_hd U7 ( .A(n287), .Y(n286) );
  nr2ad1_hd U8 ( .A(n468), .B(n483), .Y(n267) );
  mx2d1_hd U9 ( .D0(n34), .D1(n261), .S(n584), .Y(n575) );
  mx2d1_hd U10 ( .D0(n36), .D1(n262), .S(n581), .Y(n578) );
  mx2d1_hd U11 ( .D0(n35), .D1(n262), .S(n582), .Y(n577) );
  mx2d1_hd U12 ( .D0(n37), .D1(n261), .S(n583), .Y(n576) );
  mx2d1_hd U13 ( .D0(n33), .D1(n261), .S(n586), .Y(n573) );
  scg2d1_hd U14 ( .A(n105), .B(n344), .C(n96), .D(n346), .Y(n600) );
  mx2d1_hd U15 ( .D0(n160), .D1(i_ADS1292_CONTROL[2]), .S(n585), .Y(n574) );
  clknd2d1_hd U16 ( .A(n262), .B(i_ADS1292_CONTROL[0]), .Y(n580) );
  ivd1_hd U17 ( .A(n269), .Y(n597) );
  ivd1_hd U116 ( .A(n20), .Y(n518) );
  ad2d1_hd U118 ( .A(n267), .B(i_ADS1292_REG_ADDR[2]), .Y(n563) );
  or2d1_hd U119 ( .A(n330), .B(n331), .Y(n564) );
  scg9d1_hd U120 ( .A(n253), .B(i_ADS1292_CONTROL[1]), .C(i_ADS1292_CONTROL[2]), .Y(n581) );
  scg9d1_hd U121 ( .A(i_ADS1292_CONTROL[0]), .B(i_ADS1292_CONTROL[1]), .C(
        i_ADS1292_CONTROL[2]), .Y(n582) );
  scg9d1_hd U122 ( .A(i_ADS1292_CONTROL[0]), .B(i_ADS1292_CONTROL[2]), .C(
        i_ADS1292_CONTROL[1]), .Y(n583) );
  scg16d1_hd U123 ( .A(i_ADS1292_CONTROL[2]), .B(n262), .C(n579), .Y(n584) );
  nd3d1_hd U124 ( .A(n262), .B(n261), .C(n253), .Y(n579) );
  ao22d1_hd U125 ( .A(n261), .B(n580), .C(n262), .D(i_ADS1292_CONTROL[2]), .Y(
        n585) );
  scg9d1_hd U126 ( .A(n253), .B(i_ADS1292_CONTROL[2]), .C(i_ADS1292_CONTROL[1]), .Y(n586) );
  nd4d1_hd U127 ( .A(n17), .B(n15), .C(n16), .D(n19), .Y(n588) );
  ad2d1_hd U128 ( .A(n267), .B(i_ADS1292_REG_ADDR[6]), .Y(n590) );
  ad2d1_hd U129 ( .A(n267), .B(i_ADS1292_REG_ADDR[7]), .Y(n591) );
  ad2d1_hd U130 ( .A(n267), .B(i_ADS1292_REG_ADDR[5]), .Y(n592) );
  ad2d1_hd U131 ( .A(n267), .B(i_ADS1292_REG_ADDR[1]), .Y(n593) );
  nd2bd1_hd U132 ( .AN(n596), .B(n266), .Y(n594) );
  or3d1_hd U133 ( .A(n330), .B(i_ADS1292_REG_ADDR[4]), .C(n596), .Y(n595) );
  ivd1_hd U134 ( .A(n322), .Y(n596) );
  nd2bd1_hd U135 ( .AN(n564), .B(n269), .Y(n599) );
endmodule


module khu_sensor_top ( i_CLK, i_RSTN, UART_RXD, UART_TXD, MPR121_SCL_IN, 
        MPR121_SDA_IN, MPR121_SCL_OUT, MPR121_SDA_OUT, MPR121_SCL_EN, 
        MPR121_SDA_EN, ADS1292_SCLK, ADS1292_MISO, ADS1292_MOSI, ADS1292_DRDY, 
        ADS1292_RESET, ADS1292_START, ADS1292_CSN );
  input i_CLK, i_RSTN, UART_RXD, MPR121_SCL_IN, MPR121_SDA_IN, ADS1292_MISO,
         ADS1292_DRDY;
  output UART_TXD, MPR121_SCL_OUT, MPR121_SDA_OUT, MPR121_SCL_EN,
         MPR121_SDA_EN, ADS1292_SCLK, ADS1292_MOSI, ADS1292_RESET,
         ADS1292_START, ADS1292_CSN;
  wire   w_rstn, w_CLOCK_HALF, w_uart_data_tx_valid, w_uart_data_tx_ready,
         w_uart_data_rx_valid, w_mpr121_write_enable, w_mpr121_read_enable,
         w_mpr121_init_set, w_mpr121_busy, w_mpr121_fail, w_ads1292_init_set,
         w_ads1292_filtered_data_valid, w_ads1292_filtered_data_ack,
         w_ads1292_busy, w_ads1292_data_valid, n1, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8;
  wire   [55:0] w_uart_data_tx;
  wire   [15:0] w_uart_data_rx;
  wire   [7:0] w_mpr121_data_out;
  wire   [7:0] w_mpr121_reg_addr;
  wire   [7:0] w_mpr121_data_in;
  wire   [23:0] w_ads1292_filtered_data;
  wire   [2:0] w_ads1292_control;
  wire   [7:0] w_ads1292_reg_addr;
  wire   [7:0] w_ads1292_data_in;
  wire   [7:0] w_ads1292_reg_data_out;
  wire   [23:0] w_ads1292_data_out;

  async_rstn_glitch_synchronizer async_rstn_glitch_synchronizer ( .i_CLK(i_CLK), .i_RSTN(i_RSTN), .o_RSTN(w_rstn) );
  divider_by_2 divider_by_2 ( .i_CLK(i_CLK), .i_RSTN(w_rstn), .o_CLK_DIV_2(
        w_CLOCK_HALF) );
  uart_controller uart_controller ( .i_UART_DATA_TX({w_uart_data_tx[55:53], 
        1'b0, w_uart_data_tx[51:24], 1'b0, 1'b0, 1'b0, 1'b0, 
        w_uart_data_tx[19:7], 1'b0, w_uart_data_tx[5:3], 1'b0, 
        w_uart_data_tx[1:0]}), .i_UART_DATA_TX_VALID(w_uart_data_tx_valid), 
        .o_UART_DATA_TX_READY(w_uart_data_tx_ready), .o_UART_DATA_RX(
        w_uart_data_rx), .o_UART_DATA_RX_VALID(w_uart_data_rx_valid), 
        .i_CORE_BUSY(1'b0), .i_UART_RXD(UART_RXD), .o_UART_TXD(UART_TXD), 
        .i_CLK(w_CLOCK_HALF), .i_RSTN(n1) );
  sensor_core sensor_core ( .o_UART_DATA_TX({w_uart_data_tx[55:53], 
        SYNOPSYS_UNCONNECTED_1, w_uart_data_tx[51:24], SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        w_uart_data_tx[19:7], SYNOPSYS_UNCONNECTED_6, w_uart_data_tx[5:3], 
        SYNOPSYS_UNCONNECTED_7, w_uart_data_tx[1:0]}), .o_UART_DATA_TX_VALID(
        w_uart_data_tx_valid), .i_UART_DATA_TX_READY(w_uart_data_tx_ready), 
        .i_UART_DATA_RX(w_uart_data_rx), .i_UART_DATA_RX_VALID(
        w_uart_data_rx_valid), .i_MPR121_DATA_OUT(w_mpr121_data_out), 
        .o_MPR121_REG_ADDR(w_mpr121_reg_addr), .o_MPR121_DATA_IN({
        w_mpr121_data_in[7:6], SYNOPSYS_UNCONNECTED_8, w_mpr121_data_in[4:0]}), 
        .o_MPR121_WRITE_ENABLE(w_mpr121_write_enable), .o_MPR121_READ_ENABLE(
        w_mpr121_read_enable), .i_MPR121_INIT_SET(w_mpr121_init_set), 
        .i_MPR121_BUSY(w_mpr121_busy), .i_MPR121_FAIL(w_mpr121_fail), 
        .i_ADS1292_FILTERED_DATA_OUT(w_ads1292_filtered_data), 
        .o_ADS1292_CONTROL(w_ads1292_control), .o_ADS1292_REG_ADDR(
        w_ads1292_reg_addr), .o_ADS1292_DATA_IN(w_ads1292_data_in), 
        .i_ADS1292_REG_DATA_OUT(w_ads1292_reg_data_out), .i_ADS1292_INIT_SET(
        w_ads1292_init_set), .i_ADS1292_FILTERED_DATA_VALID(
        w_ads1292_filtered_data_valid), .o_ADS1292_FILTERED_DATA_ACK(
        w_ads1292_filtered_data_ack), .i_ADS1292_BUSY(w_ads1292_busy), .i_CLK(
        w_CLOCK_HALF), .i_RSTN(n1) );
  mpr121_controller mpr121_controller ( .o_MPR121_DATA_OUT(w_mpr121_data_out), 
        .o_MPR121_REG_ADDR(w_mpr121_reg_addr), .i_MPR121_DATA_IN({
        w_mpr121_data_in[7:6], 1'b0, w_mpr121_data_in[4:0]}), 
        .i_MPR121_WRITE_ENABLE(w_mpr121_write_enable), .i_MPR121_READ_ENABLE(
        w_mpr121_read_enable), .o_MPR121_INIT_SET(w_mpr121_init_set), 
        .o_MPR121_BUSY(w_mpr121_busy), .o_MPR121_FAIL(w_mpr121_fail), 
        .i_I2C_SCL_IN(MPR121_SCL_IN), .i_I2C_SDA_IN(MPR121_SDA_IN), 
        .o_I2C_SCL_OUT(MPR121_SCL_OUT), .o_I2C_SDA_OUT(MPR121_SDA_OUT), 
        .o_I2C_SCL_EN(MPR121_SCL_EN), .o_I2C_SDA_EN(MPR121_SDA_EN), .i_CLK(
        i_CLK), .i_RSTN(n1) );
  ads1292_filter ads1292_filter ( .i_ADS1292_DATA_OUT(w_ads1292_data_out), 
        .i_ADS1292_DATA_VALID(w_ads1292_data_valid), .o_ADS1292_FILTERED_DATA(
        w_ads1292_filtered_data), .o_ADS1292_FILTERED_DATA_VALID(
        w_ads1292_filtered_data_valid), .i_ADS1292_FILTERED_DATA_ACK(
        w_ads1292_filtered_data_ack), .i_CLK(i_CLK), .i_RSTN(w_rstn) );
  ads1292_controller ads1292_controller ( .o_ADS1292_DATA_OUT(
        w_ads1292_data_out), .i_ADS1292_CONTROL(w_ads1292_control), 
        .i_ADS1292_REG_ADDR(w_ads1292_reg_addr), .i_ADS1292_DATA_IN(
        w_ads1292_data_in), .o_ADS1292_REG_DATA_OUT(w_ads1292_reg_data_out), 
        .o_ADS1292_INIT_SET(w_ads1292_init_set), .o_ADS1292_DATA_VALID(
        w_ads1292_data_valid), .o_ADS1292_BUSY(w_ads1292_busy), .o_SPI_CLK(
        ADS1292_SCLK), .i_SPI_MISO(ADS1292_MISO), .o_SPI_MOSI(ADS1292_MOSI), 
        .i_ADS1292_DRDY(ADS1292_DRDY), .o_ADS1292_RESET(ADS1292_RESET), 
        .o_ADS1292_START(ADS1292_START), .o_SPI_CSN(ADS1292_CSN), .i_CLK(i_CLK), .i_RSTN(n1) );
  nid1_hd U1 ( .A(w_rstn), .Y(n1) );
endmodule


module khu_sensor_pad ( i_CLK, CLK_OUT, i_RSTN, UART_RXD, UART_TXD, MPR121_SCL, 
        MPR121_SDA, ADS1292_SCLK, ADS1292_MISO, ADS1292_MOSI, ADS1292_DRDY, 
        ADS1292_RESET, ADS1292_START, ADS1292_CSN );
  input i_CLK, i_RSTN, UART_RXD, ADS1292_MISO, ADS1292_DRDY;
  output CLK_OUT, UART_TXD, ADS1292_SCLK, ADS1292_MOSI, ADS1292_RESET,
         ADS1292_START, ADS1292_CSN;
  inout MPR121_SCL,  MPR121_SDA;
  wire   w_rstn_p, w_clk_p, n_2_net_, w_mpr121_scl_out_p, w_mpr121_scl_in_p,
         w_mpr121_scl_en_p, w_mpr121_sda_en_p, w_mpr121_sda_out_p,
         w_mpr121_sda_in_p, w_uart_rx_p, w_uart_tx_p, w_ads1292_sclk_p,
         w_ads1292_miso_p, w_ads1292_mosi_p, w_ads1292_drdy_p,
         w_ads1292_reset_p, w_ads1292_start_p, w_ads1292_csn_p, w_rstn, n1;

  vssoh pad1 (  );
  vssoh pad2 (  );
  vssoh pad3 (  );
  vdd33oph pad4 (  );
  vssoh pad5 (  );
  vssoh pad6 (  );
  vssoh pad7 (  );
  vssoh pad8 (  );
  vssoh pad9 (  );
  vssoh pad10 (  );
  vdd33oph pad11 (  );
  vssoh pad12 (  );
  vssoh pad13 (  );
  vssoh pad14 (  );
  vssoh pad15 (  );
  vssoh pad16 (  );
  phis pad17 ( .PAD(i_RSTN), .PI(1'b0), .Y(w_rstn_p) );
  vssoh pad18 (  );
  vssoh pad19 (  );
  vssiph pad20 (  );
  vssiph pad21 (  );
  vssiph pad22 (  );
  vdd12ih pad23 (  );
  vssiph pad24 (  );
  vssiph pad25 (  );
  vssiph pad26 (  );
  vssiph pad27 (  );
  vssiph pad28 (  );
  phsoscm3 pad29 ( .PADA(i_CLK), .E(1'b1), .PI(1'b0), .PADY(CLK_OUT), .YN(
        w_clk_p) );
  vssiph pad30 (  );
  vssiph pad31 (  );
  vssiph pad32 (  );
  vssiph pad33 (  );
  vssiph pad34 (  );
  vdd12ih pad35 (  );
  vssiph pad36 (  );
  vssiph pad37 (  );
  vssiph pad38 (  );
  vssoh pad39 (  );
  vssoh pad40 (  );
  vssoh pad41 (  );
  vdd33oph pad42 (  );
  vssoh pad43 (  );
  vssoh pad44 (  );
  vssoh pad45 (  );
  vssoh pad46 (  );
  vssoh pad47 (  );
  vssoh pad48 (  );
  vdd33oph pad49 (  );
  vssoh pad50 (  );
  vssoh pad51 (  );
  vssoh pad52 (  );
  vssoh pad53 (  );
  vssoh pad54 (  );
  vssoh pad55 (  );
  vdd33oph pad56 (  );
  vssoh pad57 (  );
  vssoh pad58 (  );
  vssoh pad59 (  );
  vssoh pad60 (  );
  vssoh pad61 (  );
  vssoh pad62 (  );
  vdd33oph pad63 (  );
  vssoh pad64 (  );
  vssoh pad65 (  );
  vssoh pad66 (  );
  vssoh pad68 (  );
  vssoh pad69 (  );
  phbct12 pad70 ( .TN(n_2_net_), .EN(1'b0), .A(w_mpr121_scl_out_p), .PI(1'b0), 
        .PAD(MPR121_SCL), .Y(w_mpr121_scl_in_p) );
  vssoh pad71 (  );
  vssoh pad72 (  );
  vssiph pad73 (  );
  vssiph pad74 (  );
  vssiph pad75 (  );
  vdd12ih_core pad76 (  );
  vssiph pad77 (  );
  vssiph pad78 (  );
  vssiph pad79 (  );
  vssoh pad80 (  );
  vssoh pad81 (  );
  phbct12 pad82 ( .TN(w_mpr121_sda_en_p), .EN(1'b0), .A(w_mpr121_sda_out_p), 
        .PI(1'b0), .PAD(MPR121_SDA), .Y(w_mpr121_sda_in_p) );
  vssoh pad83 (  );
  vssoh pad84 (  );
  vssiph pad85 (  );
  vssiph pad86 (  );
  vssiph pad87 (  );
  vdd12ih pad88 (  );
  vssiph pad89 (  );
  vssiph pad90 (  );
  vssiph pad91 (  );
  vssoh pad92 (  );
  vssoh pad93 (  );
  vssoh pad94 (  );
  vdd33oph pad95 (  );
  vssoh pad96 (  );
  vssoh pad97 (  );
  vssoh pad98 (  );
  vssoh pad99 (  );
  vssoh pad100 (  );
  vssoh pad101 (  );
  vdd33oph pad102 (  );
  vssoh pad103 (  );
  vssoh pad104 (  );
  vssoh pad105 (  );
  vssoh pad106 (  );
  vssoh pad107 (  );
  vdd33oph pad108 (  );
  vssoh pad109 (  );
  vssoh pad110 (  );
  vssoh pad111 (  );
  vssoh pad112 (  );
  vssoh pad113 (  );
  vssoh pad114 (  );
  vdd33oph pad115 (  );
  vssoh pad116 (  );
  vssoh pad117 (  );
  vssoh pad118 (  );
  vssoh pad119 (  );
  vssoh pad120 (  );
  phic pad121 ( .PAD(UART_RXD), .PI(1'b0), .Y(w_uart_rx_p) );
  vssoh pad122 (  );
  vssoh pad123 (  );
  vssiph pad124 (  );
  vssiph pad125 (  );
  vssiph pad126 (  );
  vdd12ih_core pad127 (  );
  vssiph pad128 (  );
  vssiph pad129 (  );
  vssiph pad130 (  );
  vssoh pad131 (  );
  vssoh pad132 (  );
  phob12 pad133 ( .A(n1), .PAD(UART_TXD) );
  vssoh pad134 (  );
  vssoh pad135 (  );
  vssiph pad136 (  );
  vssiph pad137 (  );
  vssiph pad138 (  );
  vdd12ih pad139 (  );
  vssiph pad140 (  );
  vssiph pad141 (  );
  vssiph pad142 (  );
  vssoh pad143 (  );
  vssoh pad144 (  );
  vssoh pad145 (  );
  vdd33oph pad146 (  );
  vssoh pad147 (  );
  vssoh pad148 (  );
  vssoh pad149 (  );
  vssoh pad150 (  );
  vssoh pad151 (  );
  vdd33oph pad152 (  );
  vssoh pad153 (  );
  vdd33oph pad154 (  );
  vssoh pad155 (  );
  vssoh pad156 (  );
  vssoh pad157 (  );
  vdd33oph pad158 (  );
  vssoh pad159 (  );
  vdd33oph pad160 (  );
  vssoh pad161 (  );
  vssoh pad162 (  );
  vssoh pad163 (  );
  vssoh pad164 (  );
  phob12 pad165 ( .A(w_ads1292_sclk_p), .PAD(ADS1292_SCLK) );
  vssoh pad166 (  );
  vssoh pad167 (  );
  vssoh pad168 (  );
  vssoh pad169 (  );
  vssoh pad170 (  );
  phic pad171 ( .PAD(ADS1292_MISO), .PI(1'b0), .Y(w_ads1292_miso_p) );
  vssoh pad172 (  );
  vssoh pad173 (  );
  vssoh pad174 (  );
  vssoh pad175 (  );
  phob12 pad176 ( .A(w_ads1292_mosi_p), .PAD(ADS1292_MOSI) );
  vssoh pad177 (  );
  vssoh pad178 (  );
  vssiph pad179 (  );
  vssiph pad180 (  );
  vdd12ih_core pad181 (  );
  vssiph pad182 (  );
  vssiph pad183 (  );
  vssoh pad184 (  );
  vssoh pad185 (  );
  phic pad186 ( .PAD(ADS1292_DRDY), .PI(1'b0), .Y(w_ads1292_drdy_p) );
  vssoh pad187 (  );
  vssoh pad188 (  );
  vssiph pad189 (  );
  vssiph pad190 (  );
  vdd12ih pad191 (  );
  vssiph pad192 (  );
  vssiph pad193 (  );
  vssoh pad194 (  );
  vssoh pad195 (  );
  phob12 pad196 ( .A(w_ads1292_reset_p), .PAD(ADS1292_RESET) );
  phob12 pad197 ( .A(w_ads1292_start_p), .PAD(ADS1292_START) );
  phob12 pad198 ( .A(w_ads1292_csn_p), .PAD(ADS1292_CSN) );
  vssoh pad199 (  );
  vssoh pad200 (  );
  vssoh pad201 (  );
  vdd33oph pad202 (  );
  vssoh pad203 (  );
  vssoh pad204 (  );
  vdd33oph pad205 (  );
  vdd33oph pad206 (  );
  vssoh pad207 (  );
  vssoh pad208 (  );
  async_rstn_glitch_synchronizer async_rstn_glitch_synchronizer ( .i_CLK(i_CLK), .i_RSTN(w_rstn_p), .o_RSTN(w_rstn) );
  khu_sensor_top khu_sensor_top ( .i_CLK(w_clk_p), .i_RSTN(w_rstn), .UART_RXD(
        w_uart_rx_p), .UART_TXD(w_uart_tx_p), .MPR121_SCL_IN(w_mpr121_scl_in_p), .MPR121_SDA_IN(w_mpr121_sda_in_p), .MPR121_SCL_OUT(w_mpr121_scl_out_p), 
        .MPR121_SDA_OUT(w_mpr121_sda_out_p), .MPR121_SCL_EN(w_mpr121_scl_en_p), 
        .MPR121_SDA_EN(w_mpr121_sda_en_p), .ADS1292_SCLK(w_ads1292_sclk_p), 
        .ADS1292_MISO(w_ads1292_miso_p), .ADS1292_MOSI(w_ads1292_mosi_p), 
        .ADS1292_DRDY(w_ads1292_drdy_p), .ADS1292_RESET(w_ads1292_reset_p), 
        .ADS1292_START(w_ads1292_start_p), .ADS1292_CSN(w_ads1292_csn_p) );
  nid6_hd U3 ( .A(w_uart_tx_p), .Y(n1) );
  ivd1_hd U4 ( .A(w_mpr121_scl_en_p), .Y(n_2_net_) );
endmodule

