module FIR_FILTER(
	input RESET,CLK,WR,
	input [15:0] iDATA,
	output [38:0] oDATA);


	reg [15:0] 	coef[0:18];	  
	reg [4:0] 	coef_cnt;	   
	reg [15:0] 	DATAFLOW[0:36];
	reg [16:0]	S0[0:18];
	reg [33:0] 	S1[0:18];
	reg [34:0]	S2[0:9];
	reg [35:0]	S3[0:4];
	reg [36:0]	S4[0:2];
	reg [37:0]	S5[0:1];
	reg [38:0]	S6;
	assign	oDATA = S6;
	always @ (posedge CLK or negedge RESET)		
		begin
			if(!RESET)
				begin
					coef_cnt<=0;
                                        coef[0]<=0;
                                        coef[1]<=0;
                                        coef[2]<=0;
                                        coef[3]<=0;
                                        coef[4]<=0;
                                        coef[5]<=0;
                                        coef[6]<=0;
                                        coef[7]<=0;
                                        coef[8]<=0;
                                        coef[9]<=0;
                                        coef[10]<=0;
                                        coef[11]<=0;
                                        coef[12]<=0;
                                        coef[13]<=0;
                                        coef[14]<=0;
                                        coef[15]<=0;
                                        coef[16]<=0;
                                        coef[17]<=0;
                                        coef[18]<=0;
					DATAFLOW[0]<=0;
					DATAFLOW[1]<=0;
					DATAFLOW[2]<=0;
					DATAFLOW[3]<=0;
					DATAFLOW[4]<=0;
					DATAFLOW[5]<=0;
					DATAFLOW[6]<=0;
					DATAFLOW[7]<=0;
					DATAFLOW[8]<=0;
					DATAFLOW[9]<=0;
					DATAFLOW[10]<=0;
					DATAFLOW[11]<=0;
					DATAFLOW[12]<=0;
					DATAFLOW[13]<=0;
					DATAFLOW[14]<=0;
					DATAFLOW[15]<=0;
					DATAFLOW[16]<=0;
					DATAFLOW[17]<=0;
					DATAFLOW[18]<=0;
					DATAFLOW[19]<=0;
					DATAFLOW[20]<=0;
					DATAFLOW[21]<=0;
					DATAFLOW[22]<=0;
					DATAFLOW[23]<=0;
					DATAFLOW[24]<=0;
					DATAFLOW[25]<=0;
					DATAFLOW[26]<=0;
					DATAFLOW[27]<=0;
					DATAFLOW[28]<=0;
					DATAFLOW[29]<=0;
					DATAFLOW[30]<=0;
					DATAFLOW[31]<=0;
					DATAFLOW[32]<=0;
					DATAFLOW[33]<=0;
					DATAFLOW[34]<=0;
					DATAFLOW[35]<=0;
				end
			else
				begin	
					if(WR)
						begin
							coef[coef_cnt]<=iDATA;
                		                        if(coef_cnt==18) coef_cnt<=0;
		                                        else coef_cnt<=coef_cnt+1;	
						end
					else
						begin
							DATAFLOW[0] <= iDATA;
		                                        DATAFLOW[1] <= DATAFLOW[0];
		                                        DATAFLOW[2] <= DATAFLOW[1];
		                                        DATAFLOW[3] <= DATAFLOW[2];
		                                        DATAFLOW[4] <= DATAFLOW[3];
		                                        DATAFLOW[5] <= DATAFLOW[4];
		                                        DATAFLOW[6] <= DATAFLOW[5];
		                                        DATAFLOW[7] <= DATAFLOW[6];
		                                        DATAFLOW[8] <= DATAFLOW[7];
		                                        DATAFLOW[9] <= DATAFLOW[8];
		                                        DATAFLOW[10] <= DATAFLOW[9];
		                                        DATAFLOW[11] <= DATAFLOW[10];
		                                        DATAFLOW[12] <= DATAFLOW[11];
		                                        DATAFLOW[13] <= DATAFLOW[12];
		                                        DATAFLOW[14] <= DATAFLOW[13];
		                                        DATAFLOW[15] <= DATAFLOW[14];
		                                        DATAFLOW[16] <= DATAFLOW[15];
		                                        DATAFLOW[17] <= DATAFLOW[16];
		                                        DATAFLOW[18] <= DATAFLOW[17];
		                                        DATAFLOW[19] <= DATAFLOW[18];
		                                        DATAFLOW[20] <= DATAFLOW[19];
		                                        DATAFLOW[21] <= DATAFLOW[20];
		                                        DATAFLOW[22] <= DATAFLOW[21];
		                                        DATAFLOW[23] <= DATAFLOW[22];
                		                        DATAFLOW[24] <= DATAFLOW[23];
		                                        DATAFLOW[25] <= DATAFLOW[24];
		                                        DATAFLOW[26] <= DATAFLOW[25];
		                                        DATAFLOW[27] <= DATAFLOW[26];
                                		        DATAFLOW[28] <= DATAFLOW[27];
                		                        DATAFLOW[29] <= DATAFLOW[28];
		                                        DATAFLOW[30] <= DATAFLOW[29];
                                		        DATAFLOW[31] <= DATAFLOW[30];
                		                        DATAFLOW[32] <= DATAFLOW[31];
		                                        DATAFLOW[33] <= DATAFLOW[32];
                                		        DATAFLOW[34] <= DATAFLOW[33];
                		                        DATAFLOW[35] <= DATAFLOW[34];
		                                        DATAFLOW[36] <= DATAFLOW[35];
							DATAFLOW[0] <= iDATA;
                		                        DATAFLOW[1] <= DATAFLOW[0];
        	                	                DATAFLOW[2] <= DATAFLOW[1];
	                                	        DATAFLOW[3] <= DATAFLOW[2];
                               		        	DATAFLOW[4] <= DATAFLOW[3];
                         	 	                DATAFLOW[5] <= DATAFLOW[4];
                	                	        DATAFLOW[6] <= DATAFLOW[5];
		        	                        DATAFLOW[7] <= DATAFLOW[6];	
		                                        DATAFLOW[8] <= DATAFLOW[7];
        	                                	DATAFLOW[9] <= DATAFLOW[8];
                	                	        DATAFLOW[10] <= DATAFLOW[9];
                        		                DATAFLOW[11] <= DATAFLOW[10];
        	                	                DATAFLOW[12] <= DATAFLOW[11];
	                                	        DATAFLOW[13] <= DATAFLOW[12];
                	                        	DATAFLOW[14] <= DATAFLOW[13];
	                                	        DATAFLOW[15] <= DATAFLOW[14];
        	                	                DATAFLOW[16] <= DATAFLOW[15];
                		                        DATAFLOW[17] <= DATAFLOW[16];
        	        	                        DATAFLOW[18] <= DATAFLOW[17];
	                        	                DATAFLOW[19] <= DATAFLOW[18];
                                        		DATAFLOW[20] <= DATAFLOW[19];
                                	        	DATAFLOW[21] <= DATAFLOW[20];
	                        	                DATAFLOW[22] <= DATAFLOW[21];
        	        	                        DATAFLOW[23] <= DATAFLOW[22];
        		                                DATAFLOW[24] <= DATAFLOW[23];
	                	                        DATAFLOW[25] <= DATAFLOW[24];
                                		        DATAFLOW[26] <= DATAFLOW[25];
                        	        	        DATAFLOW[27] <= DATAFLOW[26];
	                	                        DATAFLOW[28] <= DATAFLOW[27];
        		                                DATAFLOW[29] <= DATAFLOW[28];
	        	                                DATAFLOW[30] <= DATAFLOW[29];
                        	                	DATAFLOW[31] <= DATAFLOW[30];
                                		        DATAFLOW[32] <= DATAFLOW[31];
	                        	                DATAFLOW[33] <= DATAFLOW[32];
        	        	                        DATAFLOW[34] <= DATAFLOW[33];
        		                                DATAFLOW[35] <= DATAFLOW[34];
	                	                        DATAFLOW[36] <= DATAFLOW[35];
                                		        S0[0] <= DATAFLOW[0] + DATAFLOW[36];
                        	        	        S0[1] <= DATAFLOW[1] + DATAFLOW[35];
	                	                        S0[2] <= DATAFLOW[2] + DATAFLOW[34];
        		                                S0[3] <= DATAFLOW[3] + DATAFLOW[33];
	        	                                S0[4] <= DATAFLOW[4] + DATAFLOW[32];
                        	                	S0[5] <= DATAFLOW[5] + DATAFLOW[31];
							S0[6] <= DATAFLOW[6] + DATAFLOW[30];
							S0[7] <= DATAFLOW[7] + DATAFLOW[29];
							S0[8] <= DATAFLOW[8] + DATAFLOW[28];
							S0[9] <= DATAFLOW[9] + DATAFLOW[27];
							S0[10] <= DATAFLOW[10] + DATAFLOW[26];
							S0[11] <= DATAFLOW[11] + DATAFLOW[25];
							S0[12] <= DATAFLOW[12] + DATAFLOW[24];
							S0[13] <= DATAFLOW[13] + DATAFLOW[23];
							S0[14] <= DATAFLOW[14] + DATAFLOW[22];
							S0[15] <= DATAFLOW[15] + DATAFLOW[21];
							S0[16] <= DATAFLOW[16] + DATAFLOW[20];
							S0[17] <= DATAFLOW[17] + DATAFLOW[19];
							S0[18] <= DATAFLOW[18];
							S1[0] <= S0[0] * coef[0];
							S1[1] <= S0[1] * coef[1];
							S1[2] <= S0[2] * coef[2];
							S1[3] <= S0[3] * coef[3];
							S1[4] <= S0[4] * coef[4];
							S1[5] <= S0[5] * coef[5];
							S1[6] <= S0[6] * coef[6];
							S1[7] <= S0[7] * coef[7];
							S1[8] <= S0[8] * coef[8];
							S1[9] <= S0[9] * coef[9];
							S1[10] <= S0[10] * coef[10];
							S1[11] <= S0[11] * coef[11];
							S1[12] <= S0[12] * coef[12];
							S1[13] <= S0[13] * coef[13];
							S1[14] <= S0[14] * coef[14];
							S1[15] <= S0[15] * coef[15];
							S1[16] <= S0[16] * coef[16];
							S1[17] <= S0[17] * coef[17];	
							S1[18] <= S0[18] * coef[18];	
							S2[0] <= S1[0]+S1[1];
							S2[1] <= S1[2]+S1[3];
							S2[2] <= S1[4]+S1[5];
							S2[3] <= S1[6]+S1[7];
							S2[4] <= S1[8]+S1[9];
							S2[5] <= S1[10]+S1[11];
							S2[6] <= S1[12]+S1[13];
							S2[7] <= S1[14]+S1[15];
							S2[8] <= S1[16]+S1[17];
							S2[9] <= S1[18];		
							S3[0] <= S2[0]+S2[1];
							S3[1] <= S2[2]+S2[3];
							S3[2] <= S2[4]+S2[5];
							S3[3] <= S2[6]+S2[7];
							S3[4] <= S2[8]+S2[9];
							S4[0] <= S3[0]+S3[1];
							S4[1] <= S3[2]+S3[3];
							S4[2] <= S3[4];			
							S5[0] <= S4[0]+S4[1];
							S5[1] <= S4[2];
							S6    <= S5[0]+S5[1];
						end
				end					
		end	   	
endmodule
