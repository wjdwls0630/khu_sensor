
module converter_i2f ( i_A, i_A_STB, o_A_ACK, o_Z, o_Z_STB, i_Z_ACK, i_CLK, 
        i_RST );
  input [31:0] i_A;
  output [31:0] o_Z;
  input i_A_STB, i_Z_ACK, i_CLK, i_RST;
  output o_A_ACK, o_Z_STB;
  wire   z_s, N117, N166, N167, N168, N169, N170, N171, N172, N232, n13, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n222,
         n223, n224, n225, n226, n227, n228, n262, n597, n875, n876, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n181, n182, n183, n184, n185, n186, n187,
         n188, n213, n214, n215, n216, n217, n218, n219, n220, n221, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350;
  wire   [2:0] state;
  wire   [30:8] a;
  wire   [31:8] value;
  wire   [7:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U229 ( .A(i_RST), .Y(N232) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n4), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n4), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n4), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n4), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n4), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n4), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n228), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n228), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n4), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n4), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n4), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n4), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n4), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n4), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n4), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n4), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n4), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n4), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n4), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n4), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n4), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n228), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n228), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n228), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n4), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n4), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n4), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n4), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n4), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n4), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n4), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n4), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd z_reg_23_ ( .D(n597), .E(n5), .CK(i_CLK), .Q(z[23]) );
  fd1eqd1_hd z_reg_24_ ( .D(N166), .E(n5), .CK(i_CLK), .Q(z[24]) );
  fd1eqd1_hd z_reg_25_ ( .D(N167), .E(n5), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd z_reg_26_ ( .D(N168), .E(n5), .CK(i_CLK), .Q(z[26]) );
  fd1eqd1_hd z_reg_27_ ( .D(N169), .E(n5), .CK(i_CLK), .Q(z[27]) );
  fd1eqd1_hd z_reg_28_ ( .D(N170), .E(n5), .CK(i_CLK), .Q(z[28]) );
  fd1eqd1_hd z_reg_29_ ( .D(N171), .E(n227), .CK(i_CLK), .Q(z[29]) );
  fd1eqd1_hd z_reg_30_ ( .D(N172), .E(n227), .CK(i_CLK), .Q(z[30]) );
  fd1eqd1_hd z_s_reg ( .D(N117), .E(n876), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd z_reg_31_ ( .D(z_s), .E(n5), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd z_reg_0_ ( .D(z_m[0]), .E(n5), .CK(i_CLK), .Q(z[0]) );
  fd1eqd1_hd z_reg_1_ ( .D(z_m[1]), .E(n227), .CK(i_CLK), .Q(z[1]) );
  fd1eqd1_hd z_reg_2_ ( .D(z_m[2]), .E(n227), .CK(i_CLK), .Q(z[2]) );
  fd1eqd1_hd z_reg_3_ ( .D(z_m[3]), .E(n227), .CK(i_CLK), .Q(z[3]) );
  fd1eqd1_hd z_reg_4_ ( .D(z_m[4]), .E(n227), .CK(i_CLK), .Q(z[4]) );
  fd1eqd1_hd z_reg_5_ ( .D(z_m[5]), .E(n227), .CK(i_CLK), .Q(z[5]) );
  fd1eqd1_hd z_reg_6_ ( .D(z_m[6]), .E(n5), .CK(i_CLK), .Q(z[6]) );
  fd1eqd1_hd z_reg_7_ ( .D(z_m[7]), .E(n5), .CK(i_CLK), .Q(z[7]) );
  fd1eqd1_hd z_reg_8_ ( .D(z_m[8]), .E(n5), .CK(i_CLK), .Q(z[8]) );
  fd1eqd1_hd z_reg_9_ ( .D(z_m[9]), .E(n5), .CK(i_CLK), .Q(z[9]) );
  fd1eqd1_hd z_reg_10_ ( .D(z_m[10]), .E(n5), .CK(i_CLK), .Q(z[10]) );
  fd1eqd1_hd z_reg_11_ ( .D(z_m[11]), .E(n5), .CK(i_CLK), .Q(z[11]) );
  fd1eqd1_hd z_reg_12_ ( .D(z_m[12]), .E(n5), .CK(i_CLK), .Q(z[12]) );
  fd1eqd1_hd z_reg_13_ ( .D(z_m[13]), .E(n5), .CK(i_CLK), .Q(z[13]) );
  fd1eqd1_hd z_reg_14_ ( .D(z_m[14]), .E(n5), .CK(i_CLK), .Q(z[14]) );
  fd1eqd1_hd z_reg_15_ ( .D(z_m[15]), .E(n5), .CK(i_CLK), .Q(z[15]) );
  fd1eqd1_hd z_reg_16_ ( .D(z_m[16]), .E(n5), .CK(i_CLK), .Q(z[16]) );
  fd1eqd1_hd z_reg_17_ ( .D(z_m[17]), .E(n5), .CK(i_CLK), .Q(z[17]) );
  fd1eqd1_hd z_reg_18_ ( .D(z_m[18]), .E(n5), .CK(i_CLK), .Q(z[18]) );
  fd1eqd1_hd z_reg_19_ ( .D(z_m[19]), .E(n5), .CK(i_CLK), .Q(z[19]) );
  fd1eqd1_hd z_reg_20_ ( .D(z_m[20]), .E(n5), .CK(i_CLK), .Q(z[20]) );
  fd1eqd1_hd z_reg_21_ ( .D(z_m[21]), .E(n5), .CK(i_CLK), .Q(z[21]) );
  fd1eqd1_hd z_reg_22_ ( .D(z_m[22]), .E(n5), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd value_reg_30_ ( .D(n191), .CK(i_CLK), .Q(value[30]) );
  fd1qd1_hd value_reg_10_ ( .D(n211), .CK(i_CLK), .Q(value[10]) );
  fd1qd1_hd value_reg_31_ ( .D(n190), .CK(i_CLK), .Q(value[31]) );
  fd1qd1_hd value_reg_8_ ( .D(n1), .CK(i_CLK), .Q(value[8]) );
  fd1qd1_hd value_reg_12_ ( .D(n209), .CK(i_CLK), .Q(value[12]) );
  fd1qd1_hd value_reg_14_ ( .D(n207), .CK(i_CLK), .Q(value[14]) );
  fd1qd1_hd value_reg_16_ ( .D(n205), .CK(i_CLK), .Q(value[16]) );
  fd1qd1_hd value_reg_18_ ( .D(n203), .CK(i_CLK), .Q(value[18]) );
  fd1qd1_hd value_reg_20_ ( .D(n201), .CK(i_CLK), .Q(value[20]) );
  fd1qd1_hd value_reg_22_ ( .D(n199), .CK(i_CLK), .Q(value[22]) );
  fd1qd1_hd value_reg_24_ ( .D(n197), .CK(i_CLK), .Q(value[24]) );
  fd1qd1_hd value_reg_26_ ( .D(n195), .CK(i_CLK), .Q(value[26]) );
  fd1qd1_hd value_reg_28_ ( .D(n193), .CK(i_CLK), .Q(value[28]) );
  fd1qd1_hd value_reg_9_ ( .D(n212), .CK(i_CLK), .Q(value[9]) );
  fd1qd1_hd value_reg_11_ ( .D(n210), .CK(i_CLK), .Q(value[11]) );
  fd1qd1_hd value_reg_13_ ( .D(n208), .CK(i_CLK), .Q(value[13]) );
  fd1qd1_hd value_reg_15_ ( .D(n206), .CK(i_CLK), .Q(value[15]) );
  fd1qd1_hd value_reg_17_ ( .D(n204), .CK(i_CLK), .Q(value[17]) );
  fd1qd1_hd value_reg_19_ ( .D(n202), .CK(i_CLK), .Q(value[19]) );
  fd1qd1_hd value_reg_21_ ( .D(n200), .CK(i_CLK), .Q(value[21]) );
  fd1qd1_hd value_reg_23_ ( .D(n198), .CK(i_CLK), .Q(value[23]) );
  fd1qd1_hd value_reg_25_ ( .D(n196), .CK(i_CLK), .Q(value[25]) );
  fd1qd1_hd value_reg_27_ ( .D(n194), .CK(i_CLK), .Q(value[27]) );
  fd1qd1_hd value_reg_29_ ( .D(n192), .CK(i_CLK), .Q(value[29]) );
  fd1qd1_hd o_Z_STB_reg ( .D(n189), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_e_reg_4_ ( .D(n150), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n157), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n155), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n156), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_e_reg_0_ ( .D(n154), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd o_A_ACK_reg ( .D(n222), .CK(i_CLK), .Q(o_A_ACK) );
  fd1qd1_hd z_e_reg_3_ ( .D(n151), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n153), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n152), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n163), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n162), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n158), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n875), .CK(i_CLK), .Q(N117) );
  fd1qd1_hd z_m_reg_9_ ( .D(n171), .CK(i_CLK), .Q(z_m[9]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n875), .CK(i_CLK), .Q(a[30]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n226), .CK(i_CLK), .Q(z_m[23]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n875), .CK(i_CLK), .Q(a[29]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n175), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n167), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n170), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n172), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n168), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n164), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n160), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n173), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n169), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n165), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n161), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n174), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n166), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n159), .CK(i_CLK), .Q(z_m[21]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n875), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n875), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n875), .CK(i_CLK), .Q(a[24]) );
  fd1qd1_hd state_reg_2_ ( .D(n225), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_0_ ( .D(n224), .CK(i_CLK), .Q(state[0]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n875), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n875), .CK(i_CLK), .Q(a[25]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n180), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd state_reg_1_ ( .D(n223), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n176), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n177), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n179), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n178), .CK(i_CLK), .Q(z_m[2]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n875), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n875), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n875), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n875), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n875), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n875), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n875), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n875), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n875), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n875), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n875), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n875), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n875), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n875), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n875), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n875), .CK(i_CLK), .Q(a[8]) );
  ivd1_hd U435 ( .A(N232), .Y(n262) );
  clknd2d1_hd U231 ( .A(n35), .B(z_e[4]), .Y(n37) );
  clknd2d1_hd U232 ( .A(z_m[0]), .B(n345), .Y(n148) );
  clknd2d1_hd U233 ( .A(n16), .B(n188), .Y(n184) );
  clknd2d1_hd U234 ( .A(n139), .B(n345), .Y(n146) );
  clknd2d1_hd U235 ( .A(n345), .B(n214), .Y(n188) );
  clknd2d1_hd U236 ( .A(n332), .B(n339), .Y(n330) );
  clknd2d1_hd U237 ( .A(n876), .B(n15), .Y(n335) );
  clknd2d1_hd U238 ( .A(n65), .B(n345), .Y(n72) );
  clknd2d1_hd U239 ( .A(n83), .B(n345), .Y(n90) );
  clknd2d1_hd U240 ( .A(n101), .B(n345), .Y(n108) );
  clknd2d1_hd U241 ( .A(n119), .B(n345), .Y(n126) );
  clknd2d2_hd U242 ( .A(n130), .B(n16), .Y(n181) );
  clknd2d1_hd U243 ( .A(n28), .B(z_e[2]), .Y(n23) );
  clknd2d1_hd U244 ( .A(z_e[5]), .B(n41), .Y(n48) );
  clknd2d1_hd U245 ( .A(n876), .B(n39), .Y(n53) );
  clknd2d1_hd U246 ( .A(n130), .B(n39), .Y(n38) );
  clknd2d1_hd U247 ( .A(n47), .B(n24), .Y(n22) );
  clknd2d1_hd U248 ( .A(n39), .B(n323), .Y(n33) );
  clknd2d1_hd U249 ( .A(n235), .B(n237), .Y(n232) );
  clknd2d1_hd U250 ( .A(n243), .B(n245), .Y(n239) );
  clknd2d1_hd U251 ( .A(n251), .B(n253), .Y(n247) );
  clknd2d1_hd U252 ( .A(n259), .B(n261), .Y(n255) );
  clknd2d1_hd U253 ( .A(n268), .B(n270), .Y(n264) );
  clknd2d1_hd U254 ( .A(n276), .B(n278), .Y(n272) );
  clknd2d1_hd U255 ( .A(n284), .B(n286), .Y(n280) );
  clknd2d1_hd U256 ( .A(n292), .B(n294), .Y(n288) );
  clknd2d1_hd U257 ( .A(n300), .B(n302), .Y(n296) );
  clknd2d1_hd U258 ( .A(n308), .B(n310), .Y(n304) );
  clknd2d1_hd U259 ( .A(n231), .B(n219), .Y(n218) );
  clknd2d1_hd U260 ( .A(state[0]), .B(n339), .Y(n14) );
  clknd2d1_hd U261 ( .A(state[2]), .B(n327), .Y(n334) );
  clknd2d1_hd U262 ( .A(n10), .B(n49), .Y(n11) );
  clknd2d1_hd U263 ( .A(n8), .B(n18), .Y(n9) );
  clknd2d1_hd U264 ( .A(n6), .B(n27), .Y(n7) );
  clknd2d1_hd U265 ( .A(n183), .B(n182), .Y(n178) );
  clknd2d1_hd U266 ( .A(n187), .B(n186), .Y(n179) );
  clknd2d1_hd U267 ( .A(z_m[3]), .B(n143), .Y(n144) );
  clknd2d1_hd U268 ( .A(n3), .B(value[8]), .Y(n213) );
  clknd2d1_hd U269 ( .A(n338), .B(n331), .Y(n333) );
  clknd2d1_hd U270 ( .A(n60), .B(n63), .Y(n61) );
  clknd2d1_hd U271 ( .A(z_m[19]), .B(n69), .Y(n70) );
  clknd2d1_hd U272 ( .A(z_m[15]), .B(n87), .Y(n88) );
  clknd2d1_hd U273 ( .A(z_m[11]), .B(n105), .Y(n106) );
  clknd2d1_hd U274 ( .A(z_m[7]), .B(n123), .Y(n124) );
  clknd2d1_hd U275 ( .A(n96), .B(n99), .Y(n97) );
  clknd2d1_hd U276 ( .A(n134), .B(n137), .Y(n135) );
  clknd2d1_hd U277 ( .A(n114), .B(n117), .Y(n115) );
  clknd2d1_hd U278 ( .A(n78), .B(n81), .Y(n79) );
  clknd2d1_hd U279 ( .A(n28), .B(n27), .Y(n31) );
  clknd2d1_hd U280 ( .A(n35), .B(n18), .Y(n21) );
  clknd2d1_hd U281 ( .A(n25), .B(n22), .Y(n19) );
  clknd2d1_hd U282 ( .A(n234), .B(n233), .Y(n192) );
  clknd2d1_hd U283 ( .A(a[27]), .B(n239), .Y(n240) );
  clknd2d1_hd U284 ( .A(a[25]), .B(n247), .Y(n248) );
  clknd2d1_hd U285 ( .A(a[23]), .B(n255), .Y(n256) );
  clknd2d1_hd U286 ( .A(a[21]), .B(n264), .Y(n265) );
  clknd2d1_hd U287 ( .A(a[19]), .B(n272), .Y(n273) );
  clknd2d1_hd U288 ( .A(a[17]), .B(n280), .Y(n281) );
  clknd2d1_hd U289 ( .A(a[15]), .B(n288), .Y(n289) );
  clknd2d1_hd U290 ( .A(a[13]), .B(n296), .Y(n297) );
  clknd2d1_hd U291 ( .A(a[11]), .B(n304), .Y(n305) );
  clknd2d1_hd U292 ( .A(n315), .B(n314), .Y(n212) );
  clknd2d1_hd U293 ( .A(n318), .B(n317), .Y(n319) );
  clknd2d1_hd U294 ( .A(n230), .B(n229), .Y(n191) );
  ivd1_hd U295 ( .A(n16), .Y(n128) );
  clknd2d1_hd U296 ( .A(n215), .B(n335), .Y(n16) );
  nr2d1_hd U297 ( .A(a[29]), .B(n232), .Y(n231) );
  ad2d1_hd U298 ( .A(z_e[1]), .B(z_e[0]), .Y(n28) );
  scg2d1_hd U299 ( .A(a[8]), .B(n319), .C(value[8]), .D(n321), .Y(n1) );
  or2bd2_hd U300 ( .B(n15), .AN(n876), .Y(n321) );
  or2d1_hd U301 ( .A(n3), .B(n876), .Y(n323) );
  scg9d1_hd U302 ( .A(n4), .B(o_Z_STB), .C(n326), .Y(n189) );
  ivd2_hd U303 ( .A(n324), .Y(n875) );
  ad3d1_hd U304 ( .A(n228), .B(i_Z_ACK), .C(o_Z_STB), .Y(n217) );
  or2d1_hd U305 ( .A(n28), .B(n6), .Y(N166) );
  ad3d1_hd U306 ( .A(z_m[2]), .B(z_m[1]), .C(z_m[0]), .Y(n139) );
  nr2ad1_hd U307 ( .A(state[0]), .B(n334), .Y(n130) );
  nr2d2_hd U308 ( .A(n128), .B(n56), .Y(n343) );
  nr2d2_hd U309 ( .A(N117), .B(n321), .Y(n316) );
  ivd1_hd U310 ( .A(n321), .Y(n2) );
  ivd1_hd U311 ( .A(n181), .Y(n345) );
  nr2d1_hd U312 ( .A(a[27]), .B(n239), .Y(n235) );
  nr2d1_hd U313 ( .A(a[25]), .B(n247), .Y(n243) );
  nr2d1_hd U314 ( .A(a[23]), .B(n255), .Y(n251) );
  nr2d1_hd U315 ( .A(a[21]), .B(n264), .Y(n259) );
  nr2d1_hd U316 ( .A(a[19]), .B(n272), .Y(n268) );
  nr2d1_hd U317 ( .A(a[17]), .B(n280), .Y(n276) );
  nr2d1_hd U318 ( .A(a[15]), .B(n288), .Y(n284) );
  nr2d1_hd U319 ( .A(a[13]), .B(n296), .Y(n292) );
  nr2d1_hd U320 ( .A(a[11]), .B(n304), .Y(n300) );
  ivd1_hd U321 ( .A(n318), .Y(n320) );
  nr2d1_hd U322 ( .A(n56), .B(n36), .Y(n45) );
  ivd1_hd U323 ( .A(n39), .Y(n36) );
  nr2d1_hd U324 ( .A(n128), .B(n17), .Y(n39) );
  ivd1_hd U325 ( .A(n343), .Y(n147) );
  nr2d1_hd U326 ( .A(N117), .B(n218), .Y(n15) );
  ivd1_hd U327 ( .A(a[12]), .Y(n302) );
  ivd1_hd U328 ( .A(a[10]), .Y(n310) );
  nr2d1_hd U329 ( .A(a[9]), .B(a[8]), .Y(n308) );
  nr2d1_hd U330 ( .A(n3), .B(n216), .Y(n215) );
  ivd1_hd U331 ( .A(n336), .Y(n56) );
  nid2_hd U332 ( .A(n344), .Y(n3) );
  nr2d1_hd U333 ( .A(n327), .B(n330), .Y(n344) );
  ivd1_hd U334 ( .A(n130), .Y(n329) );
  nid2_hd U335 ( .A(n228), .Y(n4) );
  nd2d1_hd U336 ( .A(n876), .B(N117), .Y(n318) );
  nid2_hd U337 ( .A(n227), .Y(n5) );
  ivd1_hd U338 ( .A(a[30]), .Y(n219) );
  ivd1_hd U339 ( .A(a[28]), .Y(n237) );
  ivd1_hd U340 ( .A(a[26]), .Y(n245) );
  ivd1_hd U341 ( .A(a[24]), .Y(n253) );
  ivd1_hd U342 ( .A(a[22]), .Y(n261) );
  ivd1_hd U343 ( .A(a[20]), .Y(n270) );
  ivd1_hd U344 ( .A(a[18]), .Y(n278) );
  ivd1_hd U345 ( .A(a[16]), .Y(n286) );
  ivd1_hd U346 ( .A(a[14]), .Y(n294) );
  nr2d1_hd U347 ( .A(state[1]), .B(n14), .Y(n876) );
  nr2d1_hd U348 ( .A(z_m[23]), .B(n56), .Y(n216) );
  ivd1_hd U349 ( .A(state[2]), .Y(n339) );
  ivd1_hd U350 ( .A(state[1]), .Y(n327) );
  nr3d1_hd U351 ( .A(state[0]), .B(n339), .C(n327), .Y(n228) );
  nr2d1_hd U352 ( .A(n332), .B(n334), .Y(n227) );
  scg6d1_hd U353 ( .A(z_e[3]), .B(n7), .C(n8), .Y(N168) );
  scg6d1_hd U354 ( .A(z_e[5]), .B(n9), .C(n10), .Y(N170) );
  ivd1_hd U355 ( .A(z_e[0]), .Y(n597) );
  ivd1_hd U356 ( .A(z_m[23]), .Y(n349) );
  ivd1_hd U357 ( .A(n45), .Y(n55) );
  ivd1_hd U358 ( .A(z_e[6]), .Y(n49) );
  ivd1_hd U359 ( .A(z_e[4]), .Y(n18) );
  ivd1_hd U360 ( .A(z_e[2]), .Y(n27) );
  ivd1_hd U361 ( .A(z_m[21]), .Y(n63) );
  ivd1_hd U362 ( .A(z_m[22]), .Y(n342) );
  ivd1_hd U363 ( .A(z_m[17]), .Y(n81) );
  ivd1_hd U364 ( .A(z_m[13]), .Y(n99) );
  ivd1_hd U365 ( .A(z_m[9]), .Y(n117) );
  ivd1_hd U366 ( .A(z_m[5]), .Y(n137) );
  ivd1_hd U367 ( .A(state[0]), .Y(n332) );
  nr2d1_hd U368 ( .A(z_e[0]), .B(z_e[1]), .Y(n6) );
  nr2d1_hd U369 ( .A(n327), .B(n14), .Y(n336) );
  ivd1_hd U370 ( .A(a[8]), .Y(n313) );
  oa21d1_hd U371 ( .A(n6), .B(n27), .C(n7), .Y(N167) );
  nr2d1_hd U372 ( .A(z_e[3]), .B(n7), .Y(n8) );
  oa21d1_hd U373 ( .A(n8), .B(n18), .C(n9), .Y(N169) );
  nr2d1_hd U374 ( .A(z_e[5]), .B(n9), .Y(n10) );
  oa21d1_hd U375 ( .A(n10), .B(n49), .C(n11), .Y(N171) );
  ivd1_hd U376 ( .A(n11), .Y(n12) );
  ivd1_hd U377 ( .A(z_e[7]), .Y(n50) );
  ao22d1_hd U378 ( .A(n12), .B(n50), .C(z_e[7]), .D(n11), .Y(N172) );
  nr2d1_hd U379 ( .A(n349), .B(n56), .Y(n13) );
  nd3d1_hd U380 ( .A(n139), .B(z_m[3]), .C(z_m[4]), .Y(n129) );
  ivd1_hd U381 ( .A(z_m[6]), .Y(n127) );
  nr3d1_hd U382 ( .A(n129), .B(n137), .C(n127), .Y(n119) );
  nd3d1_hd U383 ( .A(n119), .B(z_m[7]), .C(z_m[8]), .Y(n110) );
  ivd1_hd U384 ( .A(z_m[10]), .Y(n109) );
  nr3d1_hd U385 ( .A(n110), .B(n117), .C(n109), .Y(n101) );
  nd3d1_hd U386 ( .A(n101), .B(z_m[11]), .C(z_m[12]), .Y(n92) );
  ivd1_hd U387 ( .A(z_m[14]), .Y(n91) );
  nr3d1_hd U388 ( .A(n92), .B(n99), .C(n91), .Y(n83) );
  nd3d1_hd U389 ( .A(n83), .B(z_m[15]), .C(z_m[16]), .Y(n74) );
  ivd1_hd U390 ( .A(z_m[18]), .Y(n73) );
  nr3d1_hd U391 ( .A(n74), .B(n81), .C(n73), .Y(n65) );
  nd3d1_hd U392 ( .A(n65), .B(z_m[19]), .C(z_m[20]), .Y(n57) );
  nr3d1_hd U393 ( .A(n342), .B(n63), .C(n57), .Y(n346) );
  ao21d1_hd U394 ( .A(n346), .B(z_m[23]), .C(n16), .Y(n17) );
  ivd1_hd U395 ( .A(z_e[3]), .Y(n24) );
  nr2d1_hd U396 ( .A(n23), .B(n24), .Y(n35) );
  ao21d1_hd U397 ( .A(n130), .B(n23), .C(n36), .Y(n25) );
  ivd1_hd U398 ( .A(n38), .Y(n47) );
  ao22d1_hd U399 ( .A(z_e[4]), .B(n19), .C(n45), .D(N169), .Y(n20) );
  oa211d1_hd U400 ( .A(n38), .B(n21), .C(n20), .D(n33), .Y(n150) );
  oa22d1_hd U401 ( .A(n25), .B(n24), .C(n23), .D(n22), .Y(n26) );
  scg17d1_hd U402 ( .A(n45), .B(N168), .C(n26), .D(n33), .Y(n151) );
  oa21d1_hd U403 ( .A(n28), .B(n329), .C(n39), .Y(n29) );
  ao22d1_hd U404 ( .A(z_e[2]), .B(n29), .C(n45), .D(N167), .Y(n30) );
  oa211d1_hd U405 ( .A(n38), .B(n31), .C(n30), .D(n33), .Y(n152) );
  ao22d1_hd U406 ( .A(n45), .B(N166), .C(z_e[1]), .D(n36), .Y(n32) );
  oa211d1_hd U407 ( .A(n38), .B(N166), .C(n32), .D(n33), .Y(n153) );
  oa21d1_hd U408 ( .A(n47), .B(n45), .C(n597), .Y(n34) );
  oa211d1_hd U409 ( .A(n39), .B(n597), .C(n34), .D(n33), .Y(n154) );
  nr2d1_hd U410 ( .A(n38), .B(n37), .Y(n41) );
  ao21d1_hd U411 ( .A(n130), .B(n37), .C(n36), .Y(n44) );
  oa21d1_hd U412 ( .A(z_e[5]), .B(n38), .C(n44), .Y(n46) );
  ao22d1_hd U413 ( .A(z_e[6]), .B(n46), .C(n45), .D(N171), .Y(n40) );
  oa211d1_hd U414 ( .A(z_e[6]), .B(n48), .C(n40), .D(n53), .Y(n155) );
  ivd1_hd U415 ( .A(z_e[5]), .Y(n43) );
  ao22d1_hd U416 ( .A(n45), .B(N170), .C(n41), .D(n43), .Y(n42) );
  oa211d1_hd U417 ( .A(n44), .B(n43), .C(n42), .D(n53), .Y(n156) );
  scg6d1_hd U418 ( .A(n49), .B(n47), .C(n46), .Y(n52) );
  nr2d1_hd U419 ( .A(n49), .B(n48), .Y(n51) );
  ao22d1_hd U420 ( .A(z_e[7]), .B(n52), .C(n51), .D(n50), .Y(n54) );
  oa211d1_hd U421 ( .A(n55), .B(N172), .C(n54), .D(n53), .Y(n157) );
  nr2d1_hd U422 ( .A(n57), .B(n181), .Y(n60) );
  ao21d1_hd U423 ( .A(n60), .B(n342), .C(n343), .Y(n59) );
  ao21d1_hd U424 ( .A(n130), .B(n57), .C(n128), .Y(n64) );
  oa21d1_hd U425 ( .A(z_m[21]), .B(n181), .C(n64), .Y(n341) );
  ao22d1_hd U426 ( .A(n3), .B(value[30]), .C(z_m[22]), .D(n341), .Y(n58) );
  oa21d1_hd U427 ( .A(n59), .B(n63), .C(n58), .Y(n158) );
  ao22d1_hd U428 ( .A(n3), .B(value[29]), .C(z_m[20]), .D(n343), .Y(n62) );
  oa211d1_hd U429 ( .A(n64), .B(n63), .C(n62), .D(n61), .Y(n159) );
  oa21d1_hd U430 ( .A(n65), .B(n329), .C(n16), .Y(n69) );
  scg20d1_hd U431 ( .A(n181), .B(z_m[19]), .C(n69), .Y(n68) );
  oa21d1_hd U432 ( .A(z_m[20]), .B(n72), .C(n147), .Y(n66) );
  ao22d1_hd U433 ( .A(n3), .B(value[28]), .C(z_m[19]), .D(n66), .Y(n67) );
  scg16d1_hd U434 ( .A(z_m[20]), .B(n68), .C(n67), .Y(n160) );
  ao22d1_hd U436 ( .A(n3), .B(value[27]), .C(z_m[18]), .D(n343), .Y(n71) );
  oa211d1_hd U437 ( .A(z_m[19]), .B(n72), .C(n71), .D(n70), .Y(n161) );
  nr2d1_hd U438 ( .A(n74), .B(n181), .Y(n78) );
  ao21d1_hd U439 ( .A(n78), .B(n73), .C(n343), .Y(n77) );
  ao21d1_hd U440 ( .A(n130), .B(n74), .C(n128), .Y(n82) );
  oa21d1_hd U441 ( .A(z_m[17]), .B(n181), .C(n82), .Y(n75) );
  ao22d1_hd U442 ( .A(n344), .B(value[26]), .C(z_m[18]), .D(n75), .Y(n76) );
  oa21d1_hd U443 ( .A(n77), .B(n81), .C(n76), .Y(n162) );
  ao22d1_hd U444 ( .A(n3), .B(value[25]), .C(z_m[16]), .D(n343), .Y(n80) );
  oa211d1_hd U445 ( .A(n82), .B(n81), .C(n80), .D(n79), .Y(n163) );
  oa21d1_hd U446 ( .A(n83), .B(n329), .C(n16), .Y(n87) );
  scg20d1_hd U447 ( .A(n181), .B(z_m[15]), .C(n87), .Y(n86) );
  oa21d1_hd U448 ( .A(z_m[16]), .B(n90), .C(n147), .Y(n84) );
  ao22d1_hd U449 ( .A(n344), .B(value[24]), .C(z_m[15]), .D(n84), .Y(n85) );
  scg16d1_hd U450 ( .A(z_m[16]), .B(n86), .C(n85), .Y(n164) );
  ao22d1_hd U451 ( .A(n3), .B(value[23]), .C(z_m[14]), .D(n343), .Y(n89) );
  oa211d1_hd U452 ( .A(z_m[15]), .B(n90), .C(n89), .D(n88), .Y(n165) );
  nr2d1_hd U453 ( .A(n92), .B(n181), .Y(n96) );
  ao21d1_hd U454 ( .A(n96), .B(n91), .C(n343), .Y(n95) );
  ao21d1_hd U455 ( .A(n130), .B(n92), .C(n128), .Y(n100) );
  oa21d1_hd U456 ( .A(z_m[13]), .B(n181), .C(n100), .Y(n93) );
  ao22d1_hd U457 ( .A(n344), .B(value[22]), .C(z_m[14]), .D(n93), .Y(n94) );
  oa21d1_hd U458 ( .A(n95), .B(n99), .C(n94), .Y(n166) );
  ao22d1_hd U459 ( .A(n3), .B(value[21]), .C(z_m[12]), .D(n343), .Y(n98) );
  oa211d1_hd U460 ( .A(n100), .B(n99), .C(n98), .D(n97), .Y(n167) );
  oa21d1_hd U461 ( .A(n101), .B(n329), .C(n16), .Y(n105) );
  scg20d1_hd U462 ( .A(n181), .B(z_m[11]), .C(n105), .Y(n104) );
  oa21d1_hd U463 ( .A(z_m[12]), .B(n108), .C(n147), .Y(n102) );
  ao22d1_hd U464 ( .A(n344), .B(value[20]), .C(z_m[11]), .D(n102), .Y(n103) );
  scg16d1_hd U465 ( .A(z_m[12]), .B(n104), .C(n103), .Y(n168) );
  ao22d1_hd U466 ( .A(n3), .B(value[19]), .C(z_m[10]), .D(n343), .Y(n107) );
  oa211d1_hd U467 ( .A(z_m[11]), .B(n108), .C(n107), .D(n106), .Y(n169) );
  nr2d1_hd U468 ( .A(n110), .B(n181), .Y(n114) );
  ao21d1_hd U469 ( .A(n114), .B(n109), .C(n343), .Y(n113) );
  ao21d1_hd U470 ( .A(n130), .B(n110), .C(n128), .Y(n118) );
  oa21d1_hd U471 ( .A(z_m[9]), .B(n181), .C(n118), .Y(n111) );
  ao22d1_hd U472 ( .A(n3), .B(value[18]), .C(z_m[10]), .D(n111), .Y(n112) );
  oa21d1_hd U473 ( .A(n113), .B(n117), .C(n112), .Y(n170) );
  ao22d1_hd U474 ( .A(n3), .B(value[17]), .C(z_m[8]), .D(n343), .Y(n116) );
  oa211d1_hd U475 ( .A(n118), .B(n117), .C(n116), .D(n115), .Y(n171) );
  oa21d1_hd U476 ( .A(n119), .B(n329), .C(n16), .Y(n123) );
  scg20d1_hd U477 ( .A(n181), .B(z_m[7]), .C(n123), .Y(n122) );
  oa21d1_hd U478 ( .A(z_m[8]), .B(n126), .C(n147), .Y(n120) );
  ao22d1_hd U479 ( .A(n344), .B(value[16]), .C(z_m[7]), .D(n120), .Y(n121) );
  scg16d1_hd U480 ( .A(z_m[8]), .B(n122), .C(n121), .Y(n172) );
  ao22d1_hd U481 ( .A(n3), .B(value[15]), .C(z_m[6]), .D(n343), .Y(n125) );
  oa211d1_hd U482 ( .A(z_m[7]), .B(n126), .C(n125), .D(n124), .Y(n173) );
  nr2d1_hd U483 ( .A(n129), .B(n181), .Y(n134) );
  ao21d1_hd U484 ( .A(n134), .B(n127), .C(n343), .Y(n133) );
  ao21d1_hd U485 ( .A(n130), .B(n129), .C(n128), .Y(n138) );
  oa21d1_hd U486 ( .A(z_m[5]), .B(n181), .C(n138), .Y(n131) );
  ao22d1_hd U487 ( .A(n3), .B(value[14]), .C(z_m[6]), .D(n131), .Y(n132) );
  oa21d1_hd U488 ( .A(n133), .B(n137), .C(n132), .Y(n174) );
  ao22d1_hd U489 ( .A(n344), .B(value[13]), .C(z_m[4]), .D(n343), .Y(n136) );
  oa211d1_hd U490 ( .A(n138), .B(n137), .C(n136), .D(n135), .Y(n175) );
  oa21d1_hd U491 ( .A(n139), .B(n329), .C(n16), .Y(n143) );
  scg20d1_hd U492 ( .A(n181), .B(z_m[3]), .C(n143), .Y(n142) );
  oa21d1_hd U493 ( .A(z_m[4]), .B(n146), .C(n147), .Y(n140) );
  ao22d1_hd U494 ( .A(n3), .B(value[12]), .C(z_m[3]), .D(n140), .Y(n141) );
  scg16d1_hd U495 ( .A(z_m[4]), .B(n142), .C(n141), .Y(n176) );
  ao22d1_hd U496 ( .A(n344), .B(value[11]), .C(z_m[2]), .D(n343), .Y(n145) );
  oa211d1_hd U497 ( .A(z_m[3]), .B(n146), .C(n145), .D(n144), .Y(n177) );
  oa21d1_hd U498 ( .A(z_m[2]), .B(n148), .C(n147), .Y(n149) );
  ao22d1_hd U499 ( .A(n3), .B(value[10]), .C(z_m[1]), .D(n149), .Y(n183) );
  ivd1_hd U500 ( .A(z_m[0]), .Y(n214) );
  nr2d1_hd U501 ( .A(z_m[1]), .B(n181), .Y(n185) );
  oa21d1_hd U502 ( .A(n184), .B(n185), .C(z_m[2]), .Y(n182) );
  ao22d1_hd U503 ( .A(n3), .B(value[9]), .C(z_m[1]), .D(n184), .Y(n187) );
  oa21d1_hd U504 ( .A(n343), .B(n185), .C(z_m[0]), .Y(n186) );
  oa211d1_hd U505 ( .A(n16), .B(n214), .C(n213), .D(n188), .Y(n180) );
  nr2d1_hd U506 ( .A(n217), .B(i_RST), .Y(n326) );
  oa22ad1_hd U507 ( .A(n218), .B(n318), .C(n321), .D(value[31]), .Y(n190) );
  nr2d1_hd U508 ( .A(n231), .B(n318), .Y(n220) );
  ao22d1_hd U509 ( .A(value[30]), .B(n321), .C(n220), .D(n219), .Y(n230) );
  ivd1_hd U510 ( .A(N117), .Y(n221) );
  oa211d1_hd U511 ( .A(n231), .B(n221), .C(n876), .D(a[30]), .Y(n229) );
  ao22d1_hd U512 ( .A(a[29]), .B(n316), .C(value[29]), .D(n321), .Y(n234) );
  scg17d1_hd U513 ( .A(a[29]), .B(n232), .C(n231), .D(n320), .Y(n233) );
  ao21d1_hd U514 ( .A(n235), .B(n320), .C(n316), .Y(n238) );
  nr2d1_hd U515 ( .A(n235), .B(n318), .Y(n241) );
  ao22d1_hd U516 ( .A(value[28]), .B(n321), .C(n241), .D(n237), .Y(n236) );
  oa21d1_hd U517 ( .A(n238), .B(n237), .C(n236), .Y(n193) );
  ao22d1_hd U518 ( .A(value[27]), .B(n321), .C(n241), .D(n240), .Y(n242) );
  scg14d1_hd U519 ( .A(a[27]), .B(n316), .C(n242), .Y(n194) );
  ao21d1_hd U520 ( .A(n243), .B(n320), .C(n316), .Y(n246) );
  nr2d1_hd U521 ( .A(n243), .B(n318), .Y(n249) );
  ao22d1_hd U522 ( .A(value[26]), .B(n321), .C(n249), .D(n245), .Y(n244) );
  oa21d1_hd U523 ( .A(n246), .B(n245), .C(n244), .Y(n195) );
  ao22d1_hd U524 ( .A(value[25]), .B(n321), .C(n249), .D(n248), .Y(n250) );
  scg14d1_hd U525 ( .A(a[25]), .B(n316), .C(n250), .Y(n196) );
  ao21d1_hd U526 ( .A(n251), .B(n320), .C(n316), .Y(n254) );
  nr2d1_hd U527 ( .A(n251), .B(n318), .Y(n257) );
  ao22d1_hd U528 ( .A(value[24]), .B(n321), .C(n257), .D(n253), .Y(n252) );
  oa21d1_hd U529 ( .A(n254), .B(n253), .C(n252), .Y(n197) );
  ao22d1_hd U530 ( .A(value[23]), .B(n321), .C(n257), .D(n256), .Y(n258) );
  scg14d1_hd U531 ( .A(a[23]), .B(n316), .C(n258), .Y(n198) );
  ao21d1_hd U532 ( .A(n259), .B(n320), .C(n316), .Y(n263) );
  nr2d1_hd U533 ( .A(n259), .B(n318), .Y(n266) );
  ao22d1_hd U534 ( .A(value[22]), .B(n321), .C(n266), .D(n261), .Y(n260) );
  oa21d1_hd U535 ( .A(n263), .B(n261), .C(n260), .Y(n199) );
  ao22d1_hd U536 ( .A(value[21]), .B(n321), .C(n266), .D(n265), .Y(n267) );
  scg14d1_hd U537 ( .A(a[21]), .B(n316), .C(n267), .Y(n200) );
  ao21d1_hd U538 ( .A(n268), .B(n320), .C(n316), .Y(n271) );
  nr2d1_hd U539 ( .A(n268), .B(n318), .Y(n274) );
  ao22d1_hd U540 ( .A(value[20]), .B(n321), .C(n274), .D(n270), .Y(n269) );
  oa21d1_hd U541 ( .A(n271), .B(n270), .C(n269), .Y(n201) );
  ao22d1_hd U542 ( .A(value[19]), .B(n321), .C(n274), .D(n273), .Y(n275) );
  scg14d1_hd U543 ( .A(a[19]), .B(n316), .C(n275), .Y(n202) );
  ao21d1_hd U544 ( .A(n276), .B(n320), .C(n316), .Y(n279) );
  nr2d1_hd U545 ( .A(n276), .B(n318), .Y(n282) );
  ao22d1_hd U546 ( .A(value[18]), .B(n321), .C(n282), .D(n278), .Y(n277) );
  oa21d1_hd U547 ( .A(n279), .B(n278), .C(n277), .Y(n203) );
  ao22d1_hd U548 ( .A(value[17]), .B(n321), .C(n282), .D(n281), .Y(n283) );
  scg14d1_hd U549 ( .A(a[17]), .B(n316), .C(n283), .Y(n204) );
  ao21d1_hd U550 ( .A(n284), .B(n320), .C(n316), .Y(n287) );
  nr2d1_hd U551 ( .A(n284), .B(n318), .Y(n290) );
  ao22d1_hd U552 ( .A(value[16]), .B(n321), .C(n290), .D(n286), .Y(n285) );
  oa21d1_hd U553 ( .A(n287), .B(n286), .C(n285), .Y(n205) );
  ao22d1_hd U554 ( .A(value[15]), .B(n321), .C(n290), .D(n289), .Y(n291) );
  scg14d1_hd U555 ( .A(a[15]), .B(n316), .C(n291), .Y(n206) );
  ao21d1_hd U556 ( .A(n292), .B(n320), .C(n316), .Y(n295) );
  nr2d1_hd U557 ( .A(n292), .B(n318), .Y(n298) );
  ao22d1_hd U558 ( .A(value[14]), .B(n321), .C(n298), .D(n294), .Y(n293) );
  oa21d1_hd U559 ( .A(n295), .B(n294), .C(n293), .Y(n207) );
  ao22d1_hd U560 ( .A(value[13]), .B(n321), .C(n298), .D(n297), .Y(n299) );
  scg14d1_hd U561 ( .A(a[13]), .B(n316), .C(n299), .Y(n208) );
  ao21d1_hd U562 ( .A(n300), .B(n320), .C(n316), .Y(n303) );
  nr2d1_hd U563 ( .A(n300), .B(n318), .Y(n306) );
  ao22d1_hd U564 ( .A(value[12]), .B(n321), .C(n306), .D(n302), .Y(n301) );
  oa21d1_hd U565 ( .A(n303), .B(n302), .C(n301), .Y(n209) );
  ao22d1_hd U566 ( .A(value[11]), .B(n321), .C(n306), .D(n305), .Y(n307) );
  scg14d1_hd U567 ( .A(a[11]), .B(n316), .C(n307), .Y(n210) );
  ao21d1_hd U568 ( .A(n308), .B(n320), .C(n316), .Y(n311) );
  nr2d1_hd U569 ( .A(n308), .B(n318), .Y(n312) );
  ao22d1_hd U570 ( .A(value[10]), .B(n321), .C(n312), .D(n310), .Y(n309) );
  oa21d1_hd U571 ( .A(n311), .B(n310), .C(n309), .Y(n211) );
  ao22d1_hd U572 ( .A(a[9]), .B(n316), .C(value[9]), .D(n321), .Y(n315) );
  scg16d1_hd U573 ( .A(a[9]), .B(n313), .C(n312), .Y(n314) );
  ivd1_hd U574 ( .A(n316), .Y(n317) );
  nr2d1_hd U575 ( .A(state[1]), .B(n330), .Y(n322) );
  nd3d1_hd U576 ( .A(n322), .B(i_A_STB), .C(o_A_ACK), .Y(n324) );
  scg21d1_hd U577 ( .A(n322), .B(o_A_ACK), .C(i_RST), .D(n875), .Y(n222) );
  nr3d1_hd U578 ( .A(n3), .B(n2), .C(n5), .Y(n328) );
  nr2d1_hd U579 ( .A(n13), .B(n323), .Y(n325) );
  nd4d1_hd U580 ( .A(n326), .B(n325), .C(n334), .D(n324), .Y(n338) );
  oa22d1_hd U581 ( .A(n262), .B(n328), .C(n327), .D(n338), .Y(n223) );
  nd3d1_hd U582 ( .A(n335), .B(n330), .C(n329), .Y(n331) );
  oa22d1_hd U583 ( .A(n262), .B(n333), .C(n338), .D(n332), .Y(n224) );
  scg15d1_hd U584 ( .A(n336), .B(n338), .C(n335), .D(n334), .Y(n337) );
  ivd1_hd U585 ( .A(n337), .Y(n340) );
  oa22d1_hd U586 ( .A(n262), .B(n340), .C(n339), .D(n338), .Y(n225) );
  ao21d1_hd U587 ( .A(n345), .B(n342), .C(n341), .Y(n350) );
  ao22d1_hd U588 ( .A(n344), .B(value[31]), .C(z_m[22]), .D(n343), .Y(n348) );
  nd3d1_hd U589 ( .A(n346), .B(n345), .C(n349), .Y(n347) );
  oa211d1_hd U590 ( .A(n350), .B(n349), .C(n348), .D(n347), .Y(n226) );
endmodule


module float_adder_3 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3, C91_DATA2_4,
         C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8, n1, n2, n27, n265,
         n266, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n509, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23,
         C2_Z_22, C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16,
         C2_Z_15, C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_43J4_124_6938_n58, DP_OP_43J4_124_6938_n57,
         DP_OP_43J4_124_6938_n56, DP_OP_43J4_124_6938_n55,
         DP_OP_43J4_124_6938_n54, DP_OP_43J4_124_6938_n53,
         DP_OP_43J4_124_6938_n52, DP_OP_43J4_124_6938_n51,
         DP_OP_43J4_124_6938_n50, DP_OP_43J4_124_6938_n49,
         DP_OP_43J4_124_6938_n48, DP_OP_43J4_124_6938_n47,
         DP_OP_43J4_124_6938_n46, DP_OP_43J4_124_6938_n45,
         DP_OP_43J4_124_6938_n44, DP_OP_43J4_124_6938_n43,
         DP_OP_43J4_124_6938_n42, DP_OP_43J4_124_6938_n41,
         DP_OP_43J4_124_6938_n40, DP_OP_43J4_124_6938_n39,
         DP_OP_43J4_124_6938_n38, DP_OP_43J4_124_6938_n37,
         DP_OP_43J4_124_6938_n36, DP_OP_43J4_124_6938_n35,
         DP_OP_43J4_124_6938_n34, DP_OP_43J4_124_6938_n33,
         DP_OP_43J4_124_6938_n32, DP_OP_43J4_124_6938_n27,
         DP_OP_43J4_124_6938_n26, DP_OP_43J4_124_6938_n25,
         DP_OP_43J4_124_6938_n24, DP_OP_43J4_124_6938_n23,
         DP_OP_43J4_124_6938_n22, DP_OP_43J4_124_6938_n21,
         DP_OP_43J4_124_6938_n20, DP_OP_43J4_124_6938_n19,
         DP_OP_43J4_124_6938_n18, DP_OP_43J4_124_6938_n17,
         DP_OP_43J4_124_6938_n16, DP_OP_43J4_124_6938_n15,
         DP_OP_43J4_124_6938_n14, DP_OP_43J4_124_6938_n13,
         DP_OP_43J4_124_6938_n12, DP_OP_43J4_124_6938_n11,
         DP_OP_43J4_124_6938_n10, DP_OP_43J4_124_6938_n9,
         DP_OP_43J4_124_6938_n8, DP_OP_43J4_124_6938_n7,
         DP_OP_43J4_124_6938_n6, DP_OP_43J4_124_6938_n5,
         DP_OP_43J4_124_6938_n4, DP_OP_43J4_124_6938_n3,
         DP_OP_43J4_124_6938_n2, DP_OP_43J4_124_6938_n1,
         DP_OP_154J4_137_6175_n9, DP_OP_154J4_137_6175_n8,
         DP_OP_154J4_137_6175_n7, DP_OP_154J4_137_6175_n6,
         DP_OP_154J4_137_6175_n5, DP_OP_154J4_137_6175_n4,
         DP_OP_154J4_137_6175_n3, DP_OP_154J4_137_6175_n2, n1282, n1283, n1286,
         n1287, n1311, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J4_137_6175_U10 ( .A(n1287), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J4_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J4_137_6175_U9 ( .A(n1287), .B(z_e[2]), .CI(
        DP_OP_154J4_137_6175_n9), .CO(DP_OP_154J4_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J4_137_6175_U8 ( .A(n1287), .B(z_e[3]), .CI(
        DP_OP_154J4_137_6175_n8), .CO(DP_OP_154J4_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J4_137_6175_U7 ( .A(n1287), .B(z_e[4]), .CI(
        DP_OP_154J4_137_6175_n7), .CO(DP_OP_154J4_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J4_137_6175_U6 ( .A(n1287), .B(z_e[5]), .CI(
        DP_OP_154J4_137_6175_n6), .CO(DP_OP_154J4_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J4_137_6175_U5 ( .A(n1287), .B(z_e[6]), .CI(
        DP_OP_154J4_137_6175_n5), .CO(DP_OP_154J4_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J4_137_6175_U4 ( .A(n1287), .B(z_e[7]), .CI(
        DP_OP_154J4_137_6175_n4), .CO(DP_OP_154J4_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J4_137_6175_U3 ( .A(n1287), .B(z_e[8]), .CI(
        DP_OP_154J4_137_6175_n3), .CO(DP_OP_154J4_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1581), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n509), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n509), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1581), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1581), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1581), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1581), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1581), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n1581), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n1581), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n1581), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n1581), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n1581), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n1581), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n1581), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n1581), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1581), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1581), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1581), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1581), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1581), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n509), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n509), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n509), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n509), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1581), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1581), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n1581), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1581), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1581), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1581), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n1571), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n1571), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n1571), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n1571), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n1570), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n1570), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n1571), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n1571), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n1571), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n1571), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n1571), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n1571), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n1571), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n1571), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n1571), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n1571), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n1571), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n1571), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n1571), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n1571), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n1571), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n1571), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n1571), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n1571), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n1571), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n1571), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n1571), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n1571), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n1571), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n1571), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n1571), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n1571), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n1571), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n1571), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n1571), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n1571), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n1571), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n1571), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n1571), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n1571), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n1571), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n1571), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n1571), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n1571), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n1571), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n1571), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n1571), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n1571), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n1571), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n1571), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n1571), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n1571), .CK(i_CLK), .Q(b[22]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n1570), .CK(i_CLK), .Q(sum[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n1570), .CK(i_CLK), .Q(sum[2]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n1570), .CK(i_CLK), .Q(sum[26]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n1570), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n1570), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n1570), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n1570), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n1570), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n1570), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n1570), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n1570), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n1570), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n1570), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n1570), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n1570), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n1570), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n1570), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n1570), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n1570), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n1570), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n1570), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n1570), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n1570), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n1570), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n1570), .CK(i_CLK), .Q(sum[25]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n1570), .CK(i_CLK), .Q(sum[1]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n1571), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n1571), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n1571), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n1571), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n1570), .CK(i_CLK), .Q(sum[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n1571), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n1571), .CK(i_CLK), .Q(b[28]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n1571), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n1571), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n1571), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n1571), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n1571), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n1571), .CK(i_CLK), .Q(b[26]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n1571), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n1571), .CK(i_CLK), .Q(b[23]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n265), .CK(i_CLK), .Q(guard) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1578), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1578), .CK(i_CLK), .Q(a_s) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n1286), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n1286), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J4_124_6938_U28 ( .A(C2_Z_0), .B(n1311), .CI(
        DP_OP_43J4_124_6938_n58), .CO(DP_OP_43J4_124_6938_n27), .S(N310) );
  fad1_hd DP_OP_43J4_124_6938_U27 ( .A(DP_OP_43J4_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J4_124_6938_n27), .CO(DP_OP_43J4_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J4_124_6938_U26 ( .A(DP_OP_43J4_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J4_124_6938_n26), .CO(DP_OP_43J4_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J4_124_6938_U25 ( .A(DP_OP_43J4_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J4_124_6938_n25), .CO(DP_OP_43J4_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J4_124_6938_U24 ( .A(DP_OP_43J4_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J4_124_6938_n24), .CO(DP_OP_43J4_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J4_124_6938_U23 ( .A(DP_OP_43J4_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J4_124_6938_n23), .CO(DP_OP_43J4_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J4_124_6938_U2 ( .A(DP_OP_43J4_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J4_124_6938_n2), .CO(DP_OP_43J4_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J4_124_6938_U3 ( .A(DP_OP_43J4_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J4_124_6938_n3), .CO(DP_OP_43J4_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J4_124_6938_U4 ( .A(DP_OP_43J4_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J4_124_6938_n4), .CO(DP_OP_43J4_124_6938_n3), .S(N334) );
  fad1_hd DP_OP_43J4_124_6938_U14 ( .A(DP_OP_43J4_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J4_124_6938_n14), .CO(DP_OP_43J4_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J4_124_6938_U15 ( .A(DP_OP_43J4_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J4_124_6938_n15), .CO(DP_OP_43J4_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J4_124_6938_U16 ( .A(DP_OP_43J4_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J4_124_6938_n16), .CO(DP_OP_43J4_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J4_124_6938_U17 ( .A(DP_OP_43J4_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J4_124_6938_n17), .CO(DP_OP_43J4_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J4_124_6938_U18 ( .A(DP_OP_43J4_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J4_124_6938_n18), .CO(DP_OP_43J4_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J4_124_6938_U19 ( .A(DP_OP_43J4_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J4_124_6938_n19), .CO(DP_OP_43J4_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J4_124_6938_U20 ( .A(DP_OP_43J4_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J4_124_6938_n20), .CO(DP_OP_43J4_124_6938_n19), .S(N318)
         );
  fad1_hd DP_OP_43J4_124_6938_U21 ( .A(DP_OP_43J4_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J4_124_6938_n21), .CO(DP_OP_43J4_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J4_124_6938_U22 ( .A(DP_OP_43J4_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J4_124_6938_n22), .CO(DP_OP_43J4_124_6938_n21), .S(N316)
         );
  fad1_hd DP_OP_43J4_124_6938_U13 ( .A(DP_OP_43J4_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J4_124_6938_n13), .CO(DP_OP_43J4_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J4_124_6938_U12 ( .A(DP_OP_43J4_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J4_124_6938_n12), .CO(DP_OP_43J4_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J4_124_6938_U11 ( .A(DP_OP_43J4_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J4_124_6938_n11), .CO(DP_OP_43J4_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J4_124_6938_U10 ( .A(DP_OP_43J4_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J4_124_6938_n10), .CO(DP_OP_43J4_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J4_124_6938_U9 ( .A(DP_OP_43J4_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J4_124_6938_n9), .CO(DP_OP_43J4_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J4_124_6938_U8 ( .A(DP_OP_43J4_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J4_124_6938_n8), .CO(DP_OP_43J4_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J4_124_6938_U7 ( .A(DP_OP_43J4_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J4_124_6938_n7), .CO(DP_OP_43J4_124_6938_n6), .S(N331) );
  fad1_hd DP_OP_43J4_124_6938_U6 ( .A(DP_OP_43J4_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J4_124_6938_n6), .CO(DP_OP_43J4_124_6938_n5), .S(N332) );
  fad1_hd DP_OP_43J4_124_6938_U5 ( .A(DP_OP_43J4_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J4_124_6938_n5), .CO(DP_OP_43J4_124_6938_n4), .S(N333) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  nr2d1_hd U523 ( .A(n1988), .B(n1932), .Y(n1949) );
  clknd2d1_hd U524 ( .A(b_m[5]), .B(n2081), .Y(n1588) );
  clknd2d1_hd U525 ( .A(n1596), .B(n1595), .Y(n1597) );
  clknd2d1_hd U526 ( .A(b_m[18]), .B(n1612), .Y(n1613) );
  clknd2d1_hd U527 ( .A(b_m[8]), .B(n2075), .Y(n1593) );
  clknd2d1_hd U528 ( .A(n1591), .B(b_m[7]), .Y(n1592) );
  clknd2d1_hd U529 ( .A(b_m[12]), .B(n2067), .Y(n1601) );
  clknd2d1_hd U530 ( .A(b_m[11]), .B(n1599), .Y(n1600) );
  clknd2d1_hd U531 ( .A(b_m[17]), .B(n2057), .Y(n1611) );
  clknd2d1_hd U532 ( .A(b_e[8]), .B(n2099), .Y(n1697) );
  clknd2d1_hd U533 ( .A(n1680), .B(n1679), .Y(n1688) );
  clknd2d1_hd U534 ( .A(b_e[6]), .B(n2097), .Y(n1679) );
  clknd2d1_hd U535 ( .A(a_e[9]), .B(n1683), .Y(n1700) );
  clknd2d1_hd U536 ( .A(b_m[19]), .B(n2053), .Y(n1614) );
  clknd2d1_hd U537 ( .A(n1717), .B(n1715), .Y(n1719) );
  clknd2d1_hd U538 ( .A(n1750), .B(n1792), .Y(n1716) );
  clknd2d1_hd U539 ( .A(n1700), .B(n1699), .Y(n1701) );
  clknd2d1_hd U540 ( .A(a_e[8]), .B(n2166), .Y(n1694) );
  clknd2d1_hd U541 ( .A(n2186), .B(n1701), .Y(n2232) );
  clknd2d1_hd U542 ( .A(n1705), .B(n1727), .Y(n2228) );
  clknd2d1_hd U543 ( .A(n1712), .B(n2094), .Y(n1715) );
  clknd2d1_hd U544 ( .A(n2160), .B(n1711), .Y(n1717) );
  clknd2d1_hd U545 ( .A(n1703), .B(z_e[1]), .Y(n1727) );
  clknd2d1_hd U546 ( .A(a_e[4]), .B(n2118), .Y(n2096) );
  clknd2d1_hd U547 ( .A(state[0]), .B(n2240), .Y(n2225) );
  clknd2d1_hd U548 ( .A(n1971), .B(guard), .Y(n1963) );
  clknd2d1_hd U549 ( .A(n1576), .B(n2186), .Y(n2249) );
  clknd2d1_hd U550 ( .A(n1718), .B(n2260), .Y(n1707) );
  clknd2d1_hd U551 ( .A(n1574), .B(n2186), .Y(n2091) );
  clknd2d1_hd U552 ( .A(n2185), .B(n2163), .Y(n2170) );
  clknd2d1_hd U553 ( .A(n2246), .B(n2240), .Y(n2243) );
  clknd2d1_hd U554 ( .A(n2202), .B(n2212), .Y(n2210) );
  clknd2d1_hd U555 ( .A(b_e[2]), .B(n2201), .Y(n2195) );
  clknd2d1_hd U556 ( .A(a_e[2]), .B(n2133), .Y(n2127) );
  clknd2d1_hd U557 ( .A(n2136), .B(n2128), .Y(n2126) );
  clknd2d1_hd U558 ( .A(n2136), .B(n2145), .Y(n2143) );
  clknd2d1_hd U559 ( .A(n2117), .B(n2095), .Y(n2103) );
  clknd2d1_hd U560 ( .A(n2177), .B(n2173), .Y(n2253) );
  clknd2d1_hd U561 ( .A(b_e[5]), .B(n2180), .Y(n2179) );
  clknd2d1_hd U562 ( .A(n2191), .B(b_e[4]), .Y(n2162) );
  clknd2d1_hd U563 ( .A(n2187), .B(b[28]), .Y(n2181) );
  clknd2d1_hd U564 ( .A(state[2]), .B(n2260), .Y(n2244) );
  clknd2d1_hd U565 ( .A(N41), .B(n2259), .Y(n2261) );
  clknd2d1_hd U566 ( .A(n1955), .B(n1946), .Y(n1937) );
  clknd2d1_hd U567 ( .A(n1942), .B(n1937), .Y(n1933) );
  clknd2d1_hd U568 ( .A(n1955), .B(n1918), .Y(n1925) );
  clknd2d1_hd U569 ( .A(z_m[21]), .B(n1964), .Y(n1957) );
  clknd2d1_hd U570 ( .A(n1972), .B(sum[27]), .Y(n1969) );
  clknd2d1_hd U571 ( .A(n1955), .B(n1893), .Y(n1900) );
  clknd2d1_hd U572 ( .A(n1955), .B(n1869), .Y(n1876) );
  clknd2d1_hd U573 ( .A(n1955), .B(n1967), .Y(n1827) );
  clknd2d1_hd U574 ( .A(n1955), .B(n1845), .Y(n1852) );
  clknd2d1_hd U575 ( .A(z_m[20]), .B(n1823), .Y(n1958) );
  clknd2d1_hd U576 ( .A(z_m[19]), .B(z_m[20]), .Y(n1813) );
  clknd2d1_hd U577 ( .A(n2190), .B(n2121), .Y(n1758) );
  clknd2d1_hd U578 ( .A(n2164), .B(n2097), .Y(n1743) );
  clknd2d1_hd U579 ( .A(b_e[0]), .B(a_e[0]), .Y(n1786) );
  clknd2d1_hd U580 ( .A(n1751), .B(n1750), .Y(n1779) );
  clknd2d1_hd U581 ( .A(n1778), .B(n1773), .Y(n1772) );
  clknd2d1_hd U582 ( .A(n1764), .B(n1760), .Y(n1759) );
  clknd2d1_hd U583 ( .A(b_e[7]), .B(a_e[7]), .Y(n1738) );
  clknd2d1_hd U584 ( .A(n1749), .B(n1745), .Y(n1744) );
  clknd2d1_hd U585 ( .A(n1796), .B(n1735), .Y(n1790) );
  clknd2d1_hd U586 ( .A(n1726), .B(n1725), .Y(n1729) );
  nid1_hd U587 ( .A(n1802), .Y(n1572) );
  clknd2d1_hd U588 ( .A(state[1]), .B(n2246), .Y(n2222) );
  clknd2d1_hd U589 ( .A(state[3]), .B(n1718), .Y(n2221) );
  clknd2d1_hd U590 ( .A(a[23]), .B(a[24]), .Y(n2147) );
  clknd2d1_hd U591 ( .A(n2134), .B(a[26]), .Y(n2130) );
  clknd2d1_hd U592 ( .A(b[23]), .B(b[24]), .Y(n2214) );
  clknd2d1_hd U593 ( .A(n2213), .B(n2210), .Y(n2206) );
  clknd2d1_hd U594 ( .A(a_e[5]), .B(n2112), .Y(n2111) );
  clknd2d1_hd U595 ( .A(n2119), .B(a[28]), .Y(n2113) );
  clknd2d1_hd U596 ( .A(b_e[4]), .B(n2202), .Y(n2194) );
  clknd2d1_hd U597 ( .A(n2203), .B(b[26]), .Y(n2198) );
  clknd2d1_hd U598 ( .A(n1808), .B(n1807), .Y(n393) );
  clknd2d1_hd U599 ( .A(n1580), .B(n2167), .Y(n2172) );
  clknd2d1_hd U600 ( .A(n2200), .B(n2199), .Y(n495) );
  clknd2d1_hd U601 ( .A(a[30]), .B(n2100), .Y(n2105) );
  clknd2d1_hd U602 ( .A(n2181), .B(n2174), .Y(n2176) );
  clknd2d1_hd U603 ( .A(n1956), .B(n1937), .Y(n1939) );
  clknd2d1_hd U604 ( .A(n1993), .B(n1992), .Y(n428) );
  clknd2d1_hd U605 ( .A(DP_OP_154J4_137_6175_n2), .B(n1991), .Y(n1989) );
  clknd2d1_hd U606 ( .A(n1970), .B(n1805), .Y(n265) );
  clknd2d1_hd U607 ( .A(n1789), .B(n1741), .Y(n362) );
  clknd2d1_hd U608 ( .A(n2136), .B(n2133), .Y(n2142) );
  clknd2d1_hd U609 ( .A(n2136), .B(n2118), .Y(n2125) );
  clknd2d1_hd U610 ( .A(n2202), .B(n2201), .Y(n2209) );
  clknd2d1_hd U611 ( .A(n2113), .B(n2106), .Y(n2107) );
  ad2d4_hd U612 ( .A(n1311), .B(n1627), .Y(n1568) );
  ivd4_hd U613 ( .A(n1568), .Y(n1569) );
  ivd2_hd U614 ( .A(n1791), .Y(n1311) );
  ivd1_hd U615 ( .A(b_m[1]), .Y(n2040) );
  ivd1_hd U616 ( .A(b_m[2]), .Y(n2039) );
  ivd1_hd U617 ( .A(b_m[23]), .Y(n1997) );
  nr2d4_hd U618 ( .A(n1568), .B(n1791), .Y(n1655) );
  oa21d1_hd U619 ( .A(n1624), .B(n1623), .C(n1622), .Y(n1625) );
  ao21d1_hd U620 ( .A(a_m[23]), .B(n1997), .C(n1621), .Y(n1624) );
  ivd3_hd U621 ( .A(n1282), .Y(n1570) );
  ivd1_hd U622 ( .A(b_m[26]), .Y(n2250) );
  xo2d1_hd U623 ( .A(n1311), .B(DP_OP_43J4_124_6938_n1), .Y(N337) );
  nid6_hd U624 ( .A(n27), .Y(n1571) );
  ad3d1_hd U625 ( .A(n2220), .B(i_AB_STB), .C(o_AB_ACK), .Y(n27) );
  or2d2_hd U626 ( .A(n1707), .B(n2225), .Y(n1283) );
  scg9d1_hd U627 ( .A(n2238), .B(n1701), .C(n1283), .Y(n2158) );
  scg2d1_hd U628 ( .A(b_e[9]), .B(n1698), .C(n1697), .D(n1696), .Y(n1699) );
  ad3d1_hd U629 ( .A(n2258), .B(n1577), .C(n2256), .Y(n2262) );
  ivd2_hd U630 ( .A(n1779), .Y(n1804) );
  ivd2_hd U631 ( .A(n1969), .Y(n1943) );
  or4d1_hd U632 ( .A(z_m[23]), .B(z_e[0]), .C(n1728), .D(n1727), .Y(n1735) );
  or2d1_hd U633 ( .A(n2243), .B(n2244), .Y(n1282) );
  or4d1_hd U634 ( .A(n1678), .B(a_e[9]), .C(a_e[0]), .D(a_e[8]), .Y(n1792) );
  oa22d4_hd U635 ( .A(n1657), .B(n1709), .C(a_s), .D(b_s), .Y(n1791) );
  or2d1_hd U636 ( .A(b_e[2]), .B(a_e[2]), .Y(n1771) );
  ivd1_hd U637 ( .A(b_m[0]), .Y(n2041) );
  nr2d2_hd U638 ( .A(n1797), .B(n2224), .Y(n1803) );
  ivd2_hd U639 ( .A(n1949), .Y(n1956) );
  nr2ad1_hd U640 ( .A(n1973), .B(n1986), .Y(n1990) );
  nr2ad1_hd U641 ( .A(n2256), .B(n1932), .Y(n1938) );
  nr2ad1_hd U642 ( .A(n2222), .B(n2244), .Y(n1287) );
  oa22ad1_hd U643 ( .A(n1590), .B(a_m[6]), .C(n1589), .D(b_m[6]), .Y(n1591) );
  ivd1_hd U644 ( .A(b_m[3]), .Y(n2038) );
  ivd1_hd U645 ( .A(b_m[4]), .Y(n2035) );
  ao22d1_hd U646 ( .A(a_m[26]), .B(n2250), .C(n1626), .D(n1625), .Y(n1627) );
  ivd1_hd U647 ( .A(a_m[3]), .Y(n2086) );
  ivd1_hd U648 ( .A(a_m[5]), .Y(n2081) );
  ivd1_hd U649 ( .A(b_m[5]), .Y(n2033) );
  nid2_hd U650 ( .A(n2257), .Y(n1577) );
  ivd1_hd U651 ( .A(n1955), .Y(n1931) );
  ivd1_hd U652 ( .A(n1984), .Y(n1986) );
  ivd1_hd U653 ( .A(n2093), .Y(n1575) );
  oa21d1_hd U654 ( .A(a_m[21]), .B(n2001), .C(n1618), .Y(n1619) );
  ivd1_hd U655 ( .A(a_m[4]), .Y(n2083) );
  ivd1_hd U656 ( .A(n1787), .Y(n1800) );
  ivd1_hd U657 ( .A(n1283), .Y(n1578) );
  nr2d1_hd U658 ( .A(n2258), .B(n1932), .Y(n1955) );
  ivd1_hd U659 ( .A(n1971), .Y(n2258) );
  nid2_hd U660 ( .A(n1944), .Y(n1573) );
  ivd1_hd U661 ( .A(n1938), .Y(n1945) );
  nr2d1_hd U662 ( .A(n2221), .B(n2243), .Y(n1971) );
  ivd1_hd U663 ( .A(n1287), .Y(n1988) );
  ivd2_hd U664 ( .A(n2158), .Y(n1576) );
  ivd2_hd U665 ( .A(n1575), .Y(n1574) );
  ivd1_hd U666 ( .A(n1286), .Y(n2223) );
  ivd1_hd U667 ( .A(n2238), .Y(n2186) );
  nd2bd1_hd U668 ( .AN(n1707), .B(n2234), .Y(n2238) );
  ivd1_hd U669 ( .A(b_m[24]), .Y(n1995) );
  ivd1_hd U670 ( .A(a_m[16]), .Y(n2059) );
  ivd1_hd U671 ( .A(b_m[10]), .Y(n2023) );
  ivd1_hd U672 ( .A(b_m[13]), .Y(n2017) );
  ivd1_hd U673 ( .A(a_m[15]), .Y(n2061) );
  ivd1_hd U674 ( .A(b_m[14]), .Y(n2015) );
  ivd1_hd U675 ( .A(a_m[17]), .Y(n2057) );
  ivd1_hd U676 ( .A(b_m[17]), .Y(n2009) );
  ivd1_hd U677 ( .A(b_m[21]), .Y(n2001) );
  nid2_hd U678 ( .A(n509), .Y(n1581) );
  nr3d1_hd U679 ( .A(n1751), .B(n1717), .C(n1716), .Y(n1802) );
  ivd1_hd U680 ( .A(n1715), .Y(n1751) );
  ivd2_hd U681 ( .A(n2249), .Y(n2036) );
  scg20d2_hd U682 ( .A(n1812), .B(n1963), .C(n265), .Y(n1932) );
  ivd1_hd U683 ( .A(n1972), .Y(n1805) );
  ivd2_hd U684 ( .A(n1283), .Y(n1579) );
  ivd2_hd U685 ( .A(n2091), .Y(n2084) );
  nr2d1_hd U686 ( .A(n2225), .B(n2244), .Y(n1972) );
  nd2bd1_hd U687 ( .AN(n2244), .B(n2234), .Y(n2256) );
  ivd1_hd U688 ( .A(n2202), .Y(n2252) );
  nr2d1_hd U689 ( .A(n2218), .B(n2238), .Y(n2202) );
  ao21d1_hd U690 ( .A(n2160), .B(n2159), .C(n1576), .Y(n2218) );
  ivd1_hd U691 ( .A(n1283), .Y(n1580) );
  ivd1_hd U692 ( .A(n2136), .Y(n2154) );
  nr2d1_hd U693 ( .A(n2151), .B(n2238), .Y(n2136) );
  ao21d1_hd U694 ( .A(n2094), .B(n2159), .C(n1574), .Y(n2151) );
  scg16d1_hd U695 ( .A(n2233), .B(n2232), .C(n1283), .Y(n2093) );
  ivd1_hd U696 ( .A(b_e[1]), .Y(n2212) );
  nr2d1_hd U697 ( .A(n1719), .B(n1716), .Y(n2159) );
  nr2d1_hd U698 ( .A(n1707), .B(n2222), .Y(n1286) );
  ivd1_hd U699 ( .A(b_e[6]), .Y(n2164) );
  ivd1_hd U700 ( .A(a_e[8]), .Y(n2099) );
  ivd1_hd U701 ( .A(a_e[5]), .Y(n2116) );
  ivd1_hd U702 ( .A(a_e[6]), .Y(n2097) );
  nr2d1_hd U703 ( .A(n2246), .B(n2240), .Y(n2234) );
  ivd1_hd U704 ( .A(state[0]), .Y(n2246) );
  ivd1_hd U705 ( .A(state[1]), .Y(n2240) );
  ivd1_hd U706 ( .A(state[3]), .Y(n2260) );
  ivd1_hd U707 ( .A(b_m[25]), .Y(n1629) );
  ivd1_hd U708 ( .A(b_m[19]), .Y(n2005) );
  ivd1_hd U709 ( .A(b_m[20]), .Y(n2003) );
  ivd1_hd U710 ( .A(a_m[20]), .Y(n2051) );
  ivd1_hd U711 ( .A(b_m[22]), .Y(n1999) );
  ivd1_hd U712 ( .A(a_m[22]), .Y(n2047) );
  ivd1_hd U713 ( .A(a_m[25]), .Y(n1668) );
  ivd1_hd U714 ( .A(n2159), .Y(n2242) );
  nr2d1_hd U715 ( .A(n2222), .B(n2221), .Y(n509) );
  ivd1_hd U716 ( .A(n1796), .Y(n2224) );
  ivd1_hd U717 ( .A(z_m[1]), .Y(n1946) );
  ao21d1_hd U718 ( .A(n1796), .B(n1797), .C(n1734), .Y(n1789) );
  ivd1_hd U719 ( .A(n1710), .Y(n1793) );
  nr2d1_hd U720 ( .A(n2225), .B(n2221), .Y(n1796) );
  ivd1_hd U721 ( .A(z_m[20]), .Y(n1832) );
  ivd1_hd U722 ( .A(z_m[21]), .Y(n1826) );
  ivd1_hd U723 ( .A(n1932), .Y(n1952) );
  ivd1_hd U724 ( .A(z_m[22]), .Y(n1965) );
  ivd1_hd U725 ( .A(z_m[17]), .Y(n1850) );
  ivd1_hd U726 ( .A(z_m[18]), .Y(n1838) );
  ivd1_hd U727 ( .A(z_m[13]), .Y(n1874) );
  ivd1_hd U728 ( .A(z_m[14]), .Y(n1862) );
  ivd1_hd U729 ( .A(z_m[10]), .Y(n1886) );
  ivd1_hd U730 ( .A(z_m[9]), .Y(n1898) );
  ivd1_hd U731 ( .A(z_m[5]), .Y(n1923) );
  ivd1_hd U732 ( .A(z_m[6]), .Y(n1910) );
  ivd1_hd U733 ( .A(z_m[23]), .Y(n1964) );
  ivd1_hd U734 ( .A(z_e[8]), .Y(n1975) );
  ivd1_hd U735 ( .A(z_e[7]), .Y(n1733) );
  ivd1_hd U736 ( .A(z_e[0]), .Y(n1985) );
  ivd1_hd U737 ( .A(n2254), .Y(n2207) );
  nr2d1_hd U738 ( .A(n2223), .B(n2218), .Y(n2254) );
  ivd1_hd U739 ( .A(b[30]), .Y(n2173) );
  ivd1_hd U740 ( .A(n2156), .Y(n2140) );
  nr2d1_hd U741 ( .A(n2223), .B(n2151), .Y(n2156) );
  ivd1_hd U742 ( .A(a_e[7]), .Y(n2101) );
  ivd1_hd U743 ( .A(a_e[4]), .Y(n2121) );
  ivd1_hd U744 ( .A(a_e[2]), .Y(n2137) );
  ivd1_hd U745 ( .A(b_e[7]), .Y(n2168) );
  nr3d1_hd U746 ( .A(n1676), .B(n1675), .C(n1674), .Y(n1712) );
  ivd1_hd U747 ( .A(b_e[9]), .Y(n1683) );
  ivd1_hd U748 ( .A(b_e[0]), .Y(n2211) );
  ivd1_hd U749 ( .A(b_e[5]), .Y(n2184) );
  ivd1_hd U750 ( .A(b_e[8]), .Y(n2166) );
  ivd1_hd U751 ( .A(a_e[0]), .Y(n2144) );
  ivd1_hd U752 ( .A(a_e[1]), .Y(n2145) );
  ivd1_hd U753 ( .A(a_e[3]), .Y(n2128) );
  ivd1_hd U754 ( .A(state[2]), .Y(n1718) );
  ivd1_hd U755 ( .A(a_m[1]), .Y(n2088) );
  ivd1_hd U756 ( .A(a_m[2]), .Y(n2087) );
  ivd1_hd U757 ( .A(a_m[6]), .Y(n2079) );
  ivd1_hd U758 ( .A(b_m[6]), .Y(n2031) );
  ivd1_hd U759 ( .A(a_m[7]), .Y(n2077) );
  ivd1_hd U760 ( .A(b_m[7]), .Y(n2029) );
  ivd1_hd U761 ( .A(a_m[11]), .Y(n2069) );
  ivd1_hd U762 ( .A(b_m[11]), .Y(n2021) );
  ivd1_hd U763 ( .A(a_m[13]), .Y(n2065) );
  ivd1_hd U764 ( .A(a_m[14]), .Y(n2063) );
  ivd1_hd U765 ( .A(a_m[18]), .Y(n2055) );
  ivd1_hd U766 ( .A(b_m[18]), .Y(n2007) );
  ivd1_hd U767 ( .A(a_m[21]), .Y(n2049) );
  ivd1_hd U768 ( .A(a_m[23]), .Y(n2045) );
  ivd1_hd U769 ( .A(a_m[24]), .Y(n2043) );
  ivd1_hd U770 ( .A(a_m[19]), .Y(n2053) );
  ivd1_hd U771 ( .A(b_m[15]), .Y(n2013) );
  ivd1_hd U772 ( .A(b_m[16]), .Y(n2011) );
  ivd1_hd U773 ( .A(a_m[12]), .Y(n2067) );
  ivd1_hd U774 ( .A(a_m[8]), .Y(n2075) );
  ivd1_hd U775 ( .A(b_m[8]), .Y(n2027) );
  ivd1_hd U776 ( .A(b_m[9]), .Y(n2025) );
  ivd1_hd U777 ( .A(a_m[10]), .Y(n2071) );
  ivd1_hd U778 ( .A(a_m[9]), .Y(n2073) );
  ivd1_hd U779 ( .A(b_m[12]), .Y(n2019) );
  ivd1_hd U780 ( .A(a_m[26]), .Y(n2092) );
  ivd1_hd U781 ( .A(a_s), .Y(n1709) );
  ivd1_hd U782 ( .A(b_s), .Y(n1657) );
  ivd1_hd U783 ( .A(z_m[0]), .Y(n1953) );
  nr2d1_hd U784 ( .A(n1577), .B(n2223), .Y(n1787) );
  nd2bd1_hd U785 ( .AN(a[30]), .B(n2108), .Y(n2155) );
  ivd1_hd U786 ( .A(a_e[9]), .Y(n1698) );
  nr2d1_hd U787 ( .A(sum[27]), .B(n1805), .Y(n1944) );
  ao22d1_hd U788 ( .A(b_m[25]), .B(n1668), .C(b_m[26]), .D(n2092), .Y(n1626)
         );
  ao22d1_hd U789 ( .A(a_m[21]), .B(n2001), .C(a_m[22]), .D(n1999), .Y(n1620)
         );
  ao22d1_hd U790 ( .A(a_m[20]), .B(n2003), .C(a_m[19]), .D(n2005), .Y(n1617)
         );
  nr2d1_hd U791 ( .A(b_m[15]), .B(n2061), .Y(n1607) );
  ao22d1_hd U792 ( .A(a_m[13]), .B(n2017), .C(a_m[12]), .D(n2019), .Y(n1605)
         );
  ao22d1_hd U793 ( .A(b_m[9]), .B(n2073), .C(b_m[10]), .D(n2071), .Y(n1598) );
  ao22d1_hd U794 ( .A(a_m[9]), .B(n2025), .C(a_m[8]), .D(n2027), .Y(n1596) );
  ao211d1_hd U795 ( .A(a_m[1]), .B(n2040), .C(a_m[0]), .D(n2041), .Y(n1583) );
  oa22d1_hd U796 ( .A(a_m[1]), .B(n2040), .C(a_m[2]), .D(n2039), .Y(n1582) );
  oa22d1_hd U797 ( .A(b_m[3]), .B(n2086), .C(n1583), .D(n1582), .Y(n1584) );
  ao21d1_hd U798 ( .A(a_m[2]), .B(n2039), .C(n1584), .Y(n1586) );
  oa22d1_hd U799 ( .A(a_m[4]), .B(n2035), .C(a_m[3]), .D(n2038), .Y(n1585) );
  oa22d1_hd U800 ( .A(n1586), .B(n1585), .C(b_m[4]), .D(n2083), .Y(n1587) );
  ao22d1_hd U801 ( .A(a_m[5]), .B(n2033), .C(n1588), .D(n1587), .Y(n1589) );
  nr2d1_hd U802 ( .A(n1589), .B(b_m[6]), .Y(n1590) );
  nr2d1_hd U803 ( .A(n1591), .B(b_m[7]), .Y(n1594) );
  oa211d1_hd U804 ( .A(a_m[7]), .B(n1594), .C(n1593), .D(n1592), .Y(n1595) );
  ao22d1_hd U805 ( .A(a_m[10]), .B(n2023), .C(n1598), .D(n1597), .Y(n1599) );
  nr2d1_hd U806 ( .A(b_m[11]), .B(n1599), .Y(n1602) );
  oa211d1_hd U807 ( .A(a_m[11]), .B(n1602), .C(n1601), .D(n1600), .Y(n1604) );
  oa22d1_hd U808 ( .A(a_m[13]), .B(n2017), .C(a_m[14]), .D(n2015), .Y(n1603)
         );
  ao21d1_hd U809 ( .A(n1605), .B(n1604), .C(n1603), .Y(n1606) );
  ao211d1_hd U810 ( .A(a_m[14]), .B(n2015), .C(n1607), .D(n1606), .Y(n1609) );
  oa22d1_hd U811 ( .A(a_m[16]), .B(n2011), .C(a_m[15]), .D(n2013), .Y(n1608)
         );
  oa22d1_hd U812 ( .A(n1609), .B(n1608), .C(b_m[16]), .D(n2059), .Y(n1610) );
  ao22d1_hd U813 ( .A(a_m[17]), .B(n2009), .C(n1611), .D(n1610), .Y(n1612) );
  nr2d1_hd U814 ( .A(b_m[18]), .B(n1612), .Y(n1615) );
  oa211d1_hd U815 ( .A(a_m[18]), .B(n1615), .C(n1614), .D(n1613), .Y(n1616) );
  ao22d1_hd U816 ( .A(b_m[20]), .B(n2051), .C(n1617), .D(n1616), .Y(n1618) );
  ao22d1_hd U817 ( .A(b_m[22]), .B(n2047), .C(n1620), .D(n1619), .Y(n1621) );
  oa22d1_hd U818 ( .A(a_m[23]), .B(n1997), .C(a_m[24]), .D(n1995), .Y(n1623)
         );
  ao22d1_hd U819 ( .A(a_m[24]), .B(n1995), .C(a_m[25]), .D(n1629), .Y(n1622)
         );
  ivd1_hd U820 ( .A(a_m[0]), .Y(n2089) );
  ao22d1_hd U821 ( .A(n1568), .B(n2041), .C(n2089), .D(n1569), .Y(C2_Z_0) );
  ao22d1_hd U822 ( .A(n1568), .B(n2040), .C(n2088), .D(n1569), .Y(C2_Z_1) );
  ao22d1_hd U823 ( .A(n1568), .B(n2023), .C(n2071), .D(n1569), .Y(C2_Z_10) );
  ao22d1_hd U824 ( .A(n1568), .B(n2021), .C(n2069), .D(n1569), .Y(C2_Z_11) );
  ao22d1_hd U825 ( .A(n1568), .B(n2019), .C(n2067), .D(n1569), .Y(C2_Z_12) );
  ao22d1_hd U826 ( .A(n1568), .B(n2017), .C(n2065), .D(n1569), .Y(C2_Z_13) );
  ao22d1_hd U827 ( .A(n1568), .B(n2015), .C(n2063), .D(n1569), .Y(C2_Z_14) );
  ao22d1_hd U828 ( .A(n1568), .B(n2013), .C(n2061), .D(n1569), .Y(C2_Z_15) );
  ao22d1_hd U829 ( .A(n1568), .B(n2011), .C(n2059), .D(n1569), .Y(C2_Z_16) );
  ao22d1_hd U830 ( .A(n1568), .B(n2009), .C(n2057), .D(n1569), .Y(C2_Z_17) );
  ao22d1_hd U831 ( .A(n1568), .B(n2007), .C(n2055), .D(n1569), .Y(C2_Z_18) );
  ao22d1_hd U832 ( .A(n1568), .B(n2005), .C(n2053), .D(n1569), .Y(C2_Z_19) );
  ao22d1_hd U833 ( .A(n1568), .B(n2039), .C(n2087), .D(n1569), .Y(C2_Z_2) );
  ao22d1_hd U834 ( .A(n1568), .B(n2003), .C(n2051), .D(n1569), .Y(C2_Z_20) );
  ao22d1_hd U835 ( .A(n1568), .B(n2001), .C(n2049), .D(n1569), .Y(C2_Z_21) );
  ao22d1_hd U836 ( .A(n1568), .B(n1999), .C(n2047), .D(n1569), .Y(C2_Z_22) );
  ao22d1_hd U837 ( .A(n1568), .B(n1997), .C(n2045), .D(n1569), .Y(C2_Z_23) );
  ao22d1_hd U838 ( .A(n1568), .B(n1995), .C(n2043), .D(n1569), .Y(C2_Z_24) );
  ao22d1_hd U839 ( .A(n1568), .B(n1629), .C(n1668), .D(n1569), .Y(C2_Z_25) );
  oa21d1_hd U840 ( .A(n2250), .B(n1791), .C(n2092), .Y(C2_Z_26) );
  ao22d1_hd U841 ( .A(n1568), .B(n2038), .C(n2086), .D(n1569), .Y(C2_Z_3) );
  ao22d1_hd U842 ( .A(n1568), .B(n2035), .C(n2083), .D(n1569), .Y(C2_Z_4) );
  ao22d1_hd U843 ( .A(n1568), .B(n2033), .C(n2081), .D(n1569), .Y(C2_Z_5) );
  ao22d1_hd U844 ( .A(n1568), .B(n2031), .C(n2079), .D(n1569), .Y(C2_Z_6) );
  ao22d1_hd U845 ( .A(n1568), .B(n2029), .C(n2077), .D(n1569), .Y(C2_Z_7) );
  ao22d1_hd U846 ( .A(n1568), .B(n2027), .C(n2075), .D(n1569), .Y(C2_Z_8) );
  ao22d1_hd U847 ( .A(n1568), .B(n2025), .C(n2073), .D(n1569), .Y(C2_Z_9) );
  nr2d1_hd U848 ( .A(n2250), .B(n2092), .Y(n1628) );
  ao22d1_hd U849 ( .A(n1311), .B(n1628), .C(n2250), .D(n1791), .Y(
        DP_OP_43J4_124_6938_n32) );
  ao22d1_hd U850 ( .A(b_m[25]), .B(n1791), .C(n1655), .D(n1629), .Y(n1630) );
  oa21d1_hd U851 ( .A(a_m[25]), .B(n1569), .C(n1630), .Y(
        DP_OP_43J4_124_6938_n33) );
  ao22d1_hd U852 ( .A(b_m[24]), .B(n1791), .C(n1655), .D(n1995), .Y(n1631) );
  oa21d1_hd U853 ( .A(a_m[24]), .B(n1569), .C(n1631), .Y(
        DP_OP_43J4_124_6938_n34) );
  ao22d1_hd U854 ( .A(b_m[23]), .B(n1791), .C(n1655), .D(n1997), .Y(n1632) );
  oa21d1_hd U855 ( .A(a_m[23]), .B(n1569), .C(n1632), .Y(
        DP_OP_43J4_124_6938_n35) );
  ao22d1_hd U856 ( .A(n1568), .B(n2047), .C(n1655), .D(n1999), .Y(n1633) );
  oa21d1_hd U857 ( .A(n1311), .B(n1999), .C(n1633), .Y(DP_OP_43J4_124_6938_n36) );
  ao22d1_hd U858 ( .A(b_m[21]), .B(n1791), .C(n1655), .D(n2001), .Y(n1634) );
  oa21d1_hd U859 ( .A(a_m[21]), .B(n1569), .C(n1634), .Y(
        DP_OP_43J4_124_6938_n37) );
  ao22d1_hd U860 ( .A(n1568), .B(n2051), .C(n1655), .D(n2003), .Y(n1635) );
  oa21d1_hd U861 ( .A(n1311), .B(n2003), .C(n1635), .Y(DP_OP_43J4_124_6938_n38) );
  ao22d1_hd U862 ( .A(n1568), .B(n2053), .C(n1655), .D(n2005), .Y(n1636) );
  oa21d1_hd U863 ( .A(n1311), .B(n2005), .C(n1636), .Y(DP_OP_43J4_124_6938_n39) );
  ao22d1_hd U864 ( .A(b_m[18]), .B(n1791), .C(n1655), .D(n2007), .Y(n1637) );
  oa21d1_hd U865 ( .A(a_m[18]), .B(n1569), .C(n1637), .Y(
        DP_OP_43J4_124_6938_n40) );
  ao22d1_hd U866 ( .A(n1568), .B(n2057), .C(n1655), .D(n2009), .Y(n1638) );
  oa21d1_hd U867 ( .A(n1311), .B(n2009), .C(n1638), .Y(DP_OP_43J4_124_6938_n41) );
  ao22d1_hd U868 ( .A(n1568), .B(n2059), .C(n1655), .D(n2011), .Y(n1639) );
  oa21d1_hd U869 ( .A(n1311), .B(n2011), .C(n1639), .Y(DP_OP_43J4_124_6938_n42) );
  ao22d1_hd U870 ( .A(n1568), .B(n2061), .C(n1655), .D(n2013), .Y(n1640) );
  oa21d1_hd U871 ( .A(n1311), .B(n2013), .C(n1640), .Y(DP_OP_43J4_124_6938_n43) );
  ao22d1_hd U872 ( .A(b_m[14]), .B(n1791), .C(n1655), .D(n2015), .Y(n1641) );
  oa21d1_hd U873 ( .A(a_m[14]), .B(n1569), .C(n1641), .Y(
        DP_OP_43J4_124_6938_n44) );
  ao22d1_hd U874 ( .A(b_m[13]), .B(n1791), .C(n1655), .D(n2017), .Y(n1642) );
  oa21d1_hd U875 ( .A(a_m[13]), .B(n1569), .C(n1642), .Y(
        DP_OP_43J4_124_6938_n45) );
  ao22d1_hd U876 ( .A(n1568), .B(n2067), .C(n1655), .D(n2019), .Y(n1643) );
  oa21d1_hd U877 ( .A(n1311), .B(n2019), .C(n1643), .Y(DP_OP_43J4_124_6938_n46) );
  ao22d1_hd U878 ( .A(b_m[11]), .B(n1791), .C(n1655), .D(n2021), .Y(n1644) );
  oa21d1_hd U879 ( .A(a_m[11]), .B(n1569), .C(n1644), .Y(
        DP_OP_43J4_124_6938_n47) );
  ao22d1_hd U880 ( .A(n1568), .B(n2071), .C(n1655), .D(n2023), .Y(n1645) );
  oa21d1_hd U881 ( .A(n1311), .B(n2023), .C(n1645), .Y(DP_OP_43J4_124_6938_n48) );
  ao22d1_hd U882 ( .A(n1568), .B(n2073), .C(n1655), .D(n2025), .Y(n1646) );
  oa21d1_hd U883 ( .A(n1311), .B(n2025), .C(n1646), .Y(DP_OP_43J4_124_6938_n49) );
  ao22d1_hd U884 ( .A(n1568), .B(n2075), .C(n1655), .D(n2027), .Y(n1647) );
  oa21d1_hd U885 ( .A(n1311), .B(n2027), .C(n1647), .Y(DP_OP_43J4_124_6938_n50) );
  ao22d1_hd U886 ( .A(b_m[7]), .B(n1791), .C(n1655), .D(n2029), .Y(n1648) );
  oa21d1_hd U887 ( .A(a_m[7]), .B(n1569), .C(n1648), .Y(
        DP_OP_43J4_124_6938_n51) );
  ao22d1_hd U888 ( .A(b_m[6]), .B(n1791), .C(n1655), .D(n2031), .Y(n1649) );
  oa21d1_hd U889 ( .A(a_m[6]), .B(n1569), .C(n1649), .Y(
        DP_OP_43J4_124_6938_n52) );
  ao22d1_hd U890 ( .A(n1568), .B(n2081), .C(n1655), .D(n2033), .Y(n1650) );
  oa21d1_hd U891 ( .A(n1311), .B(n2033), .C(n1650), .Y(DP_OP_43J4_124_6938_n53) );
  ao22d1_hd U892 ( .A(n1568), .B(n2083), .C(n1655), .D(n2035), .Y(n1651) );
  oa21d1_hd U893 ( .A(n1311), .B(n2035), .C(n1651), .Y(DP_OP_43J4_124_6938_n54) );
  ao22d1_hd U894 ( .A(n1568), .B(n2086), .C(n1655), .D(n2038), .Y(n1652) );
  oa21d1_hd U895 ( .A(n1311), .B(n2038), .C(n1652), .Y(DP_OP_43J4_124_6938_n55) );
  ao22d1_hd U896 ( .A(b_m[2]), .B(n1791), .C(n1655), .D(n2039), .Y(n1653) );
  oa21d1_hd U897 ( .A(a_m[2]), .B(n1569), .C(n1653), .Y(
        DP_OP_43J4_124_6938_n56) );
  ao22d1_hd U898 ( .A(b_m[1]), .B(n1791), .C(n1655), .D(n2040), .Y(n1654) );
  oa21d1_hd U899 ( .A(a_m[1]), .B(n1569), .C(n1654), .Y(
        DP_OP_43J4_124_6938_n57) );
  ao22d1_hd U900 ( .A(b_m[0]), .B(n1791), .C(n1655), .D(n2041), .Y(n1656) );
  oa21d1_hd U901 ( .A(a_m[0]), .B(n1569), .C(n1656), .Y(
        DP_OP_43J4_124_6938_n58) );
  ao22d1_hd U902 ( .A(n1568), .B(n1657), .C(n1709), .D(n1569), .Y(N338) );
  nr4d1_hd U903 ( .A(a_e[1]), .B(a_e[2]), .C(a_e[3]), .D(a_e[4]), .Y(n1658) );
  nd4d1_hd U904 ( .A(a_e[7]), .B(n1658), .C(n2097), .D(n2116), .Y(n1678) );
  nr4d1_hd U905 ( .A(n1678), .B(n2144), .C(n1698), .D(n2099), .Y(n2094) );
  nr4d1_hd U906 ( .A(b_e[2]), .B(b_e[1]), .C(b_e[3]), .D(b_e[4]), .Y(n1659) );
  nd4d1_hd U907 ( .A(b_e[7]), .B(n1659), .C(n2184), .D(n2164), .Y(n1677) );
  nr4d1_hd U908 ( .A(n2166), .B(n1677), .C(n2211), .D(n1683), .Y(n2160) );
  nd4d1_hd U909 ( .A(n2033), .B(n2035), .C(n2025), .D(n2013), .Y(n1667) );
  nr4d1_hd U910 ( .A(b_m[0]), .B(b_m[1]), .C(b_m[2]), .D(b_m[3]), .Y(n1660) );
  nd4d1_hd U911 ( .A(n1660), .B(n2011), .C(n2031), .D(n2017), .Y(n1666) );
  nr4d1_hd U912 ( .A(b_m[25]), .B(b_m[23]), .C(b_m[22]), .D(b_m[26]), .Y(n1664) );
  nr4d1_hd U913 ( .A(b_m[18]), .B(b_m[11]), .C(b_m[14]), .D(b_m[24]), .Y(n1663) );
  nr4d1_hd U914 ( .A(b_m[8]), .B(b_m[7]), .C(b_m[10]), .D(b_m[12]), .Y(n1662)
         );
  nr4d1_hd U915 ( .A(b_m[17]), .B(b_m[19]), .C(b_m[20]), .D(b_m[21]), .Y(n1661) );
  nd4d1_hd U916 ( .A(n1664), .B(n1663), .C(n1662), .D(n1661), .Y(n1665) );
  nr3d1_hd U917 ( .A(n1667), .B(n1666), .C(n1665), .Y(n1711) );
  nd4d1_hd U918 ( .A(n2057), .B(n2075), .C(n2049), .D(n2043), .Y(n1676) );
  nr4d1_hd U919 ( .A(a_m[18]), .B(a_m[12]), .C(a_m[20]), .D(a_m[26]), .Y(n1669) );
  nd4d1_hd U920 ( .A(n1669), .B(n2045), .C(n2047), .D(n1668), .Y(n1675) );
  nr4d1_hd U921 ( .A(a_m[11]), .B(a_m[6]), .C(a_m[9]), .D(a_m[10]), .Y(n1673)
         );
  nr4d1_hd U922 ( .A(a_m[13]), .B(a_m[14]), .C(a_m[15]), .D(a_m[19]), .Y(n1672) );
  nr4d1_hd U923 ( .A(a_m[16]), .B(a_m[5]), .C(a_m[4]), .D(a_m[7]), .Y(n1671)
         );
  nr4d1_hd U924 ( .A(a_m[0]), .B(a_m[1]), .C(a_m[2]), .D(a_m[3]), .Y(n1670) );
  nd4d1_hd U925 ( .A(n1673), .B(n1672), .C(n1671), .D(n1670), .Y(n1674) );
  nr4d1_hd U926 ( .A(b_e[8]), .B(b_e[0]), .C(b_e[9]), .D(n1677), .Y(n1710) );
  nr2d1_hd U927 ( .A(n1710), .B(n2223), .Y(n1750) );
  ao22d1_hd U928 ( .A(b_e[2]), .B(n2137), .C(b_e[3]), .D(n2128), .Y(n1685) );
  nr2d1_hd U929 ( .A(a_e[1]), .B(n2212), .Y(n1681) );
  ao22d1_hd U930 ( .A(b_e[4]), .B(n2121), .C(b_e[5]), .D(n2116), .Y(n1680) );
  ao211d1_hd U931 ( .A(b_e[0]), .B(n2144), .C(n1681), .D(n1688), .Y(n1682) );
  oa211d1_hd U932 ( .A(a_e[7]), .B(n2168), .C(n1685), .D(n1682), .Y(n1684) );
  nd3bd1_hd U933 ( .AN(n1684), .B(n1697), .C(n1700), .Y(n2233) );
  ao211d1_hd U934 ( .A(b_e[6]), .B(n2097), .C(b_e[5]), .D(n2116), .Y(n1692) );
  ivd1_hd U935 ( .A(b_e[4]), .Y(n2190) );
  ivd1_hd U936 ( .A(b_e[3]), .Y(n2161) );
  ao22d1_hd U937 ( .A(a_e[4]), .B(n2190), .C(a_e[3]), .D(n2161), .Y(n1690) );
  ao211d1_hd U938 ( .A(b_e[1]), .B(n2145), .C(b_e[0]), .D(n2144), .Y(n1687) );
  oa22d1_hd U939 ( .A(b_e[1]), .B(n2145), .C(b_e[2]), .D(n2137), .Y(n1686) );
  oa21d1_hd U940 ( .A(n1687), .B(n1686), .C(n1685), .Y(n1689) );
  ao21d1_hd U941 ( .A(n1690), .B(n1689), .C(n1688), .Y(n1691) );
  ao211d1_hd U942 ( .A(a_e[6]), .B(n2164), .C(n1692), .D(n1691), .Y(n1695) );
  scg6d1_hd U943 ( .A(b_e[7]), .B(n1695), .C(n2101), .Y(n1693) );
  oa211d1_hd U944 ( .A(b_e[7]), .B(n1695), .C(n1694), .D(n1693), .Y(n1696) );
  oa21d1_hd U945 ( .A(n2094), .B(n2242), .C(n1575), .Y(n1) );
  oa21d1_hd U946 ( .A(n2160), .B(n2242), .C(n2158), .Y(n2) );
  nr2d1_hd U947 ( .A(n1733), .B(n1975), .Y(n1703) );
  nr4d1_hd U948 ( .A(z_e[2]), .B(z_e[3]), .C(z_e[4]), .D(z_e[5]), .Y(n1702) );
  ivd1_hd U949 ( .A(z_e[6]), .Y(n1745) );
  nd3d1_hd U950 ( .A(z_e[9]), .B(n1702), .C(n1745), .Y(n1728) );
  ivd1_hd U951 ( .A(z_e[9]), .Y(n1987) );
  ao21d1_hd U952 ( .A(n1703), .B(n1728), .C(n1987), .Y(n1705) );
  nr2d1_hd U953 ( .A(n2256), .B(n2228), .Y(n1806) );
  nr2d1_hd U954 ( .A(n1727), .B(n1985), .Y(n1704) );
  scg16d1_hd U955 ( .A(n1705), .B(n1704), .C(n1964), .Y(n2227) );
  nr2d1_hd U956 ( .A(n2227), .B(n1988), .Y(n1706) );
  nr2d1_hd U957 ( .A(n1806), .B(n1706), .Y(n1970) );
  ivd1_hd U958 ( .A(n2256), .Y(n2229) );
  scg4d1_hd U959 ( .A(n2229), .B(z_m[0]), .C(n1287), .D(round_bit), .E(n1573), 
        .F(sum[2]), .G(sum[3]), .H(n1943), .Y(n266) );
  nr2d1_hd U960 ( .A(n1707), .B(n2243), .Y(n2220) );
  nr2d1_hd U961 ( .A(a_s), .B(n1717), .Y(n1708) );
  oa21d1_hd U962 ( .A(n1715), .B(n1708), .C(n1793), .Y(n1714) );
  nr3d1_hd U963 ( .A(n1710), .B(n1792), .C(n1709), .Y(n1713) );
  oa22d1_hd U964 ( .A(n1712), .B(n1792), .C(n1711), .D(n1793), .Y(n1794) );
  ao211d1_hd U965 ( .A(b_s), .B(n1714), .C(n1713), .D(n1794), .Y(n1732) );
  ao21d1_hd U966 ( .A(n1792), .B(n1793), .C(n2223), .Y(n1734) );
  ao211d1_hd U967 ( .A(n1286), .B(n1719), .C(n1734), .D(n1796), .Y(n2257) );
  ao22d1_hd U968 ( .A(a_s), .B(n1572), .C(n1577), .D(z[31]), .Y(n1731) );
  ivd1_hd U969 ( .A(z_m[4]), .Y(n1916) );
  ivd1_hd U970 ( .A(z_m[3]), .Y(n1924) );
  nd4d1_hd U971 ( .A(n1946), .B(n1916), .C(n1924), .D(n1910), .Y(n1720) );
  nr4d1_hd U972 ( .A(z_m[0]), .B(z_m[19]), .C(z_m[2]), .D(n1720), .Y(n1726) );
  ivd1_hd U973 ( .A(z_m[12]), .Y(n1868) );
  ivd1_hd U974 ( .A(z_m[11]), .Y(n1875) );
  nd4d1_hd U975 ( .A(n1886), .B(n1868), .C(n1875), .D(n1862), .Y(n1724) );
  ivd1_hd U976 ( .A(z_m[8]), .Y(n1892) );
  ivd1_hd U977 ( .A(z_m[7]), .Y(n1899) );
  nd4d1_hd U978 ( .A(n1923), .B(n1892), .C(n1899), .D(n1898), .Y(n1723) );
  nd4d1_hd U979 ( .A(n1965), .B(n1826), .C(n1832), .D(n1850), .Y(n1722) );
  ivd1_hd U980 ( .A(z_m[16]), .Y(n1844) );
  ivd1_hd U981 ( .A(z_m[15]), .Y(n1851) );
  nd4d1_hd U982 ( .A(n1874), .B(n1844), .C(n1851), .D(n1838), .Y(n1721) );
  nr4d1_hd U983 ( .A(n1724), .B(n1723), .C(n1722), .D(n1721), .Y(n1725) );
  oa211d1_hd U984 ( .A(n1729), .B(n1735), .C(n1796), .D(z_s), .Y(n1730) );
  oa211d1_hd U985 ( .A(n1732), .B(n2223), .C(n1731), .D(n1730), .Y(n361) );
  ao21d1_hd U986 ( .A(n1733), .B(n1975), .C(z_e[9]), .Y(n1797) );
  nr2d1_hd U987 ( .A(z_e[1]), .B(z_e[0]), .Y(n1778) );
  ivd1_hd U988 ( .A(z_e[2]), .Y(n1773) );
  nr2d1_hd U989 ( .A(z_e[3]), .B(n1772), .Y(n1764) );
  ivd1_hd U990 ( .A(z_e[4]), .Y(n1760) );
  nr2d1_hd U991 ( .A(z_e[5]), .B(n1759), .Y(n1749) );
  nr2d1_hd U992 ( .A(z_e[7]), .B(n1744), .Y(n1736) );
  ao211d1_hd U993 ( .A(z_e[7]), .B(n1744), .C(n1790), .D(n1736), .Y(n1740) );
  nd3d1_hd U994 ( .A(n2212), .B(n2145), .C(n1786), .Y(n1780) );
  nr2d1_hd U995 ( .A(n1780), .B(n1771), .Y(n1770) );
  nd3d1_hd U996 ( .A(n1770), .B(n2161), .C(n2128), .Y(n1765) );
  nr2d1_hd U997 ( .A(n1765), .B(n1758), .Y(n1757) );
  nd3d1_hd U998 ( .A(n1757), .B(n2184), .C(n2116), .Y(n1752) );
  nr2d1_hd U999 ( .A(n1752), .B(n1743), .Y(n1742) );
  nr2d1_hd U1000 ( .A(n1742), .B(n1738), .Y(n1737) );
  ao211d1_hd U1001 ( .A(n1742), .B(n1738), .C(n1800), .D(n1737), .Y(n1739) );
  ao211d1_hd U1002 ( .A(n1577), .B(z[30]), .C(n1740), .D(n1739), .Y(n1741) );
  ao21d1_hd U1003 ( .A(n1752), .B(n1743), .C(n1742), .Y(n1748) );
  ivd1_hd U1004 ( .A(n1790), .Y(n1775) );
  oa21d1_hd U1005 ( .A(n1749), .B(n1745), .C(n1744), .Y(n1746) );
  ao22d1_hd U1006 ( .A(n1577), .B(z[29]), .C(n1775), .D(n1746), .Y(n1747) );
  oa211d1_hd U1007 ( .A(n1748), .B(n1800), .C(n1789), .D(n1747), .Y(n363) );
  ao21d1_hd U1008 ( .A(z_e[5]), .B(n1759), .C(n1749), .Y(n1756) );
  ao22d1_hd U1009 ( .A(b_e[5]), .B(n1804), .C(a_e[5]), .D(n1787), .Y(n1753) );
  oa22d1_hd U1010 ( .A(n1757), .B(n1753), .C(n1800), .D(n1752), .Y(n1754) );
  ao21d1_hd U1011 ( .A(n1577), .B(z[28]), .C(n1754), .Y(n1755) );
  oa211d1_hd U1012 ( .A(n1756), .B(n1790), .C(n1789), .D(n1755), .Y(n364) );
  ao21d1_hd U1013 ( .A(n1765), .B(n1758), .C(n1757), .Y(n1763) );
  oa21d1_hd U1014 ( .A(n1764), .B(n1760), .C(n1759), .Y(n1761) );
  ao22d1_hd U1015 ( .A(n1577), .B(z[27]), .C(n1775), .D(n1761), .Y(n1762) );
  oa211d1_hd U1016 ( .A(n1763), .B(n1800), .C(n1789), .D(n1762), .Y(n365) );
  ao21d1_hd U1017 ( .A(z_e[3]), .B(n1772), .C(n1764), .Y(n1769) );
  ao22d1_hd U1018 ( .A(b_e[3]), .B(n1804), .C(a_e[3]), .D(n1787), .Y(n1766) );
  oa22d1_hd U1019 ( .A(n1770), .B(n1766), .C(n1800), .D(n1765), .Y(n1767) );
  ao21d1_hd U1020 ( .A(n1577), .B(z[26]), .C(n1767), .Y(n1768) );
  oa211d1_hd U1021 ( .A(n1769), .B(n1790), .C(n1789), .D(n1768), .Y(n366) );
  ao21d1_hd U1022 ( .A(n1780), .B(n1771), .C(n1770), .Y(n1777) );
  oa21d1_hd U1023 ( .A(n1778), .B(n1773), .C(n1772), .Y(n1774) );
  ao22d1_hd U1024 ( .A(n1577), .B(z[25]), .C(n1775), .D(n1774), .Y(n1776) );
  oa211d1_hd U1025 ( .A(n1777), .B(n1800), .C(n1789), .D(n1776), .Y(n367) );
  ao21d1_hd U1026 ( .A(z_e[0]), .B(z_e[1]), .C(n1778), .Y(n1785) );
  nr3d1_hd U1027 ( .A(n2212), .B(n1786), .C(n1779), .Y(n1783) );
  nd2bd1_hd U1028 ( .AN(n1786), .B(a_e[1]), .Y(n1781) );
  ao21d1_hd U1029 ( .A(n1781), .B(n1780), .C(n1800), .Y(n1782) );
  ao211d1_hd U1030 ( .A(n1577), .B(z[24]), .C(n1783), .D(n1782), .Y(n1784) );
  oa211d1_hd U1031 ( .A(n1785), .B(n1790), .C(n1789), .D(n1784), .Y(n368) );
  ao22d1_hd U1032 ( .A(n1577), .B(z[23]), .C(n1787), .D(n1786), .Y(n1788) );
  oa211d1_hd U1033 ( .A(z_e[0]), .B(n1790), .C(n1789), .D(n1788), .Y(n369) );
  nr3d1_hd U1034 ( .A(n1793), .B(n1792), .C(n1791), .Y(n1795) );
  nr2d1_hd U1035 ( .A(n1795), .B(n1794), .Y(n1801) );
  ao22d1_hd U1036 ( .A(b_m[25]), .B(n1804), .C(z_m[22]), .D(n1803), .Y(n1799)
         );
  ao22d1_hd U1037 ( .A(a_m[25]), .B(n1572), .C(n1577), .D(z[22]), .Y(n1798) );
  oa211d1_hd U1038 ( .A(n1801), .B(n1800), .C(n1799), .D(n1798), .Y(n370) );
  scg4d1_hd U1039 ( .A(b_m[24]), .B(n1804), .C(z_m[21]), .D(n1803), .E(a_m[24]), .F(n1572), .G(n1577), .H(z[21]), .Y(n371) );
  scg4d1_hd U1040 ( .A(b_m[23]), .B(n1804), .C(z_m[20]), .D(n1803), .E(a_m[23]), .F(n1572), .G(n1577), .H(z[20]), .Y(n372) );
  scg4d1_hd U1041 ( .A(b_m[22]), .B(n1804), .C(z_m[19]), .D(n1803), .E(a_m[22]), .F(n1572), .G(n1577), .H(z[19]), .Y(n373) );
  scg4d1_hd U1042 ( .A(b_m[21]), .B(n1804), .C(z_m[18]), .D(n1803), .E(a_m[21]), .F(n1572), .G(n1577), .H(z[18]), .Y(n374) );
  scg4d1_hd U1043 ( .A(b_m[20]), .B(n1804), .C(z_m[17]), .D(n1803), .E(a_m[20]), .F(n1572), .G(n1577), .H(z[17]), .Y(n375) );
  scg4d1_hd U1044 ( .A(b_m[19]), .B(n1804), .C(z_m[16]), .D(n1803), .E(a_m[19]), .F(n1572), .G(n1577), .H(z[16]), .Y(n376) );
  scg4d1_hd U1045 ( .A(b_m[18]), .B(n1804), .C(z_m[15]), .D(n1803), .E(a_m[18]), .F(n1572), .G(n1577), .H(z[15]), .Y(n377) );
  scg4d1_hd U1046 ( .A(b_m[17]), .B(n1804), .C(z_m[14]), .D(n1803), .E(a_m[17]), .F(n1572), .G(n1577), .H(z[14]), .Y(n378) );
  scg4d1_hd U1047 ( .A(b_m[16]), .B(n1804), .C(z_m[13]), .D(n1803), .E(a_m[16]), .F(n1572), .G(n1577), .H(z[13]), .Y(n379) );
  scg4d1_hd U1048 ( .A(b_m[15]), .B(n1804), .C(z_m[12]), .D(n1803), .E(a_m[15]), .F(n1572), .G(n1577), .H(z[12]), .Y(n380) );
  scg4d1_hd U1049 ( .A(b_m[14]), .B(n1804), .C(z_m[11]), .D(n1803), .E(a_m[14]), .F(n1802), .G(n1577), .H(z[11]), .Y(n381) );
  scg4d1_hd U1050 ( .A(b_m[13]), .B(n1804), .C(z_m[10]), .D(n1803), .E(a_m[13]), .F(n1802), .G(n1577), .H(z[10]), .Y(n382) );
  scg4d1_hd U1051 ( .A(b_m[12]), .B(n1804), .C(z_m[9]), .D(n1803), .E(a_m[12]), 
        .F(n1802), .G(n1577), .H(z[9]), .Y(n383) );
  scg4d1_hd U1052 ( .A(b_m[11]), .B(n1804), .C(z_m[8]), .D(n1803), .E(a_m[11]), 
        .F(n1802), .G(n1577), .H(z[8]), .Y(n384) );
  scg4d1_hd U1053 ( .A(b_m[10]), .B(n1804), .C(z_m[7]), .D(n1803), .E(a_m[10]), 
        .F(n1802), .G(n1577), .H(z[7]), .Y(n385) );
  scg4d1_hd U1054 ( .A(b_m[9]), .B(n1804), .C(z_m[6]), .D(n1803), .E(a_m[9]), 
        .F(n1802), .G(n1577), .H(z[6]), .Y(n386) );
  scg4d1_hd U1055 ( .A(b_m[8]), .B(n1804), .C(z_m[5]), .D(n1803), .E(a_m[8]), 
        .F(n1572), .G(n1577), .H(z[5]), .Y(n387) );
  scg4d1_hd U1056 ( .A(b_m[7]), .B(n1804), .C(z_m[4]), .D(n1803), .E(a_m[7]), 
        .F(n1572), .G(n2257), .H(z[4]), .Y(n388) );
  scg4d1_hd U1057 ( .A(b_m[6]), .B(n1804), .C(z_m[3]), .D(n1803), .E(a_m[6]), 
        .F(n1572), .G(n1577), .H(z[3]), .Y(n389) );
  scg4d1_hd U1058 ( .A(b_m[5]), .B(n1804), .C(z_m[2]), .D(n1803), .E(a_m[5]), 
        .F(n1572), .G(n1577), .H(z[2]), .Y(n390) );
  scg4d1_hd U1059 ( .A(b_m[4]), .B(n1804), .C(z_m[1]), .D(n1803), .E(a_m[4]), 
        .F(n1572), .G(n1577), .H(z[1]), .Y(n391) );
  scg4d1_hd U1060 ( .A(b_m[3]), .B(n1804), .C(z_m[0]), .D(n1803), .E(a_m[3]), 
        .F(n1802), .G(n1577), .H(z[0]), .Y(n392) );
  ao22d1_hd U1061 ( .A(n1972), .B(sum[0]), .C(sticky), .D(n1805), .Y(n1808) );
  ao22d1_hd U1062 ( .A(n1806), .B(round_bit), .C(n1943), .D(sum[1]), .Y(n1807)
         );
  ivd1_hd U1063 ( .A(round_bit), .Y(n1811) );
  ao22d1_hd U1064 ( .A(n1573), .B(sum[1]), .C(n1943), .D(sum[2]), .Y(n1810) );
  nd3d1_hd U1065 ( .A(n2229), .B(guard), .C(n265), .Y(n1809) );
  oa211d1_hd U1066 ( .A(n1811), .B(n265), .C(n1810), .D(n1809), .Y(n394) );
  nr3d1_hd U1067 ( .A(z_m[0]), .B(sticky), .C(round_bit), .Y(n1812) );
  ao22d1_hd U1068 ( .A(n1573), .B(sum[25]), .C(n1943), .D(sum[26]), .Y(n1816)
         );
  nd3d1_hd U1069 ( .A(z_m[0]), .B(z_m[2]), .C(z_m[1]), .Y(n1917) );
  ivd1_hd U1070 ( .A(n1917), .Y(n1918) );
  nd3d1_hd U1071 ( .A(n1918), .B(z_m[4]), .C(z_m[3]), .Y(n1905) );
  nr3d1_hd U1072 ( .A(n1905), .B(n1910), .C(n1923), .Y(n1893) );
  nd3d1_hd U1073 ( .A(n1893), .B(z_m[8]), .C(z_m[7]), .Y(n1881) );
  nr3d1_hd U1074 ( .A(n1881), .B(n1898), .C(n1886), .Y(n1869) );
  nd3d1_hd U1075 ( .A(n1869), .B(z_m[12]), .C(z_m[11]), .Y(n1857) );
  nr3d1_hd U1076 ( .A(n1857), .B(n1862), .C(n1874), .Y(n1845) );
  nd3d1_hd U1077 ( .A(n1845), .B(z_m[16]), .C(z_m[15]), .Y(n1833) );
  nr3d1_hd U1078 ( .A(n1833), .B(n1838), .C(n1850), .Y(n1967) );
  oa21d1_hd U1079 ( .A(n1967), .B(n2258), .C(n1952), .Y(n1829) );
  ao21d1_hd U1080 ( .A(n1971), .B(n1813), .C(n1829), .Y(n1817) );
  oa21d1_hd U1081 ( .A(z_m[21]), .B(n1931), .C(n1817), .Y(n1954) );
  ivd1_hd U1082 ( .A(z_m[19]), .Y(n1962) );
  nr2d1_hd U1083 ( .A(n1962), .B(n1827), .Y(n1823) );
  oa21d1_hd U1084 ( .A(z_m[22]), .B(n1958), .C(n1956), .Y(n1814) );
  ao22d1_hd U1085 ( .A(z_m[22]), .B(n1954), .C(z_m[21]), .D(n1814), .Y(n1815)
         );
  oa211d1_hd U1086 ( .A(n1964), .B(n1945), .C(n1816), .D(n1815), .Y(n395) );
  ao22d1_hd U1087 ( .A(n1573), .B(sum[24]), .C(sum[25]), .D(n1943), .Y(n1820)
         );
  ao22d1_hd U1088 ( .A(z_m[21]), .B(n1817), .C(n1958), .D(n1826), .Y(n1818) );
  ao21d1_hd U1089 ( .A(z_m[20]), .B(n1949), .C(n1818), .Y(n1819) );
  oa211d1_hd U1090 ( .A(n1965), .B(n1945), .C(n1820), .D(n1819), .Y(n396) );
  ao22d1_hd U1091 ( .A(n1573), .B(sum[23]), .C(n1943), .D(sum[24]), .Y(n1825)
         );
  ao21d1_hd U1092 ( .A(n1955), .B(n1962), .C(n1829), .Y(n1821) );
  oa22d1_hd U1093 ( .A(n1821), .B(n1832), .C(n1962), .D(n1956), .Y(n1822) );
  ao21d1_hd U1094 ( .A(n1823), .B(n1832), .C(n1822), .Y(n1824) );
  oa211d1_hd U1095 ( .A(n1826), .B(n1945), .C(n1825), .D(n1824), .Y(n397) );
  ao22d1_hd U1096 ( .A(n1573), .B(sum[22]), .C(n1943), .D(sum[23]), .Y(n1831)
         );
  oa22d1_hd U1097 ( .A(z_m[19]), .B(n1827), .C(n1956), .D(n1838), .Y(n1828) );
  ao21d1_hd U1098 ( .A(z_m[19]), .B(n1829), .C(n1828), .Y(n1830) );
  oa211d1_hd U1099 ( .A(n1832), .B(n1945), .C(n1831), .D(n1830), .Y(n398) );
  nr2d1_hd U1100 ( .A(n1931), .B(n1833), .Y(n1841) );
  ao21d1_hd U1101 ( .A(n1841), .B(n1838), .C(n1949), .Y(n1837) );
  ao22d1_hd U1102 ( .A(n1573), .B(sum[21]), .C(n1943), .D(sum[22]), .Y(n1836)
         );
  ao21d1_hd U1103 ( .A(n1971), .B(n1833), .C(n1932), .Y(n1839) );
  oa21d1_hd U1104 ( .A(z_m[17]), .B(n1931), .C(n1839), .Y(n1834) );
  ao22d1_hd U1105 ( .A(z_m[19]), .B(n1938), .C(z_m[18]), .D(n1834), .Y(n1835)
         );
  oa211d1_hd U1106 ( .A(n1837), .B(n1850), .C(n1836), .D(n1835), .Y(n399) );
  ao22d1_hd U1107 ( .A(n1573), .B(sum[20]), .C(n1943), .D(sum[21]), .Y(n1843)
         );
  oa22d1_hd U1108 ( .A(n1839), .B(n1850), .C(n1838), .D(n1945), .Y(n1840) );
  ao21d1_hd U1109 ( .A(n1841), .B(n1850), .C(n1840), .Y(n1842) );
  oa211d1_hd U1110 ( .A(n1844), .B(n1956), .C(n1843), .D(n1842), .Y(n400) );
  ao22d1_hd U1111 ( .A(n1573), .B(sum[19]), .C(n1943), .D(sum[20]), .Y(n1849)
         );
  scg20d1_hd U1112 ( .A(n2258), .B(n1845), .C(n1932), .Y(n1853) );
  oa21d1_hd U1113 ( .A(z_m[15]), .B(n1931), .C(n1853), .Y(n1847) );
  oa21d1_hd U1114 ( .A(z_m[16]), .B(n1852), .C(n1956), .Y(n1846) );
  ao22d1_hd U1115 ( .A(z_m[16]), .B(n1847), .C(z_m[15]), .D(n1846), .Y(n1848)
         );
  oa211d1_hd U1116 ( .A(n1850), .B(n1945), .C(n1849), .D(n1848), .Y(n401) );
  ao22d1_hd U1117 ( .A(n1573), .B(sum[18]), .C(n1943), .D(sum[19]), .Y(n1856)
         );
  ao22d1_hd U1118 ( .A(z_m[15]), .B(n1853), .C(n1852), .D(n1851), .Y(n1854) );
  ao21d1_hd U1119 ( .A(z_m[16]), .B(n1938), .C(n1854), .Y(n1855) );
  oa211d1_hd U1120 ( .A(n1862), .B(n1956), .C(n1856), .D(n1855), .Y(n402) );
  nr2d1_hd U1121 ( .A(n1931), .B(n1857), .Y(n1865) );
  ao21d1_hd U1122 ( .A(n1865), .B(n1862), .C(n1949), .Y(n1861) );
  ao22d1_hd U1123 ( .A(n1573), .B(sum[17]), .C(n1943), .D(sum[18]), .Y(n1860)
         );
  ao21d1_hd U1124 ( .A(n1971), .B(n1857), .C(n1932), .Y(n1863) );
  oa21d1_hd U1125 ( .A(z_m[13]), .B(n1931), .C(n1863), .Y(n1858) );
  ao22d1_hd U1126 ( .A(z_m[14]), .B(n1858), .C(z_m[15]), .D(n1938), .Y(n1859)
         );
  oa211d1_hd U1127 ( .A(n1861), .B(n1874), .C(n1860), .D(n1859), .Y(n403) );
  ao22d1_hd U1128 ( .A(n1573), .B(sum[16]), .C(n1943), .D(sum[17]), .Y(n1867)
         );
  oa22d1_hd U1129 ( .A(n1863), .B(n1874), .C(n1862), .D(n1945), .Y(n1864) );
  ao21d1_hd U1130 ( .A(n1865), .B(n1874), .C(n1864), .Y(n1866) );
  oa211d1_hd U1131 ( .A(n1868), .B(n1956), .C(n1867), .D(n1866), .Y(n404) );
  ao22d1_hd U1132 ( .A(n1573), .B(sum[15]), .C(n1943), .D(sum[16]), .Y(n1873)
         );
  scg20d1_hd U1133 ( .A(n2258), .B(n1869), .C(n1932), .Y(n1877) );
  oa21d1_hd U1134 ( .A(z_m[11]), .B(n1931), .C(n1877), .Y(n1871) );
  oa21d1_hd U1135 ( .A(z_m[12]), .B(n1876), .C(n1956), .Y(n1870) );
  ao22d1_hd U1136 ( .A(z_m[12]), .B(n1871), .C(z_m[11]), .D(n1870), .Y(n1872)
         );
  oa211d1_hd U1137 ( .A(n1874), .B(n1945), .C(n1873), .D(n1872), .Y(n405) );
  ao22d1_hd U1138 ( .A(n1573), .B(sum[14]), .C(n1943), .D(sum[15]), .Y(n1880)
         );
  ao22d1_hd U1139 ( .A(z_m[11]), .B(n1877), .C(n1876), .D(n1875), .Y(n1878) );
  ao21d1_hd U1140 ( .A(z_m[12]), .B(n1938), .C(n1878), .Y(n1879) );
  oa211d1_hd U1141 ( .A(n1886), .B(n1956), .C(n1880), .D(n1879), .Y(n406) );
  nr2d1_hd U1142 ( .A(n1931), .B(n1881), .Y(n1889) );
  ao21d1_hd U1143 ( .A(n1889), .B(n1886), .C(n1949), .Y(n1885) );
  ao22d1_hd U1144 ( .A(n1573), .B(sum[13]), .C(n1943), .D(sum[14]), .Y(n1884)
         );
  ao21d1_hd U1145 ( .A(n1971), .B(n1881), .C(n1932), .Y(n1887) );
  oa21d1_hd U1146 ( .A(z_m[9]), .B(n1931), .C(n1887), .Y(n1882) );
  ao22d1_hd U1147 ( .A(z_m[10]), .B(n1882), .C(z_m[11]), .D(n1938), .Y(n1883)
         );
  oa211d1_hd U1148 ( .A(n1885), .B(n1898), .C(n1884), .D(n1883), .Y(n407) );
  ao22d1_hd U1149 ( .A(n1573), .B(sum[12]), .C(n1943), .D(sum[13]), .Y(n1891)
         );
  oa22d1_hd U1150 ( .A(n1887), .B(n1898), .C(n1886), .D(n1945), .Y(n1888) );
  ao21d1_hd U1151 ( .A(n1889), .B(n1898), .C(n1888), .Y(n1890) );
  oa211d1_hd U1152 ( .A(n1892), .B(n1956), .C(n1891), .D(n1890), .Y(n408) );
  ao22d1_hd U1153 ( .A(n1573), .B(sum[11]), .C(n1943), .D(sum[12]), .Y(n1897)
         );
  scg20d1_hd U1154 ( .A(n2258), .B(n1893), .C(n1932), .Y(n1901) );
  oa21d1_hd U1155 ( .A(z_m[7]), .B(n1931), .C(n1901), .Y(n1895) );
  oa21d1_hd U1156 ( .A(z_m[8]), .B(n1900), .C(n1956), .Y(n1894) );
  ao22d1_hd U1157 ( .A(z_m[8]), .B(n1895), .C(z_m[7]), .D(n1894), .Y(n1896) );
  oa211d1_hd U1158 ( .A(n1898), .B(n1945), .C(n1897), .D(n1896), .Y(n409) );
  ao22d1_hd U1159 ( .A(n1573), .B(sum[10]), .C(n1943), .D(sum[11]), .Y(n1904)
         );
  ao22d1_hd U1160 ( .A(z_m[7]), .B(n1901), .C(n1900), .D(n1899), .Y(n1902) );
  ao21d1_hd U1161 ( .A(z_m[8]), .B(n1938), .C(n1902), .Y(n1903) );
  oa211d1_hd U1162 ( .A(n1910), .B(n1956), .C(n1904), .D(n1903), .Y(n410) );
  nr2d1_hd U1163 ( .A(n1931), .B(n1905), .Y(n1913) );
  ao21d1_hd U1164 ( .A(n1913), .B(n1910), .C(n1949), .Y(n1909) );
  ao22d1_hd U1165 ( .A(n1573), .B(sum[9]), .C(n1943), .D(sum[10]), .Y(n1908)
         );
  ao21d1_hd U1166 ( .A(n1971), .B(n1905), .C(n1932), .Y(n1911) );
  oa21d1_hd U1167 ( .A(z_m[5]), .B(n1931), .C(n1911), .Y(n1906) );
  ao22d1_hd U1168 ( .A(z_m[6]), .B(n1906), .C(z_m[7]), .D(n1938), .Y(n1907) );
  oa211d1_hd U1169 ( .A(n1909), .B(n1923), .C(n1908), .D(n1907), .Y(n411) );
  ao22d1_hd U1170 ( .A(n1573), .B(sum[8]), .C(n1943), .D(sum[9]), .Y(n1915) );
  oa22d1_hd U1171 ( .A(n1911), .B(n1923), .C(n1910), .D(n1945), .Y(n1912) );
  ao21d1_hd U1172 ( .A(n1913), .B(n1923), .C(n1912), .Y(n1914) );
  oa211d1_hd U1173 ( .A(n1916), .B(n1956), .C(n1915), .D(n1914), .Y(n412) );
  ao22d1_hd U1174 ( .A(n1573), .B(sum[7]), .C(n1943), .D(sum[8]), .Y(n1922) );
  ao21d1_hd U1175 ( .A(n1971), .B(n1917), .C(n1932), .Y(n1926) );
  oa21d1_hd U1176 ( .A(z_m[3]), .B(n1931), .C(n1926), .Y(n1920) );
  oa21d1_hd U1177 ( .A(z_m[4]), .B(n1925), .C(n1956), .Y(n1919) );
  ao22d1_hd U1178 ( .A(z_m[4]), .B(n1920), .C(z_m[3]), .D(n1919), .Y(n1921) );
  oa211d1_hd U1179 ( .A(n1923), .B(n1945), .C(n1922), .D(n1921), .Y(n413) );
  ao22d1_hd U1180 ( .A(n1573), .B(sum[6]), .C(n1943), .D(sum[7]), .Y(n1929) );
  ao22d1_hd U1181 ( .A(z_m[3]), .B(n1926), .C(n1925), .D(n1924), .Y(n1927) );
  ao21d1_hd U1182 ( .A(z_m[4]), .B(n1938), .C(n1927), .Y(n1928) );
  scg15d1_hd U1183 ( .A(z_m[2]), .B(n1949), .C(n1929), .D(n1928), .Y(n414) );
  nr3d1_hd U1184 ( .A(z_m[2]), .B(n1931), .C(n1953), .Y(n1930) );
  nr2d1_hd U1185 ( .A(n1930), .B(n1949), .Y(n1936) );
  ao22d1_hd U1186 ( .A(n1573), .B(sum[5]), .C(n1943), .D(sum[6]), .Y(n1935) );
  nr2d1_hd U1187 ( .A(z_m[0]), .B(n1931), .Y(n1948) );
  nr2d1_hd U1188 ( .A(n1932), .B(n1948), .Y(n1942) );
  ao22d1_hd U1189 ( .A(z_m[2]), .B(n1933), .C(z_m[3]), .D(n1938), .Y(n1934) );
  oa211d1_hd U1190 ( .A(n1936), .B(n1946), .C(n1935), .D(n1934), .Y(n415) );
  ao22d1_hd U1191 ( .A(n1573), .B(sum[4]), .C(n1943), .D(sum[5]), .Y(n1941) );
  ao22d1_hd U1192 ( .A(z_m[0]), .B(n1939), .C(z_m[2]), .D(n1938), .Y(n1940) );
  oa211d1_hd U1193 ( .A(n1942), .B(n1946), .C(n1941), .D(n1940), .Y(n416) );
  ao22d1_hd U1194 ( .A(n1573), .B(sum[3]), .C(n1943), .D(sum[4]), .Y(n1951) );
  nr2d1_hd U1195 ( .A(n1946), .B(n1945), .Y(n1947) );
  ao211d1_hd U1196 ( .A(n1949), .B(guard), .C(n1948), .D(n1947), .Y(n1950) );
  oa211d1_hd U1197 ( .A(n1953), .B(n1952), .C(n1951), .D(n1950), .Y(n417) );
  ao21d1_hd U1198 ( .A(n1955), .B(n1965), .C(n1954), .Y(n1961) );
  oa21d1_hd U1199 ( .A(n1958), .B(n1957), .C(n1956), .Y(n1959) );
  ao22d1_hd U1200 ( .A(z_m[22]), .B(n1959), .C(n1972), .D(sum[26]), .Y(n1960)
         );
  oa211d1_hd U1201 ( .A(n1961), .B(n1964), .C(n1960), .D(n1969), .Y(n418) );
  nr4d1_hd U1202 ( .A(n1965), .B(n1964), .C(n1963), .D(n1962), .Y(n1966) );
  nd4d1_hd U1203 ( .A(z_m[21]), .B(z_m[20]), .C(n1967), .D(n1966), .Y(n1968)
         );
  nd4d1_hd U1204 ( .A(n1970), .B(n1282), .C(n1969), .D(n1968), .Y(n1984) );
  nr3d1_hd U1205 ( .A(n1972), .B(state[1]), .C(n1971), .Y(n1973) );
  ao22d1_hd U1206 ( .A(a_e[8]), .B(n1570), .C(n1990), .D(C91_DATA2_8), .Y(
        n1974) );
  oa21d1_hd U1207 ( .A(n1975), .B(n1984), .C(n1974), .Y(n419) );
  ao22d1_hd U1208 ( .A(z_e[7]), .B(n1986), .C(n1990), .D(C91_DATA2_7), .Y(
        n1976) );
  oa21d1_hd U1209 ( .A(n2101), .B(n1282), .C(n1976), .Y(n420) );
  ao22d1_hd U1210 ( .A(z_e[6]), .B(n1986), .C(n1990), .D(C91_DATA2_6), .Y(
        n1977) );
  oa21d1_hd U1211 ( .A(n2097), .B(n1282), .C(n1977), .Y(n421) );
  ao22d1_hd U1212 ( .A(z_e[5]), .B(n1986), .C(n1990), .D(C91_DATA2_5), .Y(
        n1978) );
  oa21d1_hd U1213 ( .A(n2116), .B(n1282), .C(n1978), .Y(n422) );
  ao22d1_hd U1214 ( .A(z_e[4]), .B(n1986), .C(n1990), .D(C91_DATA2_4), .Y(
        n1979) );
  oa21d1_hd U1215 ( .A(n2121), .B(n1282), .C(n1979), .Y(n423) );
  ao22d1_hd U1216 ( .A(z_e[3]), .B(n1986), .C(n1990), .D(C91_DATA2_3), .Y(
        n1980) );
  oa21d1_hd U1217 ( .A(n2128), .B(n1282), .C(n1980), .Y(n424) );
  ao22d1_hd U1218 ( .A(z_e[2]), .B(n1986), .C(n1990), .D(C91_DATA2_2), .Y(
        n1981) );
  oa21d1_hd U1219 ( .A(n2137), .B(n1282), .C(n1981), .Y(n425) );
  ao22d1_hd U1220 ( .A(z_e[1]), .B(n1986), .C(n1990), .D(C91_DATA2_1), .Y(
        n1982) );
  oa21d1_hd U1221 ( .A(n2145), .B(n1282), .C(n1982), .Y(n426) );
  ao22d1_hd U1222 ( .A(a_e[0]), .B(n1570), .C(n1990), .D(n1985), .Y(n1983) );
  oa21d1_hd U1223 ( .A(n1985), .B(n1984), .C(n1983), .Y(n427) );
  ao22d1_hd U1224 ( .A(a_e[9]), .B(n1570), .C(z_e[9]), .D(n1986), .Y(n1993) );
  ao22d1_hd U1225 ( .A(z_e[9]), .B(n1287), .C(n1988), .D(n1987), .Y(n1991) );
  oa211d1_hd U1226 ( .A(DP_OP_154J4_137_6175_n2), .B(n1991), .C(n1990), .D(
        n1989), .Y(n1992) );
  ao22d1_hd U1227 ( .A(b_m[25]), .B(n2036), .C(n1578), .D(b[21]), .Y(n1994) );
  oa21d1_hd U1228 ( .A(n1995), .B(n1576), .C(n1994), .Y(n429) );
  ao22d1_hd U1229 ( .A(b_m[24]), .B(n2036), .C(n1579), .D(b[20]), .Y(n1996) );
  oa21d1_hd U1230 ( .A(n1997), .B(n1576), .C(n1996), .Y(n430) );
  ao22d1_hd U1231 ( .A(b_m[23]), .B(n2036), .C(n1580), .D(b[19]), .Y(n1998) );
  oa21d1_hd U1232 ( .A(n1999), .B(n1576), .C(n1998), .Y(n431) );
  ao22d1_hd U1233 ( .A(b_m[22]), .B(n2036), .C(n1579), .D(b[18]), .Y(n2000) );
  oa21d1_hd U1234 ( .A(n2001), .B(n1576), .C(n2000), .Y(n432) );
  ao22d1_hd U1235 ( .A(b_m[21]), .B(n2036), .C(n1579), .D(b[17]), .Y(n2002) );
  oa21d1_hd U1236 ( .A(n2003), .B(n1576), .C(n2002), .Y(n433) );
  ao22d1_hd U1237 ( .A(b_m[20]), .B(n2036), .C(n1579), .D(b[16]), .Y(n2004) );
  oa21d1_hd U1238 ( .A(n2005), .B(n1576), .C(n2004), .Y(n434) );
  ao22d1_hd U1239 ( .A(b_m[19]), .B(n2036), .C(n1579), .D(b[15]), .Y(n2006) );
  oa21d1_hd U1240 ( .A(n2007), .B(n1576), .C(n2006), .Y(n435) );
  ao22d1_hd U1241 ( .A(b_m[18]), .B(n2036), .C(n1579), .D(b[14]), .Y(n2008) );
  oa21d1_hd U1242 ( .A(n2009), .B(n1576), .C(n2008), .Y(n436) );
  ao22d1_hd U1243 ( .A(b_m[17]), .B(n2036), .C(n1579), .D(b[13]), .Y(n2010) );
  oa21d1_hd U1244 ( .A(n2011), .B(n1576), .C(n2010), .Y(n437) );
  ao22d1_hd U1245 ( .A(b_m[16]), .B(n2036), .C(n1579), .D(b[12]), .Y(n2012) );
  oa21d1_hd U1246 ( .A(n2013), .B(n1576), .C(n2012), .Y(n438) );
  ao22d1_hd U1247 ( .A(b_m[15]), .B(n2036), .C(n1579), .D(b[11]), .Y(n2014) );
  oa21d1_hd U1248 ( .A(n2015), .B(n1576), .C(n2014), .Y(n439) );
  ao22d1_hd U1249 ( .A(b_m[14]), .B(n2036), .C(n1579), .D(b[10]), .Y(n2016) );
  oa21d1_hd U1250 ( .A(n2017), .B(n1576), .C(n2016), .Y(n440) );
  ao22d1_hd U1251 ( .A(b_m[13]), .B(n2036), .C(n1579), .D(b[9]), .Y(n2018) );
  oa21d1_hd U1252 ( .A(n2019), .B(n1576), .C(n2018), .Y(n441) );
  ao22d1_hd U1253 ( .A(b_m[12]), .B(n2036), .C(n1579), .D(b[8]), .Y(n2020) );
  oa21d1_hd U1254 ( .A(n2021), .B(n1576), .C(n2020), .Y(n442) );
  ao22d1_hd U1255 ( .A(b_m[11]), .B(n2036), .C(n1579), .D(b[7]), .Y(n2022) );
  oa21d1_hd U1256 ( .A(n2023), .B(n1576), .C(n2022), .Y(n443) );
  ao22d1_hd U1257 ( .A(b_m[10]), .B(n2036), .C(n1579), .D(b[6]), .Y(n2024) );
  oa21d1_hd U1258 ( .A(n2025), .B(n1576), .C(n2024), .Y(n444) );
  ao22d1_hd U1259 ( .A(b_m[9]), .B(n2036), .C(n1579), .D(b[5]), .Y(n2026) );
  oa21d1_hd U1260 ( .A(n2027), .B(n1576), .C(n2026), .Y(n445) );
  ao22d1_hd U1261 ( .A(b_m[8]), .B(n2036), .C(n1579), .D(b[4]), .Y(n2028) );
  oa21d1_hd U1262 ( .A(n2029), .B(n1576), .C(n2028), .Y(n446) );
  ao22d1_hd U1263 ( .A(b_m[7]), .B(n2036), .C(n1579), .D(b[3]), .Y(n2030) );
  oa21d1_hd U1264 ( .A(n2031), .B(n1576), .C(n2030), .Y(n447) );
  ao22d1_hd U1265 ( .A(b_m[6]), .B(n2036), .C(n1579), .D(b[2]), .Y(n2032) );
  oa21d1_hd U1266 ( .A(n2033), .B(n1576), .C(n2032), .Y(n448) );
  ao22d1_hd U1267 ( .A(b_m[5]), .B(n2036), .C(n1579), .D(b[1]), .Y(n2034) );
  oa21d1_hd U1268 ( .A(n2035), .B(n1576), .C(n2034), .Y(n449) );
  ao22d1_hd U1269 ( .A(b_m[4]), .B(n2036), .C(n1579), .D(b[0]), .Y(n2037) );
  oa21d1_hd U1270 ( .A(n2038), .B(n1576), .C(n2037), .Y(n450) );
  oa22d1_hd U1271 ( .A(n2039), .B(n1576), .C(n2038), .D(n2249), .Y(n451) );
  oa22d1_hd U1272 ( .A(n2040), .B(n1576), .C(n2039), .D(n2249), .Y(n452) );
  oa22d1_hd U1273 ( .A(n1580), .B(n2041), .C(n2040), .D(n2249), .Y(n453) );
  ao22d1_hd U1274 ( .A(a_m[25]), .B(n2084), .C(n1579), .D(a[21]), .Y(n2042) );
  oa21d1_hd U1275 ( .A(n2043), .B(n1574), .C(n2042), .Y(n454) );
  ao22d1_hd U1276 ( .A(a_m[24]), .B(n2084), .C(n1579), .D(a[20]), .Y(n2044) );
  oa21d1_hd U1277 ( .A(n2045), .B(n1574), .C(n2044), .Y(n455) );
  ao22d1_hd U1278 ( .A(a_m[23]), .B(n2084), .C(n1579), .D(a[19]), .Y(n2046) );
  oa21d1_hd U1279 ( .A(n2047), .B(n1574), .C(n2046), .Y(n456) );
  ao22d1_hd U1280 ( .A(a_m[22]), .B(n2084), .C(n1579), .D(a[18]), .Y(n2048) );
  oa21d1_hd U1281 ( .A(n2049), .B(n1574), .C(n2048), .Y(n457) );
  ao22d1_hd U1282 ( .A(a_m[21]), .B(n2084), .C(n1579), .D(a[17]), .Y(n2050) );
  oa21d1_hd U1283 ( .A(n2051), .B(n1574), .C(n2050), .Y(n458) );
  ao22d1_hd U1284 ( .A(a_m[20]), .B(n2084), .C(n1580), .D(a[16]), .Y(n2052) );
  oa21d1_hd U1285 ( .A(n2053), .B(n1574), .C(n2052), .Y(n459) );
  ao22d1_hd U1286 ( .A(a_m[19]), .B(n2084), .C(n1579), .D(a[15]), .Y(n2054) );
  oa21d1_hd U1287 ( .A(n2055), .B(n1574), .C(n2054), .Y(n460) );
  ao22d1_hd U1288 ( .A(a_m[18]), .B(n2084), .C(n1579), .D(a[14]), .Y(n2056) );
  oa21d1_hd U1289 ( .A(n2057), .B(n1574), .C(n2056), .Y(n461) );
  ao22d1_hd U1290 ( .A(a_m[17]), .B(n2084), .C(n1580), .D(a[13]), .Y(n2058) );
  oa21d1_hd U1291 ( .A(n2059), .B(n1574), .C(n2058), .Y(n462) );
  ao22d1_hd U1292 ( .A(a_m[16]), .B(n2084), .C(n1579), .D(a[12]), .Y(n2060) );
  oa21d1_hd U1293 ( .A(n2061), .B(n1574), .C(n2060), .Y(n463) );
  ao22d1_hd U1294 ( .A(a_m[15]), .B(n2084), .C(n1580), .D(a[11]), .Y(n2062) );
  oa21d1_hd U1295 ( .A(n2063), .B(n1574), .C(n2062), .Y(n464) );
  ao22d1_hd U1296 ( .A(a_m[14]), .B(n2084), .C(n1578), .D(a[10]), .Y(n2064) );
  oa21d1_hd U1297 ( .A(n2065), .B(n1574), .C(n2064), .Y(n465) );
  ao22d1_hd U1298 ( .A(a_m[13]), .B(n2084), .C(n1578), .D(a[9]), .Y(n2066) );
  oa21d1_hd U1299 ( .A(n2067), .B(n1574), .C(n2066), .Y(n466) );
  ao22d1_hd U1300 ( .A(a_m[12]), .B(n2084), .C(n1578), .D(a[8]), .Y(n2068) );
  oa21d1_hd U1301 ( .A(n2069), .B(n1574), .C(n2068), .Y(n467) );
  ao22d1_hd U1302 ( .A(a_m[11]), .B(n2084), .C(n1578), .D(a[7]), .Y(n2070) );
  oa21d1_hd U1303 ( .A(n2071), .B(n1574), .C(n2070), .Y(n468) );
  ao22d1_hd U1304 ( .A(a_m[10]), .B(n2084), .C(n1578), .D(a[6]), .Y(n2072) );
  oa21d1_hd U1305 ( .A(n2073), .B(n1574), .C(n2072), .Y(n469) );
  ao22d1_hd U1306 ( .A(a_m[9]), .B(n2084), .C(n1578), .D(a[5]), .Y(n2074) );
  oa21d1_hd U1307 ( .A(n2075), .B(n1574), .C(n2074), .Y(n470) );
  ao22d1_hd U1308 ( .A(a_m[8]), .B(n2084), .C(n1578), .D(a[4]), .Y(n2076) );
  oa21d1_hd U1309 ( .A(n2077), .B(n1574), .C(n2076), .Y(n471) );
  ao22d1_hd U1310 ( .A(a_m[7]), .B(n2084), .C(n1578), .D(a[3]), .Y(n2078) );
  oa21d1_hd U1311 ( .A(n2079), .B(n1574), .C(n2078), .Y(n472) );
  ao22d1_hd U1312 ( .A(a_m[6]), .B(n2084), .C(n1579), .D(a[2]), .Y(n2080) );
  oa21d1_hd U1313 ( .A(n2081), .B(n1574), .C(n2080), .Y(n473) );
  ao22d1_hd U1314 ( .A(a_m[5]), .B(n2084), .C(n1578), .D(a[1]), .Y(n2082) );
  oa21d1_hd U1315 ( .A(n2083), .B(n1574), .C(n2082), .Y(n474) );
  ao22d1_hd U1316 ( .A(a_m[4]), .B(n2084), .C(n1578), .D(a[0]), .Y(n2085) );
  oa21d1_hd U1317 ( .A(n2086), .B(n1574), .C(n2085), .Y(n475) );
  oa22d1_hd U1318 ( .A(n2087), .B(n1574), .C(n2086), .D(n2091), .Y(n476) );
  oa22d1_hd U1319 ( .A(n2088), .B(n1574), .C(n2087), .D(n2091), .Y(n477) );
  oa22d1_hd U1320 ( .A(n1580), .B(n2089), .C(n2088), .D(n2091), .Y(n478) );
  ao22d1_hd U1321 ( .A(a_m[25]), .B(n1575), .C(n1578), .D(a[22]), .Y(n2090) );
  oa21d1_hd U1322 ( .A(n2092), .B(n2091), .C(n2090), .Y(n479) );
  nr2d1_hd U1323 ( .A(n2145), .B(n2144), .Y(n2133) );
  nr2d1_hd U1324 ( .A(n2128), .B(n2127), .Y(n2118) );
  ao21d1_hd U1325 ( .A(n2186), .B(n2096), .C(n2151), .Y(n2117) );
  oa21d1_hd U1326 ( .A(n2097), .B(n2116), .C(n2186), .Y(n2095) );
  ao21d1_hd U1327 ( .A(n2136), .B(n2101), .C(n2103), .Y(n2153) );
  ivd1_hd U1328 ( .A(a[25]), .Y(n2135) );
  nr2d1_hd U1329 ( .A(n2147), .B(n2135), .Y(n2134) );
  ivd1_hd U1330 ( .A(a[27]), .Y(n2120) );
  nr2d1_hd U1331 ( .A(n2130), .B(n2120), .Y(n2119) );
  ivd1_hd U1332 ( .A(a[29]), .Y(n2106) );
  nr2d1_hd U1333 ( .A(n2113), .B(n2106), .Y(n2100) );
  nr2d1_hd U1334 ( .A(n2100), .B(n1283), .Y(n2108) );
  nr2d1_hd U1335 ( .A(n2154), .B(n2096), .Y(n2112) );
  nr2d1_hd U1336 ( .A(n2097), .B(n2111), .Y(n2102) );
  nd3d1_hd U1337 ( .A(a_e[7]), .B(n2102), .C(n2099), .Y(n2098) );
  oa211d1_hd U1338 ( .A(n2153), .B(n2099), .C(n2155), .D(n2098), .Y(n480) );
  ao22d1_hd U1339 ( .A(a_e[7]), .B(n2103), .C(n2102), .D(n2101), .Y(n2104) );
  oa211d1_hd U1340 ( .A(n1283), .B(n2105), .C(n2104), .D(n2155), .Y(n481) );
  oa21d1_hd U1341 ( .A(a_e[5]), .B(n2154), .C(n2117), .Y(n2109) );
  ao22d1_hd U1342 ( .A(a_e[6]), .B(n2109), .C(n2108), .D(n2107), .Y(n2110) );
  oa211d1_hd U1343 ( .A(a_e[6]), .B(n2111), .C(n2110), .D(n2140), .Y(n482) );
  ao21d1_hd U1344 ( .A(n2112), .B(n2116), .C(n2156), .Y(n2115) );
  oa211d1_hd U1345 ( .A(n2119), .B(a[28]), .C(n1580), .D(n2113), .Y(n2114) );
  oa211d1_hd U1346 ( .A(n2117), .B(n2116), .C(n2115), .D(n2114), .Y(n483) );
  ao211d1_hd U1347 ( .A(n2130), .B(n2120), .C(n2119), .D(n1283), .Y(n2123) );
  ao21d1_hd U1348 ( .A(n2186), .B(n2127), .C(n2151), .Y(n2129) );
  ao21d1_hd U1349 ( .A(n2129), .B(n2126), .C(n2121), .Y(n2122) );
  nr2d1_hd U1350 ( .A(n2123), .B(n2122), .Y(n2124) );
  oa211d1_hd U1351 ( .A(a_e[4]), .B(n2125), .C(n2124), .D(n2140), .Y(n484) );
  oa22d1_hd U1352 ( .A(n2129), .B(n2128), .C(n2127), .D(n2126), .Y(n2132) );
  oa211d1_hd U1353 ( .A(n2134), .B(a[26]), .C(n1580), .D(n2130), .Y(n2131) );
  scg13d1_hd U1354 ( .A(n2132), .B(n2156), .C(n2131), .Y(n485) );
  ao211d1_hd U1355 ( .A(n2147), .B(n2135), .C(n2134), .D(n1283), .Y(n2139) );
  nr2d1_hd U1356 ( .A(a_e[0]), .B(n2154), .Y(n2150) );
  nr2d1_hd U1357 ( .A(n2151), .B(n2150), .Y(n2146) );
  ao21d1_hd U1358 ( .A(n2146), .B(n2143), .C(n2137), .Y(n2138) );
  nr2d1_hd U1359 ( .A(n2139), .B(n2138), .Y(n2141) );
  oa211d1_hd U1360 ( .A(a_e[2]), .B(n2142), .C(n2141), .D(n2140), .Y(n486) );
  oa22d1_hd U1361 ( .A(n2146), .B(n2145), .C(n2144), .D(n2143), .Y(n2149) );
  oa211d1_hd U1362 ( .A(a[23]), .B(a[24]), .C(n1580), .D(n2147), .Y(n2148) );
  scg13d1_hd U1363 ( .A(n2149), .B(n2156), .C(n2148), .Y(n487) );
  ao21d1_hd U1364 ( .A(n2151), .B(a_e[0]), .C(n2150), .Y(n2152) );
  oa21d1_hd U1365 ( .A(a[23]), .B(n1283), .C(n2152), .Y(n488) );
  oa21d1_hd U1366 ( .A(a_e[8]), .B(n2154), .C(n2153), .Y(n2157) );
  scg17d1_hd U1367 ( .A(a_e[9]), .B(n2157), .C(n2156), .D(n2155), .Y(n489) );
  nr2d1_hd U1368 ( .A(n2212), .B(n2211), .Y(n2201) );
  nr2d1_hd U1369 ( .A(n2161), .B(n2195), .Y(n2191) );
  ao21d1_hd U1370 ( .A(n2162), .B(n2186), .C(n2218), .Y(n2185) );
  oa21d1_hd U1371 ( .A(n2164), .B(n2184), .C(n2186), .Y(n2163) );
  ao21d1_hd U1372 ( .A(n2202), .B(n2168), .C(n2170), .Y(n2251) );
  ivd1_hd U1373 ( .A(b[25]), .Y(n2204) );
  nr2d1_hd U1374 ( .A(n2214), .B(n2204), .Y(n2203) );
  ivd1_hd U1375 ( .A(b[27]), .Y(n2188) );
  nr2d1_hd U1376 ( .A(n2198), .B(n2188), .Y(n2187) );
  ivd1_hd U1377 ( .A(b[29]), .Y(n2174) );
  nr2d1_hd U1378 ( .A(n2181), .B(n2174), .Y(n2167) );
  nr2d1_hd U1379 ( .A(n2167), .B(n1283), .Y(n2177) );
  nr2bd1_hd U1380 ( .AN(n2191), .B(n2194), .Y(n2180) );
  nr2d1_hd U1381 ( .A(n2164), .B(n2179), .Y(n2169) );
  nd3d1_hd U1382 ( .A(b_e[7]), .B(n2169), .C(n2166), .Y(n2165) );
  oa211d1_hd U1383 ( .A(n2251), .B(n2166), .C(n2253), .D(n2165), .Y(n490) );
  ao22d1_hd U1384 ( .A(b_e[7]), .B(n2170), .C(n2169), .D(n2168), .Y(n2171) );
  oa211d1_hd U1385 ( .A(n2173), .B(n2172), .C(n2171), .D(n2253), .Y(n491) );
  oa21d1_hd U1386 ( .A(b_e[5]), .B(n2252), .C(n2185), .Y(n2175) );
  ao22d1_hd U1387 ( .A(n2177), .B(n2176), .C(b_e[6]), .D(n2175), .Y(n2178) );
  oa211d1_hd U1388 ( .A(b_e[6]), .B(n2179), .C(n2178), .D(n2207), .Y(n492) );
  ao21d1_hd U1389 ( .A(n2180), .B(n2184), .C(n2254), .Y(n2183) );
  oa211d1_hd U1390 ( .A(n2187), .B(b[28]), .C(n1580), .D(n2181), .Y(n2182) );
  oa211d1_hd U1391 ( .A(n2185), .B(n2184), .C(n2183), .D(n2182), .Y(n493) );
  scg6d1_hd U1392 ( .A(n2195), .B(n2186), .C(n2218), .Y(n2197) );
  ao211d1_hd U1393 ( .A(n2198), .B(n2188), .C(n2187), .D(n1283), .Y(n2189) );
  ao211d1_hd U1394 ( .A(b_e[4]), .B(n2197), .C(n2254), .D(n2189), .Y(n2193) );
  nd3d1_hd U1395 ( .A(n2202), .B(n2191), .C(n2190), .Y(n2192) );
  oa211d1_hd U1396 ( .A(b_e[3]), .B(n2194), .C(n2193), .D(n2192), .Y(n494) );
  nr3d1_hd U1397 ( .A(b_e[3]), .B(n2252), .C(n2195), .Y(n2196) );
  ao211d1_hd U1398 ( .A(b_e[3]), .B(n2197), .C(n2254), .D(n2196), .Y(n2200) );
  oa211d1_hd U1399 ( .A(n2203), .B(b[26]), .C(n1580), .D(n2198), .Y(n2199) );
  nr2d1_hd U1400 ( .A(b_e[0]), .B(n2252), .Y(n2217) );
  nr2d1_hd U1401 ( .A(n2218), .B(n2217), .Y(n2213) );
  ao211d1_hd U1402 ( .A(n2214), .B(n2204), .C(n2203), .D(n1283), .Y(n2205) );
  ao21d1_hd U1403 ( .A(n2206), .B(b_e[2]), .C(n2205), .Y(n2208) );
  oa211d1_hd U1404 ( .A(b_e[2]), .B(n2209), .C(n2208), .D(n2207), .Y(n496) );
  oa22d1_hd U1405 ( .A(n2213), .B(n2212), .C(n2211), .D(n2210), .Y(n2216) );
  oa211d1_hd U1406 ( .A(b[23]), .B(b[24]), .C(n1580), .D(n2214), .Y(n2215) );
  scg13d1_hd U1407 ( .A(n2216), .B(n2254), .C(n2215), .Y(n497) );
  ao21d1_hd U1408 ( .A(n2218), .B(b_e[0]), .C(n2217), .Y(n2219) );
  oa21d1_hd U1409 ( .A(b[23]), .B(n1283), .C(n2219), .Y(n498) );
  scg21d1_hd U1410 ( .A(n2220), .B(o_AB_ACK), .C(i_RST), .D(n1571), .Y(n499)
         );
  oa211d1_hd U1411 ( .A(state[3]), .B(n2225), .C(n2224), .D(n2223), .Y(n2239)
         );
  nd3d1_hd U1412 ( .A(n1581), .B(o_Z_STB), .C(i_Z_ACK), .Y(n2263) );
  nd4d1_hd U1413 ( .A(N41), .B(n2258), .C(n2263), .D(n1282), .Y(n2226) );
  nr3d1_hd U1414 ( .A(n27), .B(n2239), .C(n2226), .Y(n2231) );
  ao22d1_hd U1415 ( .A(n2229), .B(n2228), .C(n1287), .D(n2227), .Y(n2230) );
  oa211d1_hd U1416 ( .A(n2233), .B(n2232), .C(n2231), .D(n2230), .Y(n2259) );
  ivd1_hd U1417 ( .A(n2259), .Y(n2236) );
  nr2d1_hd U1418 ( .A(n2234), .B(n2244), .Y(n2235) );
  ao22d1_hd U1419 ( .A(state[2]), .B(n2236), .C(N41), .D(n2235), .Y(n2237) );
  oa21d1_hd U1420 ( .A(n2238), .B(n2261), .C(n2237), .Y(n500) );
  nr2d1_hd U1421 ( .A(n1287), .B(n2239), .Y(n2241) );
  oa22d1_hd U1422 ( .A(n2241), .B(n2261), .C(n2240), .D(n2259), .Y(n501) );
  oa211d1_hd U1423 ( .A(n2244), .B(state[0]), .C(n2243), .D(n2242), .Y(n2245)
         );
  ivd1_hd U1424 ( .A(n2245), .Y(n2247) );
  oa22d1_hd U1425 ( .A(n2247), .B(n2261), .C(n2246), .D(n2259), .Y(n502) );
  ao22d1_hd U1426 ( .A(b_m[25]), .B(n2158), .C(n1578), .D(b[22]), .Y(n2248) );
  oa21d1_hd U1427 ( .A(n2250), .B(n2249), .C(n2248), .Y(n503) );
  oa21d1_hd U1428 ( .A(b_e[8]), .B(n2252), .C(n2251), .Y(n2255) );
  scg17d1_hd U1429 ( .A(b_e[9]), .B(n2255), .C(n2254), .D(n2253), .Y(n504) );
  oa22d1_hd U1430 ( .A(n2262), .B(n2261), .C(n2260), .D(n2259), .Y(n505) );
  ivd1_hd U1431 ( .A(n2263), .Y(n2264) );
  scg21d1_hd U1432 ( .A(n1581), .B(o_Z_STB), .C(i_RST), .D(n2264), .Y(n506) );
endmodule


module float_multiplier_1 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, 
        i_Z_ACK, i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N34, b_s, round_bit, sticky, z_s, N176, N177, N178, N179, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, C82_DATA2_1, C82_DATA2_2, C82_DATA2_3,
         C82_DATA2_4, C82_DATA2_5, C82_DATA2_6, C81_DATA2_1, C81_DATA2_2,
         C81_DATA2_3, C81_DATA2_4, C81_DATA2_5, C81_DATA2_6, net922, n10, n14,
         n104, n105, n110, n138, n141, n148, n151, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, DP_OP_116J3_127_7148_n3,
         DP_OP_116J3_127_7148_n4, DP_OP_116J3_127_7148_n5,
         DP_OP_116J3_127_7148_n6, DP_OP_116J3_127_7148_n7,
         DP_OP_116J3_127_7148_n8, DP_OP_113J3_124_6892_n3,
         DP_OP_113J3_124_6892_n4, DP_OP_113J3_124_6892_n5,
         DP_OP_113J3_124_6892_n6, DP_OP_113J3_124_6892_n7,
         DP_OP_113J3_124_6892_n8, C1_Z_6, C1_Z_5, C1_Z_4, C1_Z_3, C1_Z_2,
         C1_Z_1, DP_OP_125J3_130_6300_n42, DP_OP_125J3_130_6300_n41,
         DP_OP_125J3_130_6300_n40, DP_OP_125J3_130_6300_n39,
         DP_OP_125J3_130_6300_n38, DP_OP_125J3_130_6300_n37,
         DP_OP_125J3_130_6300_n36, DP_OP_125J3_130_6300_n35,
         DP_OP_125J3_130_6300_n34, DP_OP_125J3_130_6300_n32,
         DP_OP_125J3_130_6300_n31, DP_OP_125J3_130_6300_n30,
         DP_OP_125J3_130_6300_n29, DP_OP_125J3_130_6300_n28,
         DP_OP_125J3_130_6300_n27, DP_OP_125J3_130_6300_n26,
         DP_OP_125J3_130_6300_n25, DP_OP_125J3_130_6300_n20,
         DP_OP_125J3_130_6300_n19, DP_OP_125J3_130_6300_n18,
         DP_OP_125J3_130_6300_n17, DP_OP_125J3_130_6300_n16,
         DP_OP_125J3_130_6300_n15, DP_OP_125J3_130_6300_n14,
         DP_OP_125J3_130_6300_n13, DP_OP_125J3_130_6300_n12,
         DP_OP_125J3_130_6300_n9, DP_OP_125J3_130_6300_n8,
         DP_OP_125J3_130_6300_n7, DP_OP_125J3_130_6300_n6,
         DP_OP_125J3_130_6300_n5, DP_OP_125J3_130_6300_n4,
         DP_OP_125J3_130_6300_n3, DP_OP_125J3_130_6300_n2, n768, n769, n770,
         n771, n772, n773, n774, n775, n1220, n2863, n2865, intadd_3_CI,
         intadd_3_SUM_17_, intadd_3_SUM_16_, intadd_3_SUM_15_,
         intadd_3_SUM_14_, intadd_3_SUM_13_, intadd_3_SUM_12_,
         intadd_3_SUM_11_, intadd_3_SUM_10_, intadd_3_SUM_9_, intadd_3_SUM_8_,
         intadd_3_SUM_7_, intadd_3_SUM_6_, intadd_3_SUM_5_, intadd_3_SUM_4_,
         intadd_3_SUM_3_, intadd_3_SUM_2_, intadd_3_SUM_1_, intadd_3_SUM_0_,
         intadd_3_n18, intadd_3_n17, intadd_3_n16, intadd_3_n15, intadd_3_n14,
         intadd_3_n13, intadd_3_n12, intadd_3_n11, intadd_3_n10, intadd_3_n9,
         intadd_3_n8, intadd_3_n7, intadd_3_n6, intadd_3_n5, intadd_3_n4,
         intadd_3_n3, intadd_3_n2, intadd_3_n1, intadd_6_A_13_, intadd_6_A_11_,
         intadd_6_A_10_, intadd_6_A_9_, intadd_6_A_8_, intadd_6_A_7_,
         intadd_6_A_6_, intadd_6_A_5_, intadd_6_A_4_, intadd_6_A_3_,
         intadd_6_A_2_, intadd_6_A_1_, intadd_6_A_0_, intadd_6_B_13_,
         intadd_6_B_12_, intadd_6_B_11_, intadd_6_B_10_, intadd_6_B_9_,
         intadd_6_B_8_, intadd_6_B_7_, intadd_6_B_6_, intadd_6_B_5_,
         intadd_6_B_4_, intadd_6_B_3_, intadd_6_B_2_, intadd_6_B_1_,
         intadd_6_B_0_, intadd_6_CI, intadd_6_SUM_13_, intadd_6_SUM_12_,
         intadd_6_SUM_11_, intadd_6_SUM_10_, intadd_6_SUM_9_, intadd_6_SUM_8_,
         intadd_6_SUM_7_, intadd_6_SUM_6_, intadd_6_SUM_5_, intadd_6_SUM_4_,
         intadd_6_SUM_3_, intadd_6_SUM_2_, intadd_6_SUM_1_, intadd_6_SUM_0_,
         intadd_6_n14, intadd_6_n13, intadd_6_n12, intadd_6_n11, intadd_6_n10,
         intadd_6_n9, intadd_6_n8, intadd_6_n7, intadd_6_n6, intadd_6_n5,
         intadd_6_n4, intadd_6_n3, intadd_6_n2, intadd_6_n1, intadd_7_A_10_,
         intadd_7_A_8_, intadd_7_A_7_, intadd_7_A_6_, intadd_7_A_5_,
         intadd_7_A_4_, intadd_7_A_3_, intadd_7_A_2_, intadd_7_A_1_,
         intadd_7_A_0_, intadd_7_B_9_, intadd_7_B_2_, intadd_7_B_1_,
         intadd_7_B_0_, intadd_7_CI, intadd_7_SUM_10_, intadd_7_SUM_9_,
         intadd_7_SUM_8_, intadd_7_SUM_7_, intadd_7_SUM_6_, intadd_7_SUM_5_,
         intadd_7_SUM_4_, intadd_7_SUM_3_, intadd_7_SUM_2_, intadd_7_SUM_1_,
         intadd_7_SUM_0_, intadd_7_n11, intadd_7_n10, intadd_7_n9, intadd_7_n8,
         intadd_7_n7, intadd_7_n6, intadd_7_n5, intadd_7_n4, intadd_7_n3,
         intadd_7_n2, intadd_7_n1, intadd_8_A_4_, intadd_8_A_2_, intadd_8_A_1_,
         intadd_8_A_0_, intadd_8_B_8_, intadd_8_B_7_, intadd_8_B_6_,
         intadd_8_B_5_, intadd_8_B_3_, intadd_8_B_2_, intadd_8_B_1_,
         intadd_8_B_0_, intadd_8_CI, intadd_8_n9, intadd_8_n8, intadd_8_n7,
         intadd_8_n6, intadd_8_n5, intadd_8_n4, intadd_8_n3, intadd_8_n2,
         intadd_8_n1, intadd_10_A_5_, intadd_10_A_4_, intadd_10_A_3_,
         intadd_10_A_2_, intadd_10_B_7_, intadd_10_B_6_, intadd_10_B_4_,
         intadd_10_B_3_, intadd_10_B_2_, intadd_10_B_1_, intadd_10_CI,
         intadd_10_SUM_7_, intadd_10_SUM_6_, intadd_10_SUM_5_,
         intadd_10_SUM_4_, intadd_10_SUM_3_, intadd_10_SUM_2_,
         intadd_10_SUM_1_, intadd_10_SUM_0_, intadd_10_n8, intadd_10_n7,
         intadd_10_n6, intadd_10_n5, intadd_10_n4, intadd_10_n3, intadd_10_n2,
         intadd_10_n1, intadd_11_A_4_, intadd_11_A_3_, intadd_11_A_2_,
         intadd_11_A_1_, intadd_11_B_5_, intadd_11_B_3_, intadd_11_B_2_,
         intadd_11_B_1_, intadd_11_B_0_, intadd_11_CI, intadd_11_SUM_5_,
         intadd_11_SUM_4_, intadd_11_SUM_3_, intadd_11_SUM_2_,
         intadd_11_SUM_1_, intadd_11_SUM_0_, intadd_11_n6, intadd_11_n5,
         intadd_11_n4, intadd_11_n3, intadd_11_n2, intadd_11_n1,
         intadd_12_A_1_, intadd_12_B_4_, intadd_12_B_2_, intadd_12_B_1_,
         intadd_12_B_0_, intadd_12_CI, intadd_12_SUM_4_, intadd_12_SUM_3_,
         intadd_12_SUM_2_, intadd_12_SUM_1_, intadd_12_SUM_0_, intadd_12_n5,
         intadd_12_n4, intadd_12_n3, intadd_12_n2, intadd_12_n1,
         intadd_13_A_1_, intadd_13_A_0_, intadd_13_B_2_, intadd_13_B_1_,
         intadd_13_B_0_, intadd_13_CI, intadd_13_SUM_2_, intadd_13_SUM_1_,
         intadd_13_SUM_0_, intadd_13_n3, intadd_13_n2, intadd_13_n1,
         intadd_14_A_1_, intadd_14_B_2_, intadd_14_B_0_, intadd_14_CI,
         intadd_14_SUM_2_, intadd_14_SUM_1_, intadd_14_SUM_0_, intadd_14_n3,
         intadd_14_n2, intadd_14_n1, intadd_15_A_2_, intadd_15_A_1_,
         intadd_15_B_2_, intadd_15_B_1_, intadd_15_B_0_, intadd_15_CI,
         intadd_15_SUM_2_, intadd_15_SUM_1_, intadd_15_SUM_0_, intadd_15_n3,
         intadd_15_n2, intadd_15_n1, intadd_16_A_0_, intadd_16_B_2_,
         intadd_16_B_1_, intadd_16_B_0_, intadd_16_SUM_2_, intadd_16_SUM_1_,
         intadd_16_SUM_0_, intadd_16_n3, intadd_16_n2, intadd_16_n1,
         intadd_17_B_2_, intadd_17_B_1_, intadd_17_B_0_, intadd_17_CI,
         intadd_17_SUM_2_, intadd_17_SUM_1_, intadd_17_SUM_0_, intadd_17_n3,
         intadd_17_n2, intadd_17_n1, intadd_18_B_2_, intadd_18_B_1_,
         intadd_18_B_0_, intadd_18_CI, intadd_18_SUM_2_, intadd_18_n3,
         intadd_18_n2, intadd_18_n1, intadd_19_B_2_, intadd_19_B_1_,
         intadd_19_B_0_, intadd_19_CI, intadd_19_SUM_2_, intadd_19_SUM_1_,
         intadd_19_SUM_0_, intadd_19_n3, intadd_19_n2, intadd_19_n1,
         intadd_20_A_1_, intadd_20_A_0_, intadd_20_B_2_, intadd_20_CI,
         intadd_20_SUM_2_, intadd_20_SUM_1_, intadd_20_SUM_0_, intadd_20_n3,
         intadd_20_n2, intadd_20_n1, intadd_0_A_24_, intadd_0_A_23_,
         intadd_0_A_22_, intadd_0_A_21_, intadd_0_A_20_, intadd_0_A_19_,
         intadd_0_A_18_, intadd_0_A_17_, intadd_0_A_16_, intadd_0_A_15_,
         intadd_0_A_14_, intadd_0_A_13_, intadd_0_A_12_, intadd_0_A_11_,
         intadd_0_A_10_, intadd_0_A_9_, intadd_0_A_8_, intadd_0_A_7_,
         intadd_0_A_6_, intadd_0_A_5_, intadd_0_A_4_, intadd_0_A_3_,
         intadd_0_A_2_, intadd_0_A_1_, intadd_0_A_0_, intadd_0_B_21_,
         intadd_0_B_20_, intadd_0_B_19_, intadd_0_B_18_, intadd_0_B_17_,
         intadd_0_B_16_, intadd_0_B_15_, intadd_0_B_14_, intadd_0_B_13_,
         intadd_0_B_12_, intadd_0_B_11_, intadd_0_B_10_, intadd_0_B_9_,
         intadd_0_B_8_, intadd_0_B_7_, intadd_0_B_6_, intadd_0_B_5_,
         intadd_0_B_4_, intadd_0_B_3_, intadd_0_B_2_, intadd_0_B_1_,
         intadd_0_B_0_, intadd_0_CI, intadd_0_SUM_24_, intadd_0_SUM_23_,
         intadd_0_SUM_22_, intadd_0_SUM_21_, intadd_0_SUM_20_,
         intadd_0_SUM_19_, intadd_0_SUM_18_, intadd_0_SUM_17_,
         intadd_0_SUM_16_, intadd_0_SUM_15_, intadd_0_SUM_14_,
         intadd_0_SUM_13_, intadd_0_SUM_12_, intadd_0_SUM_11_,
         intadd_0_SUM_10_, intadd_0_SUM_9_, intadd_0_SUM_8_, intadd_0_SUM_7_,
         intadd_0_SUM_6_, intadd_0_SUM_5_, intadd_0_SUM_4_, intadd_0_SUM_3_,
         intadd_0_SUM_2_, intadd_0_SUM_1_, intadd_0_SUM_0_, intadd_0_n25,
         intadd_0_n24, intadd_0_n23, intadd_0_n22, intadd_0_n21, intadd_0_n20,
         intadd_0_n19, intadd_0_n18, intadd_0_n17, intadd_0_n16, intadd_0_n15,
         intadd_0_n14, intadd_0_n13, intadd_0_n12, intadd_0_n11, intadd_0_n10,
         intadd_0_n9, intadd_0_n8, intadd_0_n7, intadd_0_n6, intadd_0_n5,
         intadd_0_n4, intadd_0_n3, intadd_0_n2, intadd_0_n1, intadd_1_B_19_,
         intadd_1_B_8_, intadd_1_B_6_, intadd_1_B_5_, intadd_1_B_3_,
         intadd_1_B_2_, intadd_1_B_0_, intadd_1_CI, intadd_1_SUM_8_,
         intadd_1_SUM_7_, intadd_1_SUM_6_, intadd_1_SUM_5_, intadd_1_SUM_4_,
         intadd_1_SUM_3_, intadd_1_SUM_2_, intadd_1_SUM_1_, intadd_1_SUM_0_,
         intadd_1_n20, intadd_1_n19, intadd_1_n18, intadd_1_n17, intadd_1_n16,
         intadd_1_n15, intadd_1_n14, intadd_1_n13, intadd_1_n12, intadd_1_n11,
         intadd_1_n10, intadd_1_n9, intadd_1_n8, intadd_1_n7, intadd_1_n6,
         intadd_1_n5, intadd_1_n4, intadd_1_n3, intadd_1_n2, intadd_1_n1,
         intadd_2_A_18_, intadd_2_A_17_, intadd_2_A_16_, intadd_2_A_15_,
         intadd_2_A_14_, intadd_2_A_13_, intadd_2_A_12_, intadd_2_A_11_,
         intadd_2_A_10_, intadd_2_A_9_, intadd_2_A_8_, intadd_2_A_7_,
         intadd_2_A_6_, intadd_2_A_5_, intadd_2_A_4_, intadd_2_A_3_,
         intadd_2_A_2_, intadd_2_A_1_, intadd_2_A_0_, intadd_2_B_18_,
         intadd_2_B_17_, intadd_2_B_16_, intadd_2_B_15_, intadd_2_B_14_,
         intadd_2_B_13_, intadd_2_B_12_, intadd_2_B_11_, intadd_2_B_10_,
         intadd_2_B_9_, intadd_2_B_8_, intadd_2_B_7_, intadd_2_B_6_,
         intadd_2_B_5_, intadd_2_B_4_, intadd_2_B_3_, intadd_2_B_2_,
         intadd_2_B_1_, intadd_2_B_0_, intadd_2_CI, intadd_2_n19, intadd_2_n18,
         intadd_2_n17, intadd_2_n16, intadd_2_n15, intadd_2_n14, intadd_2_n13,
         intadd_2_n12, intadd_2_n11, intadd_2_n10, intadd_2_n9, intadd_2_n8,
         intadd_2_n7, intadd_2_n6, intadd_2_n5, intadd_2_n4, intadd_2_n3,
         intadd_2_n2, intadd_2_n1, intadd_4_A_16_, intadd_4_A_15_,
         intadd_4_A_14_, intadd_4_A_13_, intadd_4_A_12_, intadd_4_A_11_,
         intadd_4_A_10_, intadd_4_A_9_, intadd_4_A_8_, intadd_4_A_7_,
         intadd_4_A_6_, intadd_4_A_5_, intadd_4_A_4_, intadd_4_A_3_,
         intadd_4_A_2_, intadd_4_A_1_, intadd_4_A_0_, intadd_4_B_16_,
         intadd_4_B_15_, intadd_4_B_14_, intadd_4_B_13_, intadd_4_B_12_,
         intadd_4_B_11_, intadd_4_B_10_, intadd_4_B_9_, intadd_4_B_8_,
         intadd_4_B_7_, intadd_4_B_6_, intadd_4_B_5_, intadd_4_B_4_,
         intadd_4_B_3_, intadd_4_B_2_, intadd_4_B_1_, intadd_4_B_0_,
         intadd_4_CI, intadd_4_n17, intadd_4_n16, intadd_4_n15, intadd_4_n14,
         intadd_4_n13, intadd_4_n12, intadd_4_n11, intadd_4_n10, intadd_4_n9,
         intadd_4_n8, intadd_4_n7, intadd_4_n6, intadd_4_n5, intadd_4_n4,
         intadd_4_n3, intadd_4_n2, intadd_4_n1, intadd_5_A_13_, intadd_5_A_11_,
         intadd_5_A_9_, intadd_5_A_7_, intadd_5_A_6_, intadd_5_A_5_,
         intadd_5_A_4_, intadd_5_A_3_, intadd_5_A_2_, intadd_5_A_1_,
         intadd_5_A_0_, intadd_5_B_16_, intadd_5_B_15_, intadd_5_B_14_,
         intadd_5_B_12_, intadd_5_B_10_, intadd_5_B_8_, intadd_5_B_2_,
         intadd_5_B_1_, intadd_5_B_0_, intadd_5_CI, intadd_5_SUM_16_,
         intadd_5_SUM_15_, intadd_5_SUM_14_, intadd_5_n17, intadd_5_n16,
         intadd_5_n15, intadd_5_n14, intadd_5_n13, intadd_5_n12, intadd_5_n11,
         intadd_5_n10, intadd_5_n9, intadd_5_n8, intadd_5_n7, intadd_5_n6,
         intadd_5_n5, intadd_5_n4, intadd_5_n3, intadd_5_n2, intadd_5_n1,
         intadd_9_B_0_, intadd_9_CI, intadd_9_SUM_0_, intadd_9_n8, intadd_9_n7,
         intadd_9_n6, intadd_9_n5, intadd_9_n4, intadd_9_n3, intadd_9_n2,
         intadd_9_n1, n7, n1103, n1111, n1118, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1133, n1134, n1135,
         n1137, n1138, n1139, n1140, n1142, n1143, n1144, n1146, n1147, n1149,
         n1151, n1152, n1153, n1155, n1156, n1157, n1159, n1160, n1161, n1163,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1208, n1210, n1211, n1221, n1222, n1224, n1225, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1112, n1113, n1114, n1115, n1116, n1117, n1119, n1120, n1132,
         n1136, n1141, n1145, n1148, n1150, n1154, n1158, n1162, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1198, n1207, n1209, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1223, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
  wire   [3:0] state;
  wire   [29:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [23:0] a_m;
  wire   [9:0] b_e;
  wire   [23:1] b_m;
  wire   [49:2] product;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U364 ( .A(i_RST), .Y(N34) );
  fad1_hd DP_OP_116J3_127_7148_U7 ( .A(n1118), .B(n774), .CI(
        DP_OP_116J3_127_7148_n5), .CO(DP_OP_116J3_127_7148_n4), .S(C82_DATA2_5) );
  fad1_hd DP_OP_116J3_127_7148_U8 ( .A(n1118), .B(n773), .CI(
        DP_OP_116J3_127_7148_n6), .CO(DP_OP_116J3_127_7148_n5), .S(C82_DATA2_4) );
  fad1_hd DP_OP_116J3_127_7148_U9 ( .A(n1118), .B(n772), .CI(
        DP_OP_116J3_127_7148_n7), .CO(DP_OP_116J3_127_7148_n6), .S(C82_DATA2_3) );
  fad1_hd DP_OP_116J3_127_7148_U10 ( .A(n1118), .B(n771), .CI(
        DP_OP_116J3_127_7148_n8), .CO(DP_OP_116J3_127_7148_n7), .S(C82_DATA2_2) );
  fad1_hd DP_OP_116J3_127_7148_U11 ( .A(n1118), .B(n770), .CI(n769), .CO(
        DP_OP_116J3_127_7148_n8), .S(C82_DATA2_1) );
  fad1_hd DP_OP_113J3_124_6892_U6 ( .A(n1118), .B(C1_Z_6), .CI(
        DP_OP_113J3_124_6892_n4), .CO(DP_OP_113J3_124_6892_n3), .S(C81_DATA2_6) );
  fad1_hd DP_OP_113J3_124_6892_U7 ( .A(n1118), .B(C1_Z_5), .CI(
        DP_OP_113J3_124_6892_n5), .CO(DP_OP_113J3_124_6892_n4), .S(C81_DATA2_5) );
  fad1_hd DP_OP_113J3_124_6892_U8 ( .A(n1118), .B(C1_Z_4), .CI(
        DP_OP_113J3_124_6892_n6), .CO(DP_OP_113J3_124_6892_n5), .S(C81_DATA2_4) );
  fad1_hd DP_OP_113J3_124_6892_U9 ( .A(n1118), .B(C1_Z_3), .CI(
        DP_OP_113J3_124_6892_n7), .CO(DP_OP_113J3_124_6892_n6), .S(C81_DATA2_3) );
  fad1_hd DP_OP_113J3_124_6892_U10 ( .A(n1118), .B(C1_Z_2), .CI(
        DP_OP_113J3_124_6892_n8), .CO(DP_OP_113J3_124_6892_n7), .S(C81_DATA2_2) );
  fad1_hd DP_OP_113J3_124_6892_U11 ( .A(n1118), .B(C1_Z_1), .CI(n768), .CO(
        DP_OP_113J3_124_6892_n8), .S(C81_DATA2_1) );
  had1_hd DP_OP_125J3_130_6300_U32 ( .A(b_e[0]), .B(a_e[0]), .CO(
        DP_OP_125J3_130_6300_n20), .S(DP_OP_125J3_130_6300_n34) );
  fad1_hd DP_OP_125J3_130_6300_U31 ( .A(a_e[1]), .B(b_e[1]), .CI(
        DP_OP_125J3_130_6300_n20), .CO(DP_OP_125J3_130_6300_n19), .S(
        DP_OP_125J3_130_6300_n35) );
  fad1_hd DP_OP_125J3_130_6300_U30 ( .A(a_e[2]), .B(b_e[2]), .CI(
        DP_OP_125J3_130_6300_n19), .CO(DP_OP_125J3_130_6300_n18), .S(
        DP_OP_125J3_130_6300_n36) );
  fad1_hd DP_OP_125J3_130_6300_U29 ( .A(a_e[3]), .B(b_e[3]), .CI(
        DP_OP_125J3_130_6300_n18), .CO(DP_OP_125J3_130_6300_n17), .S(
        DP_OP_125J3_130_6300_n37) );
  fad1_hd DP_OP_125J3_130_6300_U28 ( .A(a_e[4]), .B(b_e[4]), .CI(
        DP_OP_125J3_130_6300_n17), .CO(DP_OP_125J3_130_6300_n16), .S(
        DP_OP_125J3_130_6300_n38) );
  fad1_hd DP_OP_125J3_130_6300_U27 ( .A(a_e[5]), .B(b_e[5]), .CI(
        DP_OP_125J3_130_6300_n16), .CO(DP_OP_125J3_130_6300_n15), .S(
        DP_OP_125J3_130_6300_n39) );
  fad1_hd DP_OP_125J3_130_6300_U26 ( .A(a_e[6]), .B(b_e[6]), .CI(
        DP_OP_125J3_130_6300_n15), .CO(DP_OP_125J3_130_6300_n14), .S(
        DP_OP_125J3_130_6300_n40) );
  fad1_hd DP_OP_125J3_130_6300_U25 ( .A(a_e[7]), .B(b_e[7]), .CI(
        DP_OP_125J3_130_6300_n14), .CO(DP_OP_125J3_130_6300_n13), .S(
        DP_OP_125J3_130_6300_n41) );
  fad1_hd DP_OP_125J3_130_6300_U24 ( .A(a_e[8]), .B(b_e[8]), .CI(
        DP_OP_125J3_130_6300_n13), .CO(DP_OP_125J3_130_6300_n12), .S(
        DP_OP_125J3_130_6300_n42) );
  fds2d1_hd a_e_reg_7_ ( .CRN(n141), .D(n138), .CK(i_CLK), .Q(n10), .QN(a_e[7]) );
  fds2d1_hd b_e_reg_7_ ( .CRN(n151), .D(n148), .CK(i_CLK), .Q(n14), .QN(b_e[7]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n359), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1021), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1021), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n1021), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n1021), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n1021), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n1021), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1021), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1021), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1021), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1021), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1021), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n1021), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n359), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n359), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n359), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n359), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n359), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n1021), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n1021), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1021), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n1021), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n1021), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n1021), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1021), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1021), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1021), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1021), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1021), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1021), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1021), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1021), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd product_reg_27_ ( .D(n1134), .E(n1004), .CK(i_CLK), .Q(
        product[27]) );
  fd1eqd1_hd product_reg_28_ ( .D(n1133), .E(n1004), .CK(i_CLK), .Q(
        product[28]) );
  fd1eqd1_hd product_reg_30_ ( .D(n1128), .E(n1004), .CK(i_CLK), .Q(
        product[30]) );
  fd1eqd1_hd product_reg_32_ ( .D(N206), .E(n1004), .CK(i_CLK), .Q(product[32]) );
  fd1eqd1_hd product_reg_34_ ( .D(N208), .E(n1004), .CK(i_CLK), .Q(product[34]) );
  fd1eqd1_hd product_reg_36_ ( .D(N210), .E(n1004), .CK(i_CLK), .Q(product[36]) );
  fd1eqd1_hd product_reg_38_ ( .D(N212), .E(n1004), .CK(i_CLK), .Q(product[38]) );
  fd1eqd1_hd product_reg_40_ ( .D(N214), .E(n1004), .CK(i_CLK), .Q(product[40]) );
  fd1eqd1_hd product_reg_42_ ( .D(N216), .E(n1004), .CK(i_CLK), .Q(product[42]) );
  fd1eqd1_hd product_reg_44_ ( .D(N218), .E(n1004), .CK(i_CLK), .Q(product[44]) );
  fd1eqd1_hd product_reg_46_ ( .D(N220), .E(n1004), .CK(i_CLK), .Q(product[46]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n1018), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n1018), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n1018), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd product_reg_24_ ( .D(n1138), .E(n1004), .CK(i_CLK), .Q(
        product[24]) );
  fd1eqd1_hd product_reg_26_ ( .D(n1135), .E(n1004), .CK(i_CLK), .Q(
        product[26]) );
  fd1eqd1_hd product_reg_29_ ( .D(n1131), .E(n1004), .CK(i_CLK), .Q(
        product[29]) );
  fd1eqd1_hd product_reg_31_ ( .D(N205), .E(n1004), .CK(i_CLK), .Q(product[31]) );
  fd1eqd1_hd product_reg_33_ ( .D(N207), .E(n1004), .CK(i_CLK), .Q(product[33]) );
  fd1eqd1_hd product_reg_35_ ( .D(N209), .E(n1004), .CK(i_CLK), .Q(product[35]) );
  fd1eqd1_hd product_reg_37_ ( .D(N211), .E(n1004), .CK(i_CLK), .Q(product[37]) );
  fd1eqd1_hd product_reg_39_ ( .D(N213), .E(n1004), .CK(i_CLK), .Q(product[39]) );
  fd1eqd1_hd product_reg_41_ ( .D(N215), .E(n1004), .CK(i_CLK), .Q(product[41]) );
  fd1eqd1_hd product_reg_43_ ( .D(N217), .E(n1004), .CK(i_CLK), .Q(product[43]) );
  fd1eqd1_hd product_reg_45_ ( .D(N219), .E(n1004), .CK(i_CLK), .Q(product[45]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n1018), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n1018), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n1018), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n1018), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n1018), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n1018), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n1018), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n1018), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n1018), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n1018), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n1018), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n1018), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n1018), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n1018), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n1018), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n1018), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n1018), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n1018), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n1018), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n1018), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n1018), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n1018), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n1018), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n1018), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n1018), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n1018), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n1018), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n1018), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n1018), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n1018), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n1018), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n1018), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n1018), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n1018), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n1018), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n1018), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n1018), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n1018), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n1018), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n1018), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n1018), .CK(i_CLK), .Q(b[22]) );
  fd1eqd1_hd product_reg_47_ ( .D(N221), .E(n1004), .CK(i_CLK), .Q(product[47]) );
  fd1eqd1_hd product_reg_48_ ( .D(N222), .E(n1004), .CK(i_CLK), .Q(product[48]) );
  fd1eqd1_hd product_reg_49_ ( .D(N223), .E(n1004), .CK(i_CLK), .Q(product[49]) );
  fd1eqd1_hd z_s_reg ( .D(b_s), .E(n1004), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd product_reg_25_ ( .D(n1137), .E(n1004), .CK(i_CLK), .Q(
        product[25]) );
  fd1eqd1_hd product_reg_9_ ( .D(n1159), .E(n1004), .CK(i_CLK), .Q(product[9])
         );
  fd1eqd1_hd product_reg_20_ ( .D(n1143), .E(n1004), .CK(i_CLK), .Q(
        product[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n241), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n242), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_17_ ( .D(n243), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n244), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_15_ ( .D(n245), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n246), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_13_ ( .D(n247), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n248), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_11_ ( .D(n249), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n250), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_9_ ( .D(n251), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_3_ ( .D(n257), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_2_ ( .D(n258), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_1_ ( .D(n259), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_0_ ( .D(n260), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_21_ ( .D(n239), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n240), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_29_ ( .D(n231), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n233), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n235), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd product_reg_5_ ( .D(N179), .E(n1004), .CK(i_CLK), .Q(product[5])
         );
  fd1eqd1_hd product_reg_10_ ( .D(n1157), .E(n1004), .CK(i_CLK), .Q(
        product[10]) );
  fd1eqd1_hd product_reg_18_ ( .D(n1146), .E(n1004), .CK(i_CLK), .Q(
        product[18]) );
  fd1eqd1_hd product_reg_19_ ( .D(n1144), .E(n1004), .CK(i_CLK), .Q(
        product[19]) );
  fd1eqd1_hd product_reg_23_ ( .D(n1139), .E(n1004), .CK(i_CLK), .Q(
        product[23]) );
  fd1eqd1_hd product_reg_4_ ( .D(N178), .E(n1004), .CK(i_CLK), .Q(product[4])
         );
  fd1eqd1_hd product_reg_7_ ( .D(n1161), .E(n1004), .CK(i_CLK), .Q(product[7])
         );
  fd1eqd1_hd product_reg_11_ ( .D(n1156), .E(n1004), .CK(i_CLK), .Q(
        product[11]) );
  fd1eqd1_hd product_reg_21_ ( .D(n1142), .E(n1004), .CK(i_CLK), .Q(
        product[21]) );
  fd1eqd1_hd product_reg_22_ ( .D(n1140), .E(n1004), .CK(i_CLK), .Q(
        product[22]) );
  fd1eqd1_hd product_reg_2_ ( .D(N176), .E(n1004), .CK(i_CLK), .Q(product[2])
         );
  fd1eqd1_hd product_reg_6_ ( .D(n1163), .E(n1004), .CK(i_CLK), .Q(product[6])
         );
  fd1eqd1_hd product_reg_15_ ( .D(n1151), .E(n1004), .CK(i_CLK), .Q(
        product[15]) );
  fd1eqd1_hd product_reg_16_ ( .D(n1149), .E(n1004), .CK(i_CLK), .Q(
        product[16]) );
  fd1eqd1_hd product_reg_17_ ( .D(n1147), .E(n1004), .CK(i_CLK), .Q(
        product[17]) );
  fd1eqd1_hd product_reg_3_ ( .D(N177), .E(n1004), .CK(i_CLK), .Q(product[3])
         );
  fd1eqd1_hd product_reg_8_ ( .D(n1160), .E(n1004), .CK(i_CLK), .Q(product[8])
         );
  fd1eqd1_hd product_reg_12_ ( .D(n1155), .E(n1004), .CK(i_CLK), .Q(
        product[12]) );
  fd1eqd1_hd product_reg_13_ ( .D(n1153), .E(n1004), .CK(i_CLK), .Q(
        product[13]) );
  fd1eqd1_hd product_reg_14_ ( .D(n1152), .E(n1004), .CK(i_CLK), .Q(
        product[14]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1019), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n1018), .CK(i_CLK), .Q(b[30]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n262), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n261), .CK(i_CLK), .Q(z_m[22]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n263), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n264), .CK(i_CLK), .Q(z_m[19]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n1018), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n1018), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n1018), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n1018), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n1018), .CK(i_CLK), .Q(b[28]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n1018), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd guard_reg ( .D(n104), .E(n105), .CK(i_CLK), .Q(net922) );
  fd1qd1_hd z_m_reg_16_ ( .D(n267), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n269), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n265), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n320), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n311), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n270), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n266), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n268), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n319), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n356), .CK(i_CLK), .Q(b_e[9]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n1018), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n1018), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n1018), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n1018), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n1018), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n1018), .CK(i_CLK), .Q(b[26]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n1018), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n1018), .CK(i_CLK), .Q(b[23]) );
  fd1eqd1_hd z_e_reg_8_ ( .D(N474), .E(n110), .CK(i_CLK), .Q(z_e[8]) );
  fd1eqd1_hd z_e_reg_9_ ( .D(N475), .E(n110), .CK(i_CLK), .Q(z_e[9]) );
  fd1eqd1_hd z_e_reg_2_ ( .D(N468), .E(n110), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n286), .CK(i_CLK), .Q(z_m[23]) );
  fd1eqd1_hd z_e_reg_7_ ( .D(N473), .E(n110), .CK(i_CLK), .Q(z_e[7]) );
  fd1eqd1_hd z_e_reg_1_ ( .D(N467), .E(n110), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n323), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n314), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n322), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n321), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n313), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n312), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n275), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n271), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n273), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n274), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n276), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n272), .CK(i_CLK), .Q(z_m[11]) );
  fd1eqd1_hd z_e_reg_4_ ( .D(N470), .E(n110), .CK(i_CLK), .Q(z_e[4]) );
  fd1eqd1_hd z_e_reg_6_ ( .D(N472), .E(n110), .CK(i_CLK), .Q(z_e[6]) );
  fd1eqd1_hd z_e_reg_3_ ( .D(N469), .E(n110), .CK(i_CLK), .Q(z_e[3]) );
  fd1eqd1_hd z_e_reg_5_ ( .D(N471), .E(n110), .CK(i_CLK), .Q(z_e[5]) );
  fd1eqd1_hd z_e_reg_0_ ( .D(n2863), .E(n110), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n325), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n281), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n324), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n316), .CK(i_CLK), .Q(a_e[2]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n315), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n282), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n279), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n277), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n326), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n317), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n278), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n280), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n327), .CK(i_CLK), .Q(b_e[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n318), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd state_reg_3_ ( .D(n357), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd state_reg_0_ ( .D(n353), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd state_reg_2_ ( .D(n351), .CK(i_CLK), .Q(state[2]) );
  fad1_hd DP_OP_125J3_130_6300_U10 ( .A(n1103), .B(n2865), .CI(
        DP_OP_125J3_130_6300_n25), .CO(DP_OP_125J3_130_6300_n9), .S(N467) );
  ivd1_hd U511 ( .A(N34), .Y(n1220) );
  fad1_hd intadd_6_U15 ( .A(intadd_6_A_0_), .B(intadd_6_B_0_), .CI(intadd_6_CI), .CO(intadd_6_n14), .S(intadd_6_SUM_0_) );
  fad1_hd intadd_6_U14 ( .A(intadd_6_A_1_), .B(intadd_6_B_1_), .CI(
        intadd_6_n14), .CO(intadd_6_n13), .S(intadd_6_SUM_1_) );
  fad1_hd intadd_6_U13 ( .A(intadd_6_A_2_), .B(intadd_6_B_2_), .CI(
        intadd_6_n13), .CO(intadd_6_n12), .S(intadd_6_SUM_2_) );
  fad1_hd intadd_6_U12 ( .A(intadd_6_A_3_), .B(intadd_6_B_3_), .CI(
        intadd_6_n12), .CO(intadd_6_n11), .S(intadd_6_SUM_3_) );
  fad1_hd intadd_6_U11 ( .A(intadd_6_A_4_), .B(intadd_6_B_4_), .CI(
        intadd_6_n11), .CO(intadd_6_n10), .S(intadd_6_SUM_4_) );
  fad1_hd intadd_6_U10 ( .A(intadd_6_A_5_), .B(intadd_6_B_5_), .CI(
        intadd_6_n10), .CO(intadd_6_n9), .S(intadd_6_SUM_5_) );
  fad1_hd intadd_6_U9 ( .A(intadd_6_A_6_), .B(intadd_6_B_6_), .CI(intadd_6_n9), 
        .CO(intadd_6_n8), .S(intadd_6_SUM_6_) );
  fad1_hd intadd_6_U8 ( .A(intadd_6_A_7_), .B(intadd_6_B_7_), .CI(intadd_6_n8), 
        .CO(intadd_6_n7), .S(intadd_6_SUM_7_) );
  fad1_hd intadd_6_U7 ( .A(intadd_6_A_8_), .B(intadd_6_B_8_), .CI(intadd_6_n7), 
        .CO(intadd_6_n6), .S(intadd_6_SUM_8_) );
  fad1_hd intadd_6_U6 ( .A(intadd_6_A_9_), .B(intadd_6_B_9_), .CI(intadd_6_n6), 
        .CO(intadd_6_n5), .S(intadd_6_SUM_9_) );
  fad1_hd intadd_6_U5 ( .A(intadd_6_A_10_), .B(intadd_6_B_10_), .CI(
        intadd_6_n5), .CO(intadd_6_n4), .S(intadd_6_SUM_10_) );
  fad1_hd intadd_6_U4 ( .A(intadd_6_A_11_), .B(intadd_6_B_11_), .CI(
        intadd_6_n4), .CO(intadd_6_n3), .S(intadd_6_SUM_11_) );
  fad1_hd intadd_6_U3 ( .A(intadd_8_n1), .B(intadd_6_B_12_), .CI(intadd_6_n3), 
        .CO(intadd_6_n2), .S(intadd_6_SUM_12_) );
  fad1_hd intadd_6_U2 ( .A(intadd_6_A_13_), .B(intadd_6_B_13_), .CI(
        intadd_6_n2), .CO(intadd_6_n1), .S(intadd_6_SUM_13_) );
  fad1_hd intadd_7_U12 ( .A(intadd_7_A_0_), .B(intadd_7_B_0_), .CI(intadd_7_CI), .CO(intadd_7_n11), .S(intadd_7_SUM_0_) );
  fad1_hd intadd_7_U11 ( .A(intadd_7_A_1_), .B(intadd_7_B_1_), .CI(
        intadd_7_n11), .CO(intadd_7_n10), .S(intadd_7_SUM_1_) );
  fad1_hd intadd_7_U10 ( .A(intadd_7_A_2_), .B(intadd_7_B_2_), .CI(
        intadd_7_n10), .CO(intadd_7_n9), .S(intadd_7_SUM_2_) );
  fad1_hd intadd_7_U9 ( .A(intadd_7_A_3_), .B(intadd_6_SUM_0_), .CI(
        intadd_7_n9), .CO(intadd_7_n8), .S(intadd_7_SUM_3_) );
  fad1_hd intadd_7_U8 ( .A(intadd_7_A_4_), .B(intadd_6_SUM_1_), .CI(
        intadd_7_n8), .CO(intadd_7_n7), .S(intadd_7_SUM_4_) );
  fad1_hd intadd_7_U7 ( .A(intadd_7_A_5_), .B(intadd_6_SUM_2_), .CI(
        intadd_7_n7), .CO(intadd_7_n6), .S(intadd_7_SUM_5_) );
  fad1_hd intadd_7_U6 ( .A(intadd_7_A_6_), .B(intadd_6_SUM_3_), .CI(
        intadd_7_n6), .CO(intadd_7_n5), .S(intadd_7_SUM_6_) );
  fad1_hd intadd_7_U5 ( .A(intadd_7_A_7_), .B(intadd_6_SUM_4_), .CI(
        intadd_7_n5), .CO(intadd_7_n4), .S(intadd_7_SUM_7_) );
  fad1_hd intadd_7_U4 ( .A(intadd_7_A_8_), .B(intadd_6_SUM_5_), .CI(
        intadd_7_n4), .CO(intadd_7_n3), .S(intadd_7_SUM_8_) );
  fad1_hd intadd_7_U3 ( .A(intadd_6_SUM_6_), .B(intadd_7_B_9_), .CI(
        intadd_7_n3), .CO(intadd_7_n2), .S(intadd_7_SUM_9_) );
  fad1_hd intadd_7_U2 ( .A(intadd_7_A_10_), .B(intadd_6_SUM_7_), .CI(
        intadd_7_n2), .CO(intadd_7_n1), .S(intadd_7_SUM_10_) );
  fad1_hd intadd_8_U10 ( .A(intadd_8_A_0_), .B(intadd_8_B_0_), .CI(intadd_8_CI), .CO(intadd_8_n9), .S(intadd_6_B_3_) );
  fad1_hd intadd_8_U9 ( .A(intadd_8_A_1_), .B(intadd_8_B_1_), .CI(intadd_8_n9), 
        .CO(intadd_8_n8), .S(intadd_6_B_4_) );
  fad1_hd intadd_8_U8 ( .A(intadd_8_A_2_), .B(intadd_8_B_2_), .CI(intadd_8_n8), 
        .CO(intadd_8_n7), .S(intadd_6_B_5_) );
  fad1_hd intadd_8_U7 ( .A(n2022), .B(intadd_8_B_3_), .CI(intadd_8_n7), .CO(
        intadd_8_n6), .S(intadd_6_A_6_) );
  fad1_hd intadd_8_U6 ( .A(intadd_8_A_4_), .B(n2021), .CI(intadd_8_n6), .CO(
        intadd_8_n5), .S(intadd_6_B_7_) );
  fad1_hd intadd_8_U5 ( .A(n2020), .B(intadd_8_B_5_), .CI(intadd_8_n5), .CO(
        intadd_8_n4), .S(intadd_6_B_8_) );
  fad1_hd intadd_8_U4 ( .A(n1210), .B(intadd_8_B_6_), .CI(intadd_8_n4), .CO(
        intadd_8_n3), .S(intadd_6_A_9_) );
  fad1_hd intadd_8_U3 ( .A(n1208), .B(intadd_8_B_7_), .CI(intadd_8_n3), .CO(
        intadd_8_n2), .S(intadd_6_B_10_) );
  fad1_hd intadd_8_U2 ( .A(n1201), .B(intadd_8_B_8_), .CI(intadd_8_n2), .CO(
        intadd_8_n1), .S(intadd_6_A_11_) );
  fad1_hd intadd_10_U9 ( .A(a_m[5]), .B(a_m[2]), .CI(intadd_10_CI), .CO(
        intadd_10_n8), .S(intadd_10_SUM_0_) );
  fad1_hd intadd_10_U8 ( .A(n1225), .B(intadd_10_B_1_), .CI(intadd_10_n8), 
        .CO(intadd_10_n7), .S(intadd_10_SUM_1_) );
  fad1_hd intadd_10_U7 ( .A(intadd_10_A_2_), .B(intadd_10_B_2_), .CI(
        intadd_10_n7), .CO(intadd_10_n6), .S(intadd_10_SUM_2_) );
  fad1_hd intadd_10_U6 ( .A(intadd_10_A_3_), .B(intadd_10_B_3_), .CI(
        intadd_10_n6), .CO(intadd_10_n5), .S(intadd_10_SUM_3_) );
  fad1_hd intadd_10_U5 ( .A(intadd_10_A_4_), .B(intadd_10_B_4_), .CI(
        intadd_10_n5), .CO(intadd_10_n4), .S(intadd_10_SUM_4_) );
  fad1_hd intadd_10_U4 ( .A(intadd_10_A_5_), .B(n1206), .CI(intadd_10_n4), 
        .CO(intadd_10_n3), .S(intadd_10_SUM_5_) );
  fad1_hd intadd_10_U3 ( .A(n1204), .B(intadd_10_B_6_), .CI(intadd_10_n3), 
        .CO(intadd_10_n2), .S(intadd_10_SUM_6_) );
  fad1_hd intadd_10_U2 ( .A(n1197), .B(intadd_10_B_7_), .CI(intadd_10_n2), 
        .CO(intadd_10_n1), .S(intadd_10_SUM_7_) );
  fad1_hd intadd_11_U7 ( .A(n1222), .B(intadd_11_B_0_), .CI(intadd_11_CI), 
        .CO(intadd_11_n6), .S(intadd_11_SUM_0_) );
  fad1_hd intadd_11_U6 ( .A(intadd_11_A_1_), .B(intadd_11_B_1_), .CI(
        intadd_11_n6), .CO(intadd_11_n5), .S(intadd_11_SUM_1_) );
  fad1_hd intadd_11_U5 ( .A(intadd_11_A_2_), .B(intadd_11_B_2_), .CI(
        intadd_11_n5), .CO(intadd_11_n4), .S(intadd_11_SUM_2_) );
  fad1_hd intadd_11_U4 ( .A(intadd_11_A_3_), .B(intadd_11_B_3_), .CI(
        intadd_11_n4), .CO(intadd_11_n3), .S(intadd_11_SUM_3_) );
  fad1_hd intadd_11_U3 ( .A(intadd_11_A_4_), .B(n1194), .CI(intadd_11_n3), 
        .CO(intadd_11_n2), .S(intadd_11_SUM_4_) );
  fad1_hd intadd_12_U6 ( .A(n2034), .B(intadd_12_B_0_), .CI(intadd_12_CI), 
        .CO(intadd_12_n5), .S(intadd_12_SUM_0_) );
  fad1_hd intadd_12_U5 ( .A(intadd_12_A_1_), .B(intadd_12_B_1_), .CI(
        intadd_12_n5), .CO(intadd_12_n4), .S(intadd_12_SUM_1_) );
  fad1_hd intadd_12_U4 ( .A(n1202), .B(intadd_12_B_2_), .CI(intadd_12_n4), 
        .CO(intadd_12_n3), .S(intadd_12_SUM_2_) );
  fad1_hd intadd_12_U3 ( .A(n1188), .B(n1193), .CI(intadd_12_n3), .CO(
        intadd_12_n2), .S(intadd_12_SUM_3_) );
  fad1_hd intadd_13_U4 ( .A(intadd_13_A_0_), .B(intadd_13_B_0_), .CI(
        intadd_13_CI), .CO(intadd_13_n3), .S(intadd_13_SUM_0_) );
  fad1_hd intadd_13_U3 ( .A(intadd_13_A_1_), .B(intadd_13_B_1_), .CI(
        intadd_13_n3), .CO(intadd_13_n2), .S(intadd_13_SUM_1_) );
  fad1_hd intadd_14_U4 ( .A(a_m[2]), .B(intadd_14_B_0_), .CI(intadd_14_CI), 
        .CO(intadd_14_n3), .S(intadd_14_SUM_0_) );
  fad1_hd intadd_14_U3 ( .A(intadd_14_A_1_), .B(n1224), .CI(intadd_14_n3), 
        .CO(intadd_14_n2), .S(intadd_14_SUM_1_) );
  fad1_hd intadd_14_U2 ( .A(n1211), .B(intadd_14_B_2_), .CI(intadd_14_n2), 
        .CO(intadd_14_n1), .S(intadd_14_SUM_2_) );
  fad1_hd intadd_15_U3 ( .A(intadd_15_A_1_), .B(intadd_15_B_1_), .CI(
        intadd_15_n3), .CO(intadd_15_n2), .S(intadd_15_SUM_1_) );
  fad1_hd intadd_15_U2 ( .A(intadd_15_A_2_), .B(intadd_15_B_2_), .CI(
        intadd_15_n2), .CO(intadd_15_n1), .S(intadd_15_SUM_2_) );
  fad1_hd intadd_16_U4 ( .A(intadd_16_A_0_), .B(intadd_16_B_0_), .CI(
        intadd_11_SUM_1_), .CO(intadd_16_n3), .S(intadd_16_SUM_0_) );
  fad1_hd intadd_16_U3 ( .A(intadd_11_SUM_2_), .B(intadd_16_B_1_), .CI(
        intadd_16_n3), .CO(intadd_16_n2), .S(intadd_16_SUM_1_) );
  fad1_hd intadd_17_U4 ( .A(intadd_10_SUM_5_), .B(intadd_17_B_0_), .CI(
        intadd_17_CI), .CO(intadd_17_n3), .S(intadd_17_SUM_0_) );
  fad1_hd intadd_17_U3 ( .A(intadd_10_SUM_6_), .B(intadd_17_B_1_), .CI(
        intadd_17_n3), .CO(intadd_17_n2), .S(intadd_17_SUM_1_) );
  fad1_hd intadd_18_U4 ( .A(n1200), .B(intadd_18_B_0_), .CI(intadd_18_CI), 
        .CO(intadd_18_n3), .S(intadd_6_B_12_) );
  fad1_hd intadd_18_U3 ( .A(n1199), .B(intadd_18_B_1_), .CI(intadd_18_n3), 
        .CO(intadd_18_n2), .S(intadd_6_A_13_) );
  fad1_hd intadd_19_U4 ( .A(intadd_10_SUM_2_), .B(intadd_19_B_0_), .CI(
        intadd_19_CI), .CO(intadd_19_n3), .S(intadd_19_SUM_0_) );
  fad1_hd intadd_19_U3 ( .A(intadd_10_SUM_3_), .B(intadd_19_B_1_), .CI(
        intadd_19_n3), .CO(intadd_19_n2), .S(intadd_19_SUM_1_) );
  fad1_hd intadd_19_U2 ( .A(intadd_10_SUM_4_), .B(intadd_19_B_2_), .CI(
        intadd_19_n2), .CO(intadd_19_n1), .S(intadd_19_SUM_2_) );
  fad1_hd intadd_20_U4 ( .A(intadd_20_A_0_), .B(intadd_6_SUM_9_), .CI(
        intadd_20_CI), .CO(intadd_20_n3), .S(intadd_20_SUM_0_) );
  fad1_hd intadd_20_U3 ( .A(intadd_20_A_1_), .B(intadd_6_SUM_10_), .CI(
        intadd_20_n3), .CO(intadd_20_n2), .S(intadd_20_SUM_1_) );
  fad1_hd intadd_20_U2 ( .A(intadd_6_SUM_11_), .B(intadd_20_B_2_), .CI(
        intadd_20_n2), .CO(intadd_20_n1), .S(intadd_20_SUM_2_) );
  fad1_hd intadd_0_U26 ( .A(intadd_0_A_0_), .B(intadd_0_B_0_), .CI(intadd_0_CI), .CO(intadd_0_n25), .S(intadd_0_SUM_0_) );
  fad1_hd intadd_0_U25 ( .A(intadd_0_A_1_), .B(intadd_0_B_1_), .CI(
        intadd_0_n25), .CO(intadd_0_n24), .S(intadd_0_SUM_1_) );
  fad1_hd intadd_0_U24 ( .A(intadd_0_A_2_), .B(intadd_0_B_2_), .CI(
        intadd_0_n24), .CO(intadd_0_n23), .S(intadd_0_SUM_2_) );
  fad1_hd intadd_0_U23 ( .A(intadd_0_A_3_), .B(intadd_0_B_3_), .CI(
        intadd_0_n23), .CO(intadd_0_n22), .S(intadd_0_SUM_3_) );
  fad1_hd intadd_0_U22 ( .A(intadd_0_A_4_), .B(intadd_0_B_4_), .CI(
        intadd_0_n22), .CO(intadd_0_n21), .S(intadd_0_SUM_4_) );
  fad1_hd intadd_0_U21 ( .A(intadd_0_A_5_), .B(intadd_0_B_5_), .CI(
        intadd_0_n21), .CO(intadd_0_n20), .S(intadd_0_SUM_5_) );
  fad1_hd intadd_0_U20 ( .A(intadd_0_A_6_), .B(intadd_0_B_6_), .CI(
        intadd_0_n20), .CO(intadd_0_n19), .S(intadd_0_SUM_6_) );
  fad1_hd intadd_0_U19 ( .A(intadd_0_A_7_), .B(intadd_0_B_7_), .CI(
        intadd_0_n19), .CO(intadd_0_n18), .S(intadd_0_SUM_7_) );
  fad1_hd intadd_0_U18 ( .A(intadd_0_A_8_), .B(intadd_0_B_8_), .CI(
        intadd_0_n18), .CO(intadd_0_n17), .S(intadd_0_SUM_8_) );
  fad1_hd intadd_0_U17 ( .A(intadd_0_A_9_), .B(intadd_0_B_9_), .CI(
        intadd_0_n17), .CO(intadd_0_n16), .S(intadd_0_SUM_9_) );
  fad1_hd intadd_0_U16 ( .A(intadd_0_A_10_), .B(intadd_0_B_10_), .CI(
        intadd_0_n16), .CO(intadd_0_n15), .S(intadd_0_SUM_10_) );
  fad1_hd intadd_0_U15 ( .A(intadd_0_A_11_), .B(intadd_0_B_11_), .CI(
        intadd_0_n15), .CO(intadd_0_n14), .S(intadd_0_SUM_11_) );
  fad1_hd intadd_0_U14 ( .A(intadd_0_A_12_), .B(intadd_0_B_12_), .CI(
        intadd_0_n14), .CO(intadd_0_n13), .S(intadd_0_SUM_12_) );
  fad1_hd intadd_0_U13 ( .A(intadd_0_A_13_), .B(intadd_0_B_13_), .CI(
        intadd_0_n13), .CO(intadd_0_n12), .S(intadd_0_SUM_13_) );
  fad1_hd intadd_0_U12 ( .A(intadd_0_A_14_), .B(intadd_0_B_14_), .CI(
        intadd_0_n12), .CO(intadd_0_n11), .S(intadd_0_SUM_14_) );
  fad1_hd intadd_0_U11 ( .A(intadd_0_A_15_), .B(intadd_0_B_15_), .CI(
        intadd_0_n11), .CO(intadd_0_n10), .S(intadd_0_SUM_15_) );
  fad1_hd intadd_0_U10 ( .A(intadd_0_A_16_), .B(intadd_0_B_16_), .CI(
        intadd_0_n10), .CO(intadd_0_n9), .S(intadd_0_SUM_16_) );
  fad1_hd intadd_0_U9 ( .A(intadd_0_A_17_), .B(intadd_0_B_17_), .CI(
        intadd_0_n9), .CO(intadd_0_n8), .S(intadd_0_SUM_17_) );
  fad1_hd intadd_0_U8 ( .A(intadd_0_A_18_), .B(intadd_0_B_18_), .CI(
        intadd_0_n8), .CO(intadd_0_n7), .S(intadd_0_SUM_18_) );
  fad1_hd intadd_0_U7 ( .A(intadd_0_A_19_), .B(intadd_0_B_19_), .CI(
        intadd_0_n7), .CO(intadd_0_n6), .S(intadd_0_SUM_19_) );
  fad1_hd intadd_0_U6 ( .A(intadd_0_A_20_), .B(intadd_0_B_20_), .CI(
        intadd_0_n6), .CO(intadd_0_n5), .S(intadd_0_SUM_20_) );
  fad1_hd intadd_1_U21 ( .A(a_m[2]), .B(intadd_1_B_0_), .CI(intadd_1_CI), .CO(
        intadd_1_n20), .S(intadd_1_SUM_0_) );
  fad1_hd intadd_1_U20 ( .A(n2033), .B(intadd_14_SUM_0_), .CI(intadd_1_n20), 
        .CO(intadd_1_n19), .S(intadd_1_SUM_1_) );
  fad1_hd intadd_1_U19 ( .A(intadd_14_SUM_1_), .B(intadd_1_B_2_), .CI(
        intadd_1_n19), .CO(intadd_1_n18), .S(intadd_1_SUM_2_) );
  fad1_hd intadd_1_U18 ( .A(intadd_14_SUM_2_), .B(intadd_1_B_3_), .CI(
        intadd_1_n18), .CO(intadd_1_n17), .S(intadd_1_SUM_3_) );
  fad1_hd intadd_1_U17 ( .A(intadd_14_n1), .B(n1205), .CI(intadd_1_n17), .CO(
        intadd_1_n16), .S(intadd_1_SUM_4_) );
  fad1_hd intadd_1_U16 ( .A(n1203), .B(intadd_1_B_5_), .CI(intadd_1_n16), .CO(
        intadd_1_n15), .S(intadd_1_SUM_5_) );
  fad1_hd intadd_1_U15 ( .A(n1196), .B(intadd_1_B_6_), .CI(intadd_1_n15), .CO(
        intadd_1_n14), .S(intadd_1_SUM_6_) );
  fad1_hd intadd_1_U14 ( .A(n1195), .B(n1192), .CI(intadd_1_n14), .CO(
        intadd_1_n13), .S(intadd_1_SUM_7_) );
  fad1_hd intadd_2_U20 ( .A(intadd_2_A_0_), .B(intadd_2_B_0_), .CI(intadd_2_CI), .CO(intadd_2_n19), .S(intadd_0_A_3_) );
  fad1_hd intadd_2_U19 ( .A(intadd_2_A_1_), .B(intadd_2_B_1_), .CI(
        intadd_2_n19), .CO(intadd_2_n18), .S(intadd_0_A_4_) );
  fad1_hd intadd_2_U18 ( .A(intadd_2_A_2_), .B(intadd_2_B_2_), .CI(
        intadd_2_n18), .CO(intadd_2_n17), .S(intadd_0_A_5_) );
  fad1_hd intadd_2_U17 ( .A(intadd_2_A_3_), .B(intadd_2_B_3_), .CI(
        intadd_2_n17), .CO(intadd_2_n16), .S(intadd_0_A_6_) );
  fad1_hd intadd_2_U16 ( .A(intadd_2_A_4_), .B(intadd_2_B_4_), .CI(
        intadd_2_n16), .CO(intadd_2_n15), .S(intadd_0_A_7_) );
  fad1_hd intadd_2_U15 ( .A(intadd_2_A_5_), .B(intadd_2_B_5_), .CI(
        intadd_2_n15), .CO(intadd_2_n14), .S(intadd_0_A_8_) );
  fad1_hd intadd_2_U14 ( .A(intadd_2_A_6_), .B(intadd_2_B_6_), .CI(
        intadd_2_n14), .CO(intadd_2_n13), .S(intadd_0_A_9_) );
  fad1_hd intadd_2_U13 ( .A(intadd_2_A_7_), .B(intadd_2_B_7_), .CI(
        intadd_2_n13), .CO(intadd_2_n12), .S(intadd_0_A_10_) );
  fad1_hd intadd_2_U12 ( .A(intadd_2_A_8_), .B(intadd_2_B_8_), .CI(
        intadd_2_n12), .CO(intadd_2_n11), .S(intadd_0_A_11_) );
  fad1_hd intadd_2_U11 ( .A(intadd_2_A_9_), .B(intadd_2_B_9_), .CI(
        intadd_2_n11), .CO(intadd_2_n10), .S(intadd_0_A_12_) );
  fad1_hd intadd_2_U10 ( .A(intadd_2_A_10_), .B(intadd_2_B_10_), .CI(
        intadd_2_n10), .CO(intadd_2_n9), .S(intadd_0_A_13_) );
  fad1_hd intadd_2_U8 ( .A(intadd_2_A_12_), .B(intadd_2_B_12_), .CI(
        intadd_2_n8), .CO(intadd_2_n7), .S(intadd_0_A_15_) );
  fad1_hd intadd_2_U7 ( .A(intadd_2_A_13_), .B(intadd_2_B_13_), .CI(
        intadd_2_n7), .CO(intadd_2_n6), .S(intadd_0_A_16_) );
  fad1_hd intadd_2_U6 ( .A(intadd_2_A_14_), .B(intadd_2_B_14_), .CI(
        intadd_2_n6), .CO(intadd_2_n5), .S(intadd_0_A_17_) );
  fad1_hd intadd_2_U5 ( .A(intadd_2_A_15_), .B(intadd_2_B_15_), .CI(
        intadd_2_n5), .CO(intadd_2_n4), .S(intadd_0_A_18_) );
  fad1_hd intadd_2_U4 ( .A(intadd_2_A_16_), .B(intadd_2_B_16_), .CI(
        intadd_2_n4), .CO(intadd_2_n3), .S(intadd_0_A_19_) );
  fad1_hd intadd_2_U3 ( .A(intadd_2_A_17_), .B(intadd_2_B_17_), .CI(
        intadd_2_n3), .CO(intadd_2_n2), .S(intadd_0_A_20_) );
  fad1_hd intadd_2_U2 ( .A(intadd_2_A_18_), .B(intadd_2_B_18_), .CI(
        intadd_2_n2), .CO(intadd_2_n1), .S(intadd_0_A_21_) );
  fad1_hd intadd_4_U18 ( .A(intadd_4_A_0_), .B(intadd_4_B_0_), .CI(intadd_4_CI), .CO(intadd_4_n17), .S(intadd_2_A_3_) );
  fad1_hd intadd_4_U17 ( .A(intadd_4_A_1_), .B(intadd_4_B_1_), .CI(
        intadd_4_n17), .CO(intadd_4_n16), .S(intadd_2_A_4_) );
  fad1_hd intadd_4_U16 ( .A(intadd_4_A_2_), .B(intadd_4_B_2_), .CI(
        intadd_4_n16), .CO(intadd_4_n15), .S(intadd_2_A_5_) );
  fad1_hd intadd_4_U15 ( .A(intadd_4_A_3_), .B(intadd_4_B_3_), .CI(
        intadd_4_n15), .CO(intadd_4_n14), .S(intadd_2_A_6_) );
  fad1_hd intadd_4_U14 ( .A(intadd_4_A_4_), .B(intadd_4_B_4_), .CI(
        intadd_4_n14), .CO(intadd_4_n13), .S(intadd_2_A_7_) );
  fad1_hd intadd_4_U13 ( .A(intadd_4_A_5_), .B(intadd_4_B_5_), .CI(
        intadd_4_n13), .CO(intadd_4_n12), .S(intadd_2_A_8_) );
  fad1_hd intadd_4_U12 ( .A(intadd_4_A_6_), .B(intadd_4_B_6_), .CI(
        intadd_4_n12), .CO(intadd_4_n11), .S(intadd_2_A_9_) );
  fad1_hd intadd_4_U11 ( .A(intadd_4_A_7_), .B(intadd_4_B_7_), .CI(
        intadd_4_n11), .CO(intadd_4_n10), .S(intadd_2_B_10_) );
  fad1_hd intadd_4_U10 ( .A(intadd_4_A_8_), .B(intadd_4_B_8_), .CI(
        intadd_4_n10), .CO(intadd_4_n9), .S(intadd_2_A_11_) );
  fad1_hd intadd_4_U9 ( .A(intadd_4_A_9_), .B(intadd_4_B_9_), .CI(intadd_4_n9), 
        .CO(intadd_4_n8), .S(intadd_2_A_12_) );
  fad1_hd intadd_4_U8 ( .A(intadd_4_A_10_), .B(intadd_4_B_10_), .CI(
        intadd_4_n8), .CO(intadd_4_n7), .S(intadd_2_B_13_) );
  fad1_hd intadd_4_U7 ( .A(intadd_4_A_11_), .B(intadd_4_B_11_), .CI(
        intadd_4_n7), .CO(intadd_4_n6), .S(intadd_2_A_14_) );
  fad1_hd intadd_4_U6 ( .A(intadd_4_A_12_), .B(intadd_4_B_12_), .CI(
        intadd_4_n6), .CO(intadd_4_n5), .S(intadd_2_A_15_) );
  fad1_hd intadd_4_U5 ( .A(intadd_4_A_13_), .B(intadd_4_B_13_), .CI(
        intadd_4_n5), .CO(intadd_4_n4), .S(intadd_2_A_16_) );
  fad1_hd intadd_4_U4 ( .A(intadd_4_A_14_), .B(intadd_4_B_14_), .CI(
        intadd_4_n4), .CO(intadd_4_n3), .S(intadd_2_A_17_) );
  fad1_hd intadd_4_U3 ( .A(intadd_4_A_15_), .B(intadd_4_B_15_), .CI(
        intadd_4_n3), .CO(intadd_4_n2), .S(intadd_2_B_18_) );
  fad1_hd intadd_4_U2 ( .A(intadd_4_A_16_), .B(intadd_4_B_16_), .CI(
        intadd_4_n2), .CO(intadd_4_n1), .S(intadd_0_A_22_) );
  fad1_hd intadd_5_U18 ( .A(intadd_5_A_0_), .B(intadd_5_B_0_), .CI(intadd_5_CI), .CO(intadd_5_n17), .S(intadd_4_A_3_) );
  fad1_hd intadd_5_U17 ( .A(intadd_5_A_1_), .B(intadd_5_B_1_), .CI(
        intadd_5_n17), .CO(intadd_5_n16), .S(intadd_4_A_4_) );
  fad1_hd intadd_5_U16 ( .A(intadd_5_A_2_), .B(intadd_5_B_2_), .CI(
        intadd_5_n16), .CO(intadd_5_n15), .S(intadd_4_A_5_) );
  fad1_hd intadd_5_U15 ( .A(intadd_5_A_3_), .B(intadd_7_SUM_0_), .CI(
        intadd_5_n15), .CO(intadd_5_n14), .S(intadd_4_A_6_) );
  fad1_hd intadd_5_U14 ( .A(intadd_5_A_4_), .B(intadd_7_SUM_1_), .CI(
        intadd_5_n14), .CO(intadd_5_n13), .S(intadd_4_A_7_) );
  fad1_hd intadd_5_U13 ( .A(intadd_5_A_5_), .B(intadd_7_SUM_2_), .CI(
        intadd_5_n13), .CO(intadd_5_n12), .S(intadd_4_A_8_) );
  fad1_hd intadd_5_U12 ( .A(intadd_5_A_6_), .B(intadd_7_SUM_3_), .CI(
        intadd_5_n12), .CO(intadd_5_n11), .S(intadd_4_A_9_) );
  fad1_hd intadd_5_U11 ( .A(intadd_5_A_7_), .B(intadd_7_SUM_4_), .CI(
        intadd_5_n11), .CO(intadd_5_n10), .S(intadd_4_B_10_) );
  fad1_hd intadd_5_U10 ( .A(intadd_7_SUM_5_), .B(intadd_5_B_8_), .CI(
        intadd_5_n10), .CO(intadd_5_n9), .S(intadd_4_A_11_) );
  fad1_hd intadd_5_U9 ( .A(intadd_5_A_9_), .B(intadd_7_SUM_6_), .CI(
        intadd_5_n9), .CO(intadd_5_n8), .S(intadd_4_A_12_) );
  fad1_hd intadd_5_U8 ( .A(intadd_7_SUM_7_), .B(intadd_5_B_10_), .CI(
        intadd_5_n8), .CO(intadd_5_n7), .S(intadd_4_B_13_) );
  fad1_hd intadd_5_U7 ( .A(intadd_5_A_11_), .B(intadd_7_SUM_8_), .CI(
        intadd_5_n7), .CO(intadd_5_n6), .S(intadd_4_A_14_) );
  fad1_hd intadd_5_U6 ( .A(intadd_7_SUM_9_), .B(intadd_5_B_12_), .CI(
        intadd_5_n6), .CO(intadd_5_n5), .S(intadd_4_B_15_) );
  fad1_hd intadd_5_U5 ( .A(intadd_5_A_13_), .B(intadd_7_SUM_10_), .CI(
        intadd_5_n5), .CO(intadd_5_n4), .S(intadd_4_A_16_) );
  fad1_hd intadd_5_U4 ( .A(intadd_7_n1), .B(intadd_5_B_14_), .CI(intadd_5_n4), 
        .CO(intadd_5_n3), .S(intadd_5_SUM_14_) );
  fad1_hd intadd_5_U3 ( .A(intadd_20_SUM_0_), .B(intadd_5_B_15_), .CI(
        intadd_5_n3), .CO(intadd_5_n2), .S(intadd_5_SUM_15_) );
  fad1_hd intadd_5_U2 ( .A(intadd_20_SUM_1_), .B(intadd_5_B_16_), .CI(
        intadd_5_n2), .CO(intadd_5_n1), .S(intadd_5_SUM_16_) );
  fd1d2_hd b_m_reg_0_ ( .D(n308), .CK(i_CLK), .Q(n7), .QN(n1009) );
  fad1_hd intadd_18_U2 ( .A(n1186), .B(intadd_18_B_2_), .CI(intadd_18_n2), 
        .CO(intadd_18_n1), .S(intadd_18_SUM_2_) );
  fad1_hd intadd_9_U9 ( .A(n1130), .B(intadd_9_B_0_), .CI(intadd_9_CI), .CO(
        intadd_9_n8), .S(intadd_9_SUM_0_) );
  fad1_hd intadd_0_U4 ( .A(intadd_0_A_22_), .B(intadd_2_n1), .CI(intadd_0_n4), 
        .CO(intadd_0_n3), .S(intadd_0_SUM_22_) );
  fd1qd1_hd z_reg_8_ ( .D(n252), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_7_ ( .D(n253), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n254), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_5_ ( .D(n255), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_4_ ( .D(n256), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n349), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n288), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n290), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n291), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n294), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n296), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n300), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n302), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n303), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n287), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n309), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n289), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n292), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n293), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n295), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n297), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n298), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n299), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n301), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n304), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n305), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n306), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n354), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n330), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n333), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n334), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n337), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n339), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n340), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n342), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n345), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n348), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n343), .CK(i_CLK), .Q(a_m[6]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n346), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n307), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n352), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n285), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_reg_22_ ( .D(n238), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd z_reg_30_ ( .D(n230), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n232), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n234), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n236), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n237), .CK(i_CLK), .Q(z[23]) );
  fad1_hd intadd_0_U5 ( .A(intadd_0_A_21_), .B(intadd_0_B_21_), .CI(
        intadd_0_n5), .CO(intadd_0_n4), .S(intadd_0_SUM_21_) );
  fad1_hd intadd_2_U9 ( .A(intadd_2_A_11_), .B(intadd_2_B_11_), .CI(
        intadd_2_n9), .CO(intadd_2_n8), .S(intadd_0_A_14_) );
  fd1qd1_hd a_m_reg_11_ ( .D(n338), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n332), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n341), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n344), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n347), .CK(i_CLK), .Q(a_m[2]) );
  fad1_hd DP_OP_116J3_127_7148_U6 ( .A(n1118), .B(n775), .CI(
        DP_OP_116J3_127_7148_n4), .CO(DP_OP_116J3_127_7148_n3), .S(C82_DATA2_6) );
  fad1_hd intadd_11_U2 ( .A(n1191), .B(intadd_11_B_5_), .CI(intadd_11_n2), 
        .CO(intadd_11_n1), .S(intadd_11_SUM_5_) );
  fad1_hd intadd_16_U2 ( .A(intadd_11_SUM_3_), .B(intadd_16_B_2_), .CI(
        intadd_16_n2), .CO(intadd_16_n1), .S(intadd_16_SUM_2_) );
  fad1_hd intadd_17_U2 ( .A(intadd_10_SUM_7_), .B(intadd_17_B_2_), .CI(
        intadd_17_n2), .CO(intadd_17_n1), .S(intadd_17_SUM_2_) );
  fad1_hd intadd_1_U13 ( .A(n1189), .B(intadd_1_B_8_), .CI(intadd_1_n13), .CO(
        intadd_1_n12), .S(intadd_1_SUM_8_) );
  fad1_hd DP_OP_125J3_130_6300_U9 ( .A(DP_OP_125J3_130_6300_n26), .B(n2865), 
        .CI(DP_OP_125J3_130_6300_n9), .CO(DP_OP_125J3_130_6300_n8), .S(N468)
         );
  fad1_hd DP_OP_125J3_130_6300_U8 ( .A(DP_OP_125J3_130_6300_n27), .B(n2865), 
        .CI(DP_OP_125J3_130_6300_n8), .CO(DP_OP_125J3_130_6300_n7), .S(N469)
         );
  fad1_hd DP_OP_125J3_130_6300_U7 ( .A(DP_OP_125J3_130_6300_n28), .B(n2865), 
        .CI(DP_OP_125J3_130_6300_n7), .CO(DP_OP_125J3_130_6300_n6), .S(N470)
         );
  fad1_hd DP_OP_125J3_130_6300_U6 ( .A(DP_OP_125J3_130_6300_n29), .B(n2865), 
        .CI(DP_OP_125J3_130_6300_n6), .CO(DP_OP_125J3_130_6300_n5), .S(N471)
         );
  fad1_hd DP_OP_125J3_130_6300_U5 ( .A(DP_OP_125J3_130_6300_n30), .B(n2865), 
        .CI(DP_OP_125J3_130_6300_n5), .CO(DP_OP_125J3_130_6300_n4), .S(N472)
         );
  fad1_hd DP_OP_125J3_130_6300_U4 ( .A(DP_OP_125J3_130_6300_n31), .B(n2865), 
        .CI(DP_OP_125J3_130_6300_n4), .CO(DP_OP_125J3_130_6300_n3), .S(N473)
         );
  fad1_hd DP_OP_125J3_130_6300_U3 ( .A(DP_OP_125J3_130_6300_n32), .B(n2865), 
        .CI(DP_OP_125J3_130_6300_n3), .CO(DP_OP_125J3_130_6300_n2), .S(N474)
         );
  fad1_hd intadd_13_U2 ( .A(n1187), .B(intadd_13_B_2_), .CI(intadd_13_n2), 
        .CO(intadd_13_n1), .S(intadd_13_SUM_2_) );
  fad1_hd intadd_12_U2 ( .A(n1190), .B(intadd_12_B_4_), .CI(intadd_12_n2), 
        .CO(intadd_12_n1), .S(intadd_12_SUM_4_) );
  fad1_hd intadd_15_U4 ( .A(n1221), .B(intadd_15_B_0_), .CI(intadd_15_CI), 
        .CO(intadd_15_n3), .S(intadd_15_SUM_0_) );
  fad1_hd intadd_3_U11 ( .A(n1038), .B(b_m[11]), .CI(intadd_3_n11), .CO(
        intadd_3_n10), .S(intadd_3_SUM_8_) );
  fad1_hd intadd_3_U12 ( .A(b_m[11]), .B(n1035), .CI(intadd_3_n12), .CO(
        intadd_3_n11), .S(intadd_3_SUM_7_) );
  fad1_hd intadd_3_U14 ( .A(b_m[9]), .B(n1032), .CI(intadd_3_n14), .CO(
        intadd_3_n13), .S(intadd_3_SUM_5_) );
  fad1_hd intadd_3_U13 ( .A(n1035), .B(b_m[9]), .CI(intadd_3_n13), .CO(
        intadd_3_n12), .S(intadd_3_SUM_6_) );
  fad1_hd intadd_3_U15 ( .A(n1032), .B(n1030), .CI(intadd_3_n15), .CO(
        intadd_3_n14), .S(intadd_3_SUM_4_) );
  fad1_hd intadd_3_U16 ( .A(n1030), .B(b_m[6]), .CI(intadd_3_n16), .CO(
        intadd_3_n15), .S(intadd_3_SUM_3_) );
  fad1_hd intadd_3_U17 ( .A(b_m[6]), .B(n1028), .CI(intadd_3_n17), .CO(
        intadd_3_n16), .S(intadd_3_SUM_2_) );
  fad1_hd intadd_3_U18 ( .A(n1028), .B(n1006), .CI(intadd_3_n18), .CO(
        intadd_3_n17), .S(intadd_3_SUM_1_) );
  fad1_hd intadd_3_U19 ( .A(n1006), .B(n1025), .CI(intadd_3_CI), .CO(
        intadd_3_n18), .S(intadd_3_SUM_0_) );
  fad1_hd intadd_0_U3 ( .A(intadd_0_A_23_), .B(intadd_4_n1), .CI(intadd_0_n3), 
        .CO(intadd_0_n2), .S(intadd_0_SUM_23_) );
  fad1_hd intadd_0_U2 ( .A(intadd_0_A_24_), .B(n1129), .CI(intadd_0_n2), .CO(
        intadd_0_n1), .S(intadd_0_SUM_24_) );
  fad1_hd intadd_1_U4 ( .A(n1185), .B(n2023), .CI(intadd_1_n4), .CO(
        intadd_1_n3), .S(N220) );
  fad1_hd intadd_1_U3 ( .A(n2032), .B(n1184), .CI(intadd_1_n3), .CO(
        intadd_1_n2), .S(N221) );
  fad1_hd intadd_1_U2 ( .A(n2031), .B(intadd_1_B_19_), .CI(intadd_1_n2), .CO(
        intadd_1_n1), .S(N222) );
  fad1_hd intadd_9_U7 ( .A(n1124), .B(n1125), .CI(intadd_9_n7), .CO(
        intadd_9_n6), .S(N206) );
  fad1_hd intadd_9_U6 ( .A(n2019), .B(n1123), .CI(intadd_9_n6), .CO(
        intadd_9_n5), .S(N207) );
  fad1_hd intadd_9_U5 ( .A(n1122), .B(n2018), .CI(intadd_9_n5), .CO(
        intadd_9_n4), .S(N208) );
  fad1_hd intadd_9_U4 ( .A(n1181), .B(n1121), .CI(intadd_9_n4), .CO(
        intadd_9_n3), .S(N209) );
  fad1_hd intadd_9_U3 ( .A(n2030), .B(n1180), .CI(intadd_9_n3), .CO(
        intadd_9_n2), .S(N210) );
  fad1_hd intadd_9_U2 ( .A(intadd_1_SUM_8_), .B(n2029), .CI(intadd_9_n2), .CO(
        intadd_9_n1), .S(N211) );
  fad1_hd intadd_1_U11 ( .A(n2028), .B(n1178), .CI(intadd_1_n11), .CO(
        intadd_1_n10), .S(N213) );
  fad1_hd intadd_1_U10 ( .A(intadd_12_SUM_4_), .B(n2027), .CI(intadd_1_n10), 
        .CO(intadd_1_n9), .S(N214) );
  fad1_hd intadd_1_U9 ( .A(n1177), .B(intadd_12_n1), .CI(intadd_1_n9), .CO(
        intadd_1_n8), .S(N215) );
  fad1_hd intadd_1_U8 ( .A(n2026), .B(n1176), .CI(intadd_1_n8), .CO(
        intadd_1_n7), .S(N216) );
  fad1_hd intadd_1_U7 ( .A(n1183), .B(n2025), .CI(intadd_1_n7), .CO(
        intadd_1_n6), .S(N217) );
  fad1_hd intadd_1_U6 ( .A(intadd_13_SUM_2_), .B(n1182), .CI(intadd_1_n6), 
        .CO(intadd_1_n5), .S(N218) );
  fad1_hd intadd_1_U5 ( .A(n2024), .B(intadd_13_n1), .CI(intadd_1_n5), .CO(
        intadd_1_n4), .S(N219) );
  fd1qd1_hd sticky_reg ( .D(n283), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n350), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd round_bit_reg ( .D(n284), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd o_Z_STB_reg ( .D(n358), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd a_m_reg_21_ ( .D(n328), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n331), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n336), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n310), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n355), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd z_reg_31_ ( .D(n229), .CK(i_CLK), .Q(z[31]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n335), .CK(i_CLK), .Q(a_m[14]) );
  fad1_hd intadd_1_U12 ( .A(n1179), .B(intadd_9_n1), .CI(intadd_1_n12), .CO(
        intadd_1_n11), .S(N212) );
  fad1_hd intadd_9_U8 ( .A(n1127), .B(n1126), .CI(intadd_9_n8), .CO(
        intadd_9_n7), .S(N205) );
  fad1_hd intadd_3_U5 ( .A(b_m[18]), .B(n1045), .CI(intadd_3_n5), .CO(
        intadd_3_n4), .S(intadd_3_SUM_14_) );
  fad1_hd intadd_3_U7 ( .A(n1008), .B(n1042), .CI(intadd_3_n7), .CO(
        intadd_3_n6), .S(intadd_3_SUM_12_) );
  fad1_hd intadd_3_U6 ( .A(n1045), .B(n1008), .CI(intadd_3_n6), .CO(
        intadd_3_n5), .S(intadd_3_SUM_13_) );
  fad1_hd intadd_3_U2 ( .A(n1052), .B(n1050), .CI(intadd_3_n2), .CO(
        intadd_3_n1), .S(intadd_3_SUM_17_) );
  fad1_hd intadd_3_U4 ( .A(n1048), .B(b_m[18]), .CI(intadd_3_n4), .CO(
        intadd_3_n3), .S(intadd_3_SUM_15_) );
  fad1_hd intadd_3_U3 ( .A(n1050), .B(n1048), .CI(intadd_3_n3), .CO(
        intadd_3_n2), .S(intadd_3_SUM_16_) );
  fad1_hd intadd_3_U10 ( .A(n1039), .B(n1038), .CI(intadd_3_n10), .CO(
        intadd_3_n9), .S(intadd_3_SUM_9_) );
  fad1_hd intadd_3_U9 ( .A(n1041), .B(n1039), .CI(intadd_3_n9), .CO(
        intadd_3_n8), .S(intadd_3_SUM_10_) );
  fad1_hd intadd_3_U8 ( .A(n1042), .B(n1041), .CI(intadd_3_n8), .CO(
        intadd_3_n7), .S(intadd_3_SUM_11_) );
  fd1qd1_hd a_m_reg_20_ ( .D(n329), .CK(i_CLK), .Q(a_m[20]) );
  ad2bd2_hd U367 ( .B(n1216), .AN(n1434), .Y(n1902) );
  clknd2d1_hd U368 ( .A(n1175), .B(n1857), .Y(n1148) );
  clknd2d1_hd U369 ( .A(a_m[0]), .B(n1061), .Y(n1158) );
  clknd2d1_hd U370 ( .A(n1058), .B(n7), .Y(n1909) );
  clknd2d1_hd U371 ( .A(n1432), .B(a_m[20]), .Y(n1420) );
  clknd2d1_hd U372 ( .A(n1058), .B(n1029), .Y(intadd_10_B_2_) );
  clknd2d1_hd U373 ( .A(n1058), .B(n1007), .Y(n1911) );
  clknd2d1_hd U374 ( .A(n1058), .B(n1028), .Y(intadd_10_CI) );
  clknd2d1_hd U375 ( .A(n1452), .B(a_m[17]), .Y(n1453) );
  clknd2d1_hd U376 ( .A(n7), .B(n1415), .Y(n1456) );
  clknd2d1_hd U377 ( .A(n1032), .B(intadd_10_A_2_), .Y(n1223) );
  clknd2d1_hd U378 ( .A(n7), .B(n1409), .Y(n1459) );
  clknd2d1_hd U379 ( .A(n1407), .B(a_m[14]), .Y(n1406) );
  clknd2d1_hd U380 ( .A(n1058), .B(n1038), .Y(intadd_11_B_1_) );
  clknd2d1_hd U381 ( .A(n1058), .B(n1034), .Y(n2034) );
  clknd2d1_hd U382 ( .A(n1058), .B(n1037), .Y(n1259) );
  clknd2d1_hd U383 ( .A(n1058), .B(n1524), .Y(n1219) );
  clknd2d1_hd U384 ( .A(n1033), .B(n1031), .Y(n1524) );
  clknd2d1_hd U385 ( .A(n7), .B(n1355), .Y(n1412) );
  clknd2d1_hd U386 ( .A(n1368), .B(a_m[11]), .Y(n1369) );
  clknd2d1_hd U387 ( .A(n1041), .B(intadd_11_A_1_), .Y(n1253) );
  clknd2d1_hd U388 ( .A(n7), .B(n1324), .Y(n1379) );
  clknd2d1_hd U389 ( .A(n1333), .B(a_m[8]), .Y(n1334) );
  clknd2d1_hd U390 ( .A(n1009), .B(n1022), .Y(n1070) );
  clknd2d1_hd U391 ( .A(n1024), .B(n1023), .Y(n1525) );
  clknd2d1_hd U392 ( .A(n1086), .B(n1088), .Y(n1487) );
  clknd2d1_hd U393 ( .A(n1058), .B(n1047), .Y(intadd_15_B_1_) );
  clknd2d1_hd U394 ( .A(n1046), .B(n1043), .Y(n1532) );
  clknd2d1_hd U395 ( .A(n1253), .B(n1252), .Y(n1254) );
  clknd2d1_hd U396 ( .A(n1355), .B(n1291), .Y(n1403) );
  clknd2d1_hd U397 ( .A(n1324), .B(n1312), .Y(n1357) );
  clknd2d1_hd U398 ( .A(n1056), .B(n1055), .Y(n1119) );
  clknd2d1_hd U399 ( .A(n1052), .B(intadd_3_n1), .Y(n1116) );
  clknd2d1_hd U400 ( .A(n1508), .B(n1507), .Y(n1522) );
  clknd2d1_hd U401 ( .A(n1747), .B(n1541), .Y(n1538) );
  clknd2d1_hd U402 ( .A(n1836), .B(n1539), .Y(n1540) );
  clknd2d1_hd U403 ( .A(n1763), .B(n1842), .Y(n1509) );
  clknd2d1_hd U404 ( .A(n1824), .B(n1534), .Y(n1812) );
  clknd2d1_hd U405 ( .A(n7), .B(n1168), .Y(n1344) );
  clknd2d1_hd U406 ( .A(n1165), .B(a_m[5]), .Y(n1090) );
  clknd2d1_hd U407 ( .A(n7), .B(n1086), .Y(n1213) );
  clknd2d1_hd U408 ( .A(n1495), .B(n1494), .Y(n1556) );
  clknd2d1_hd U409 ( .A(z_e[7]), .B(z_e[8]), .Y(n1555) );
  clknd2d1_hd U410 ( .A(n1054), .B(n1053), .Y(n1113) );
  clknd2d1_hd U411 ( .A(n1056), .B(n1198), .Y(n1145) );
  clknd2d1_hd U412 ( .A(n1049), .B(n1051), .Y(n1855) );
  ivd1_hd U413 ( .A(b_m[22]), .Y(n1055) );
  clknd2d1_hd U414 ( .A(n1290), .B(n1285), .Y(n1402) );
  clknd2d1_hd U415 ( .A(n1311), .B(n1293), .Y(n1356) );
  xo2d1_hd U416 ( .A(intadd_3_n1), .B(n1301), .Y(n1936) );
  xo2d1_hd U417 ( .A(n1132), .B(n1120), .Y(n1429) );
  clknd2d1_hd U418 ( .A(n1119), .B(n1117), .Y(n1120) );
  clknd2d1_hd U419 ( .A(n1116), .B(n1115), .Y(n1132) );
  clknd2d1_hd U420 ( .A(n1054), .B(n1057), .Y(n1117) );
  clknd2d1_hd U421 ( .A(n1824), .B(state[0]), .Y(n1060) );
  clknd2d1_hd U422 ( .A(n1822), .B(n1846), .Y(n1807) );
  clknd2d1_hd U423 ( .A(n1534), .B(state[1]), .Y(n1548) );
  nid2_hd U424 ( .A(a_m[23]), .Y(n1058) );
  ivd2_hd U425 ( .A(a_m[20]), .Y(n1891) );
  clknd2d1_hd U426 ( .A(n1118), .B(n1832), .Y(n1783) );
  clknd2d1_hd U427 ( .A(n105), .B(n1818), .Y(n1704) );
  clknd2d1_hd U428 ( .A(n1541), .B(n1540), .Y(n1542) );
  clknd2d1_hd U429 ( .A(n1539), .B(n1538), .Y(n1544) );
  ivd2_hd U430 ( .A(n1023), .Y(n1022) );
  nid2_hd U431 ( .A(n1791), .Y(n1013) );
  ivd2_hd U432 ( .A(a_m[14]), .Y(n1869) );
  ivd2_hd U433 ( .A(n1024), .Y(n1007) );
  ivd1_hd U434 ( .A(b_m[1]), .Y(n1023) );
  ivd1_hd U435 ( .A(b_m[2]), .Y(n1024) );
  ivd2_hd U436 ( .A(n1026), .Y(n1025) );
  ivd2_hd U437 ( .A(n1027), .Y(n1006) );
  ivd2_hd U438 ( .A(n1031), .Y(n1030) );
  ivd1_hd U439 ( .A(b_m[8]), .Y(n1033) );
  ivd2_hd U440 ( .A(n1036), .Y(n1035) );
  ivd2_hd U441 ( .A(n1040), .Y(n1039) );
  ivd2_hd U442 ( .A(n1043), .Y(n1042) );
  ivd2_hd U443 ( .A(n1044), .Y(n1008) );
  ivd2_hd U444 ( .A(n1049), .Y(n1048) );
  ivd2_hd U445 ( .A(n1053), .Y(n1052) );
  ivd2_hd U446 ( .A(n1055), .Y(n1054) );
  ivd1_hd U447 ( .A(b_m[7]), .Y(n1031) );
  ivd2_hd U448 ( .A(n1033), .Y(n1032) );
  nid2_hd U449 ( .A(b_m[12]), .Y(n1038) );
  nid2_hd U450 ( .A(b_m[14]), .Y(n1041) );
  ivd2_hd U451 ( .A(n1046), .Y(n1045) );
  ivd2_hd U452 ( .A(n1051), .Y(n1050) );
  clknd2d1_hd U453 ( .A(N34), .B(n1845), .Y(n1847) );
  clknd2d1_hd U454 ( .A(n1711), .B(n1666), .Y(n1674) );
  clknd2d1_hd U455 ( .A(n1711), .B(n1675), .Y(n1681) );
  clknd2d1_hd U456 ( .A(n1711), .B(n1648), .Y(n1656) );
  clknd2d1_hd U457 ( .A(n1711), .B(n1639), .Y(n1644) );
  clknd2d1_hd U458 ( .A(n1711), .B(n1657), .Y(n1662) );
  clknd2d1_hd U459 ( .A(n1497), .B(n1815), .Y(n1844) );
  clknd2d1_hd U460 ( .A(n1711), .B(n1612), .Y(n1620) );
  clknd2d1_hd U461 ( .A(n1711), .B(n1630), .Y(n1638) );
  clknd2d1_hd U462 ( .A(n1711), .B(n1621), .Y(n1626) );
  clknd2d1_hd U463 ( .A(n1711), .B(n1603), .Y(n1608) );
  clknd2d1_hd U464 ( .A(n1600), .B(n1598), .Y(n1714) );
  clknd2d1_hd U465 ( .A(n1711), .B(n1599), .Y(n1598) );
  or2d2_hd U466 ( .A(n1060), .B(n1807), .Y(n1118) );
  clknd2d1_hd U467 ( .A(n1068), .B(n1067), .Y(n1069) );
  clknd2d1_hd U468 ( .A(n1213), .B(n1069), .Y(n1074) );
  clknd2d1_hd U469 ( .A(n1073), .B(n1074), .Y(intadd_0_A_0_) );
  clknd2d1_hd U470 ( .A(n1582), .B(n1578), .Y(n1577) );
  clknd2d1_hd U471 ( .A(n1574), .B(n1571), .Y(n1570) );
  clknd2d1_hd U472 ( .A(n1567), .B(n1564), .Y(n1563) );
  clknd2d1_hd U473 ( .A(n1053), .B(n1057), .Y(n1526) );
  clknd2d1_hd U474 ( .A(n1055), .B(n1052), .Y(n1112) );
  clknd2d1_hd U475 ( .A(n1076), .B(n1113), .Y(n1075) );
  clknd2d1_hd U476 ( .A(n1113), .B(n1112), .Y(n1301) );
  clknd2d1_hd U477 ( .A(n1050), .B(intadd_15_A_1_), .Y(n1856) );
  clknd2d1_hd U478 ( .A(n1148), .B(n1145), .Y(n1150) );
  clknd2d1_hd U479 ( .A(state[3]), .B(n1822), .Y(n1809) );
  clknd2d1_hd U480 ( .A(state[1]), .B(state[0]), .Y(n1820) );
  clknd2d1_hd U481 ( .A(n1010), .B(n1550), .Y(n1551) );
  clknd2d1_hd U482 ( .A(n1011), .B(z[23]), .Y(n1585) );
  clknd2d1_hd U483 ( .A(n1011), .B(z[24]), .Y(n1583) );
  clknd2d1_hd U484 ( .A(n1011), .B(z[26]), .Y(n1575) );
  clknd2d1_hd U485 ( .A(n1011), .B(z[28]), .Y(n1568) );
  clknd2d1_hd U486 ( .A(z_e[7]), .B(n1563), .Y(n1561) );
  clknd2d1_hd U487 ( .A(n1011), .B(z[22]), .Y(n1590) );
  clknd2d1_hd U488 ( .A(state[2]), .B(state[3]), .Y(n1826) );
  clknd2d1_hd U489 ( .A(n1753), .B(n138), .Y(n317) );
  clknd2d1_hd U490 ( .A(n1769), .B(n148), .Y(n326) );
  clknd2d1_hd U491 ( .A(n1710), .B(n1689), .Y(n1692) );
  clknd2d1_hd U492 ( .A(n1690), .B(n1689), .Y(n1687) );
  clknd2d1_hd U493 ( .A(z_m[0]), .B(n1711), .Y(n1685) );
  clknd2d1_hd U494 ( .A(n1711), .B(n1814), .Y(n1718) );
  clknd2d1_hd U495 ( .A(z_m[23]), .B(n1593), .Y(n1501) );
  clknd2d1_hd U496 ( .A(n1840), .B(n1839), .Y(n1837) );
  clknd2d1_hd U497 ( .A(b_e[9]), .B(n1850), .Y(n1839) );
  clknd2d1_hd U498 ( .A(n1759), .B(n1758), .Y(n1756) );
  clknd2d1_hd U499 ( .A(n1752), .B(n138), .Y(n311) );
  clknd2d1_hd U500 ( .A(b_e[8]), .B(n1766), .Y(n1767) );
  clknd2d1_hd U501 ( .A(n1500), .B(n1712), .Y(n105) );
  clknd2d1_hd U502 ( .A(a_m[2]), .B(N176), .Y(n1063) );
  clknd2d1_hd U503 ( .A(n1586), .B(n1581), .Y(n235) );
  ivd1_hd U504 ( .A(intadd_0_n1), .Y(n1127) );
  ivd4_hd U505 ( .A(n1111), .Y(n1004) );
  clknd2d1_hd U506 ( .A(n1553), .B(n1843), .Y(n148) );
  clknd2d1_hd U507 ( .A(n1553), .B(n1762), .Y(n138) );
  ivd1_hd U508 ( .A(b_m[23]), .Y(n1057) );
  ivd1_hd U509 ( .A(b_m[17]), .Y(n1046) );
  ivd1_hd U510 ( .A(b_m[15]), .Y(n1043) );
  ivd1_hd U512 ( .A(b_m[3]), .Y(n1026) );
  scg16d2_hd U513 ( .A(n1116), .B(n1119), .C(n1091), .Y(n1857) );
  scg12d2_hd U514 ( .A(n1311), .B(n1312), .C(n1293), .Y(n1932) );
  nr2d2_hd U515 ( .A(n1096), .B(n1095), .Y(n1929) );
  ad2d2_hd U516 ( .A(n1434), .B(n1217), .Y(n1903) );
  oa22ad1_hd U517 ( .A(n1059), .B(a_m[22]), .C(a_m[22]), .D(n1059), .Y(n1216)
         );
  ivd1_hd U518 ( .A(b_m[10]), .Y(n1036) );
  ivd1_hd U519 ( .A(a_m[11]), .Y(n1938) );
  ivd1_hd U520 ( .A(b_m[21]), .Y(n1053) );
  ivd1_hd U521 ( .A(b_m[19]), .Y(n1049) );
  xo2d1_hd U522 ( .A(n1014), .B(n1093), .Y(n1099) );
  xo2d1_hd U523 ( .A(n1016), .B(n1136), .Y(intadd_0_B_19_) );
  xo2d1_hd U524 ( .A(n1014), .B(n1367), .Y(intadd_4_B_16_) );
  xo2d1_hd U525 ( .A(n1303), .B(n1302), .Y(intadd_1_B_19_) );
  xo2d1_hd U526 ( .A(n1014), .B(n1321), .Y(intadd_2_A_18_) );
  xo2d1_hd U527 ( .A(n1014), .B(n1332), .Y(intadd_2_B_17_) );
  xo2d1_hd U528 ( .A(n1013), .B(n1385), .Y(intadd_5_A_13_) );
  xo2d1_hd U529 ( .A(n1381), .B(n1380), .Y(intadd_4_CI) );
  xo2d1_hd U530 ( .A(n1414), .B(n1413), .Y(intadd_5_CI) );
  xo2d1_hd U531 ( .A(n1461), .B(n1460), .Y(intadd_7_CI) );
  xo2d1_hd U532 ( .A(n1215), .B(n1214), .Y(intadd_0_CI) );
  ivd2_hd U533 ( .A(n1357), .Y(n1935) );
  xo2d1_hd U534 ( .A(n1026), .B(n1071), .Y(n1475) );
  nid6_hd U535 ( .A(n2017), .Y(n1018) );
  xo2d1_hd U536 ( .A(n1013), .B(n1232), .Y(intadd_10_B_3_) );
  ivd2_hd U537 ( .A(n1403), .Y(n1875) );
  ad2d2_hd U538 ( .A(n1235), .B(n1415), .Y(n1918) );
  ivd2_hd U539 ( .A(n1487), .Y(n1364) );
  ivd2_hd U540 ( .A(n1158), .Y(n1175) );
  ad2d2_hd U541 ( .A(n1094), .B(n1096), .Y(n1491) );
  nr2d2_hd U542 ( .A(n1086), .B(n1085), .Y(n1366) );
  ivd1_hd U543 ( .A(b_m[20]), .Y(n1051) );
  ivd1_hd U544 ( .A(b_m[13]), .Y(n1040) );
  ivd1_hd U545 ( .A(a_m[17]), .Y(n1881) );
  ivd1_hd U546 ( .A(b_m[16]), .Y(n1044) );
  xo2d1_hd U547 ( .A(n1059), .B(n1275), .Y(intadd_15_B_2_) );
  xo2d1_hd U548 ( .A(n1015), .B(n1282), .Y(intadd_16_B_2_) );
  xo2d1_hd U549 ( .A(a_m[5]), .B(n1489), .Y(intadd_9_B_0_) );
  xo2d1_hd U550 ( .A(n1059), .B(n1859), .Y(n1861) );
  xo2d1_hd U551 ( .A(n1017), .B(n1430), .Y(intadd_6_B_13_) );
  xo2d1_hd U552 ( .A(a_m[20]), .B(n1267), .Y(intadd_13_B_2_) );
  xo2d1_hd U553 ( .A(n1013), .B(n1315), .Y(intadd_20_B_2_) );
  xo2d1_hd U554 ( .A(n1891), .B(n1256), .Y(intadd_11_B_5_) );
  xo2d1_hd U555 ( .A(n1013), .B(n1401), .Y(intadd_5_B_16_) );
  xo2d1_hd U556 ( .A(a_m[17]), .B(n1262), .Y(intadd_12_B_4_) );
  xo2d1_hd U557 ( .A(n1938), .B(n1295), .Y(intadd_18_B_2_) );
  xo2d1_hd U558 ( .A(n1869), .B(n1287), .Y(intadd_17_B_2_) );
  xo2d1_hd U559 ( .A(a_m[14]), .B(n1308), .Y(intadd_1_B_8_) );
  xo2d1_hd U560 ( .A(a_m[20]), .B(n1896), .Y(n1900) );
  xo2d1_hd U561 ( .A(a_m[8]), .B(n1931), .Y(n1941) );
  xo2d1_hd U562 ( .A(a_m[11]), .B(n1865), .Y(n1872) );
  xo2d1_hd U563 ( .A(a_m[14]), .B(n1877), .Y(n1884) );
  xo2d1_hd U564 ( .A(a_m[17]), .B(n1889), .Y(n1894) );
  xo2d1_hd U565 ( .A(n1891), .B(n1890), .Y(n1893) );
  xo2d1_hd U566 ( .A(n1059), .B(n1897), .Y(n1899) );
  xo2d1_hd U567 ( .A(n1015), .B(n1880), .Y(n1883) );
  xo2d1_hd U568 ( .A(a_m[8]), .B(n1492), .Y(intadd_9_CI) );
  xo2d1_hd U569 ( .A(n1869), .B(n1868), .Y(n1871) );
  xo2d1_hd U570 ( .A(n1017), .B(n1937), .Y(n1940) );
  xo2d1_hd U571 ( .A(n1016), .B(n1114), .Y(intadd_0_B_18_) );
  xo2d1_hd U572 ( .A(a_m[14]), .B(n1307), .Y(intadd_1_B_6_) );
  xo2d1_hd U573 ( .A(n1013), .B(n1097), .Y(n1098) );
  xo2d1_hd U574 ( .A(n1015), .B(n1241), .Y(intadd_10_B_7_) );
  xo2d1_hd U575 ( .A(n1017), .B(n1428), .Y(intadd_6_B_11_) );
  xo2d1_hd U576 ( .A(n1016), .B(n1110), .Y(intadd_0_B_17_) );
  xo2d1_hd U577 ( .A(n1891), .B(n1255), .Y(intadd_11_B_3_) );
  xo2d1_hd U578 ( .A(n1059), .B(n1276), .Y(intadd_15_CI) );
  xo2d1_hd U579 ( .A(n1016), .B(n1109), .Y(intadd_0_B_16_) );
  xo2d1_hd U580 ( .A(n1017), .B(n1313), .Y(intadd_20_A_1_) );
  xo2d1_hd U581 ( .A(n1869), .B(n1292), .Y(intadd_18_B_1_) );
  xo2d1_hd U582 ( .A(n1014), .B(n1331), .Y(intadd_2_B_16_) );
  xo2d1_hd U583 ( .A(n1891), .B(n1279), .Y(intadd_16_B_1_) );
  xo2d1_hd U584 ( .A(n1015), .B(n1284), .Y(intadd_17_B_1_) );
  xo2d1_hd U585 ( .A(n1058), .B(n1264), .Y(intadd_13_A_1_) );
  xo2d1_hd U586 ( .A(n1013), .B(n1352), .Y(intadd_4_A_15_) );
  xo2d1_hd U587 ( .A(n1058), .B(n1268), .Y(intadd_13_CI) );
  xo2d1_hd U588 ( .A(n1015), .B(n1288), .Y(intadd_17_CI) );
  xo2d1_hd U589 ( .A(n1869), .B(n1296), .Y(intadd_18_CI) );
  xo2d1_hd U590 ( .A(n1014), .B(n1330), .Y(intadd_2_B_15_) );
  xo2d1_hd U591 ( .A(n1891), .B(n1278), .Y(intadd_16_B_0_) );
  xo2d1_hd U592 ( .A(n1016), .B(n1108), .Y(intadd_0_B_15_) );
  xo2d1_hd U593 ( .A(n1017), .B(n1316), .Y(intadd_20_CI) );
  xo2d1_hd U594 ( .A(n1013), .B(n1362), .Y(intadd_4_B_14_) );
  xo2d1_hd U595 ( .A(n1869), .B(n1482), .Y(intadd_8_B_8_) );
  xo2d1_hd U596 ( .A(n1014), .B(n1329), .Y(intadd_2_B_14_) );
  xo2d1_hd U597 ( .A(a_m[20]), .B(n1261), .Y(intadd_12_B_2_) );
  xo2d1_hd U598 ( .A(n1017), .B(n1397), .Y(n1400) );
  xo2d1_hd U599 ( .A(n1058), .B(n1245), .Y(n1247) );
  xo2d1_hd U600 ( .A(n1016), .B(n1107), .Y(intadd_0_B_14_) );
  xo2d1_hd U601 ( .A(n1015), .B(n1299), .Y(intadd_19_B_2_) );
  xo2d1_hd U602 ( .A(n1013), .B(n1351), .Y(intadd_4_A_13_) );
  xo2d1_hd U603 ( .A(n1869), .B(n1418), .Y(intadd_6_A_10_) );
  xo2d1_hd U604 ( .A(n1017), .B(n1442), .Y(intadd_7_A_10_) );
  xo2d1_hd U605 ( .A(n1891), .B(n1237), .Y(intadd_10_B_6_) );
  xo2d1_hd U606 ( .A(n1059), .B(n1242), .Y(intadd_11_A_2_) );
  xo2d1_hd U607 ( .A(n1016), .B(n1106), .Y(intadd_0_B_13_) );
  xo2d1_hd U608 ( .A(a_m[17]), .B(n1306), .Y(intadd_1_B_5_) );
  xo2d1_hd U609 ( .A(n1014), .B(n1320), .Y(intadd_2_A_13_) );
  xo2d1_hd U610 ( .A(n1891), .B(n1283), .Y(intadd_17_B_0_) );
  xo2d1_hd U611 ( .A(n1017), .B(n1396), .Y(intadd_5_B_12_) );
  xo2d1_hd U612 ( .A(n1016), .B(n1105), .Y(intadd_0_B_12_) );
  xo2d1_hd U613 ( .A(n1869), .B(n1310), .Y(intadd_20_A_0_) );
  xo2d1_hd U614 ( .A(n1013), .B(n1361), .Y(intadd_4_B_12_) );
  xo2d1_hd U615 ( .A(n1059), .B(n1277), .Y(intadd_16_A_0_) );
  xo2d1_hd U616 ( .A(n1015), .B(n1289), .Y(intadd_18_B_0_) );
  xo2d1_hd U617 ( .A(n1014), .B(n1328), .Y(intadd_2_B_12_) );
  xo2d1_hd U618 ( .A(n1891), .B(n1236), .Y(intadd_10_B_4_) );
  xo2d1_hd U619 ( .A(n1869), .B(n1398), .Y(n1399) );
  xo2d1_hd U620 ( .A(n1084), .B(n1815), .Y(N475) );
  xo2d1_hd U621 ( .A(n1016), .B(n1104), .Y(intadd_0_B_11_) );
  xo2d1_hd U622 ( .A(n1014), .B(n1327), .Y(intadd_2_B_11_) );
  xo2d1_hd U623 ( .A(n1059), .B(n1257), .Y(intadd_11_CI) );
  xo2d1_hd U624 ( .A(a_m[17]), .B(n1305), .Y(intadd_1_B_3_) );
  xo2d1_hd U625 ( .A(n1017), .B(n1384), .Y(intadd_5_A_11_) );
  xo2d1_hd U626 ( .A(n1013), .B(n1360), .Y(intadd_4_B_11_) );
  xo2d1_hd U627 ( .A(n1869), .B(n1425), .Y(intadd_6_A_7_) );
  xo2d1_hd U628 ( .A(n1013), .B(n1350), .Y(intadd_4_A_10_) );
  xo2d1_hd U629 ( .A(n1014), .B(n1319), .Y(intadd_2_A_10_) );
  xo2d1_hd U630 ( .A(n1015), .B(n1481), .Y(intadd_8_B_7_) );
  xo2d1_hd U631 ( .A(n1017), .B(n1395), .Y(intadd_5_B_10_) );
  xo2d1_hd U632 ( .A(DP_OP_125J3_130_6300_n2), .B(n1083), .Y(n1084) );
  xo2d1_hd U633 ( .A(n1058), .B(n1258), .Y(intadd_12_A_1_) );
  xo2d1_hd U634 ( .A(n1016), .B(n1102), .Y(intadd_0_B_10_) );
  xo2d1_hd U635 ( .A(n1891), .B(n1298), .Y(intadd_19_B_1_) );
  xo2d1_hd U636 ( .A(n1058), .B(n1263), .Y(intadd_12_CI) );
  xo2d1_hd U637 ( .A(n1016), .B(n1212), .Y(intadd_0_B_9_) );
  xo2d1_hd U638 ( .A(n1013), .B(n1378), .Y(intadd_4_B_9_) );
  xo2d1_hd U639 ( .A(n1017), .B(n1393), .Y(intadd_5_A_9_) );
  xo2d1_hd U640 ( .A(n1891), .B(n1300), .Y(intadd_19_CI) );
  xo2d1_hd U641 ( .A(n1869), .B(n1458), .Y(intadd_7_B_9_) );
  xo2d1_hd U642 ( .A(n1014), .B(n1343), .Y(intadd_2_B_9_) );
  xo2d1_hd U643 ( .A(n1015), .B(n1437), .Y(intadd_6_B_9_) );
  xo2d1_hd U644 ( .A(n1017), .B(n1411), .Y(intadd_5_B_8_) );
  xo2d1_hd U645 ( .A(n1014), .B(n1342), .Y(intadd_2_B_8_) );
  xo2d1_hd U646 ( .A(n1869), .B(n1450), .Y(intadd_7_A_8_) );
  xo2d1_hd U647 ( .A(a_m[20]), .B(n1270), .Y(intadd_14_B_2_) );
  xo2d1_hd U648 ( .A(n1016), .B(n1174), .Y(intadd_0_B_8_) );
  xo2d1_hd U649 ( .A(n1058), .B(n1226), .Y(n1228) );
  xo2d1_hd U650 ( .A(n1015), .B(n1426), .Y(intadd_6_A_8_) );
  xo2d1_hd U651 ( .A(n1017), .B(n1392), .Y(intadd_5_A_7_) );
  xo2d1_hd U652 ( .A(n1015), .B(n1472), .Y(intadd_8_A_4_) );
  xo2d1_hd U653 ( .A(n1059), .B(n1218), .Y(intadd_10_A_3_) );
  xo2d1_hd U654 ( .A(n1869), .B(n1449), .Y(intadd_7_A_7_) );
  xo2d1_hd U655 ( .A(a_m[20]), .B(n1304), .Y(intadd_1_B_2_) );
  xo2d1_hd U656 ( .A(n1014), .B(n1341), .Y(intadd_2_B_7_) );
  xo2d1_hd U657 ( .A(n1016), .B(n1173), .Y(intadd_0_B_7_) );
  xo2d1_hd U658 ( .A(n1869), .B(n1448), .Y(intadd_7_A_6_) );
  xo2d1_hd U659 ( .A(n1014), .B(n1340), .Y(intadd_2_B_6_) );
  xo2d1_hd U660 ( .A(n1059), .B(n1297), .Y(intadd_19_B_0_) );
  xo2d1_hd U661 ( .A(n1015), .B(n1436), .Y(intadd_6_B_6_) );
  xo2d1_hd U662 ( .A(n1891), .B(n1480), .Y(intadd_8_B_6_) );
  xo2d1_hd U663 ( .A(n1017), .B(n1391), .Y(intadd_5_A_6_) );
  xo2d1_hd U664 ( .A(n1016), .B(n1172), .Y(intadd_0_B_6_) );
  xo2d1_hd U665 ( .A(n1014), .B(n1339), .Y(intadd_2_B_5_) );
  xo2d1_hd U666 ( .A(n1869), .B(n1447), .Y(intadd_7_A_5_) );
  xo2d1_hd U667 ( .A(n1017), .B(n1390), .Y(intadd_5_A_5_) );
  xo2d1_hd U668 ( .A(n1015), .B(n1424), .Y(intadd_6_A_5_) );
  xo2d1_hd U669 ( .A(n1059), .B(n1231), .Y(intadd_10_B_1_) );
  xo2d1_hd U670 ( .A(n1891), .B(n1479), .Y(n1851) );
  xo2d1_hd U671 ( .A(n1014), .B(n1338), .Y(intadd_2_B_4_) );
  xo2d1_hd U672 ( .A(a_m[20]), .B(n1922), .Y(n1924) );
  xo2d1_hd U673 ( .A(n1017), .B(n1389), .Y(intadd_5_A_4_) );
  xo2d1_hd U674 ( .A(n1058), .B(n1269), .Y(intadd_14_A_1_) );
  xo2d1_hd U675 ( .A(n1869), .B(n1446), .Y(intadd_7_A_4_) );
  xo2d1_hd U676 ( .A(n1015), .B(n1423), .Y(intadd_6_A_4_) );
  xo2d1_hd U677 ( .A(n1433), .B(n1420), .Y(intadd_6_A_1_) );
  xo2d1_hd U678 ( .A(n1370), .B(n1369), .Y(intadd_4_B_1_) );
  xo2d1_hd U679 ( .A(n1408), .B(n1406), .Y(intadd_5_B_1_) );
  xo2d1_hd U680 ( .A(n1015), .B(n1422), .Y(intadd_6_A_3_) );
  xo2d1_hd U681 ( .A(n1014), .B(n1337), .Y(intadd_2_B_3_) );
  xo2d1_hd U682 ( .A(n1869), .B(n1445), .Y(intadd_7_A_3_) );
  xo2d1_hd U683 ( .A(n1058), .B(n1271), .Y(intadd_14_CI) );
  xo2d1_hd U684 ( .A(n1166), .B(n1090), .Y(intadd_0_A_1_) );
  xo2d1_hd U685 ( .A(n1891), .B(n1477), .Y(intadd_8_B_3_) );
  xo2d1_hd U686 ( .A(n1891), .B(n1471), .Y(intadd_8_A_2_) );
  xo2d1_hd U687 ( .A(n1014), .B(n1336), .Y(intadd_2_B_2_) );
  xo2d1_hd U688 ( .A(n1058), .B(n1309), .Y(intadd_1_CI) );
  xo2d1_hd U689 ( .A(n1869), .B(n1444), .Y(intadd_7_A_2_) );
  xo2d1_hd U690 ( .A(n1454), .B(n1453), .Y(intadd_7_B_1_) );
  xo2d1_hd U691 ( .A(n1335), .B(n1334), .Y(intadd_2_B_1_) );
  xo2d1_hd U692 ( .A(n1015), .B(n1421), .Y(intadd_6_A_2_) );
  xo2d1_hd U693 ( .A(n1891), .B(n1474), .Y(intadd_8_B_1_) );
  xo2d1_hd U694 ( .A(n1014), .B(n1322), .Y(intadd_2_A_1_) );
  scg6d1_hd U695 ( .A(n1553), .B(n1549), .C(n1558), .Y(n1010) );
  xo2d1_hd U696 ( .A(n1439), .B(n1438), .Y(intadd_6_CI) );
  xo2d1_hd U697 ( .A(n1015), .B(n1431), .Y(intadd_6_B_1_) );
  xo2d1_hd U698 ( .A(n1059), .B(n1478), .Y(n1912) );
  xo2d1_hd U699 ( .A(n1891), .B(n1473), .Y(intadd_8_B_0_) );
  xo2d1_hd U700 ( .A(n1485), .B(n1484), .Y(intadd_8_CI) );
  xo2d1_hd U701 ( .A(n1059), .B(n1476), .Y(n1907) );
  xo2d1_hd U702 ( .A(n1058), .B(n1906), .Y(n1917) );
  xo2d1_hd U703 ( .A(n1059), .B(n1466), .Y(n1470) );
  xo2d1_hd U704 ( .A(n1015), .B(n1427), .Y(intadd_6_B_0_) );
  xo2d1_hd U705 ( .A(n1346), .B(n1345), .Y(intadd_2_CI) );
  xo2d1_hd U706 ( .A(n1014), .B(n1326), .Y(intadd_2_B_0_) );
  xo2d1_hd U707 ( .A(a_m[5]), .B(n1167), .Y(n1317) );
  xo2d1_hd U708 ( .A(n1869), .B(n1254), .Y(intadd_11_B_2_) );
  scg2d1_hd U709 ( .A(n1467), .B(n1364), .C(n1022), .D(n1365), .Y(n1089) );
  nid2_hd U710 ( .A(n1930), .Y(n1005) );
  scg2d1_hd U711 ( .A(n1467), .B(n1929), .C(n1022), .D(n1490), .Y(n1325) );
  xo2d1_hd U712 ( .A(n1017), .B(n1260), .Y(intadd_12_B_1_) );
  ao21d1_hd U713 ( .A(n7), .B(n1022), .C(n1007), .Y(n1347) );
  ivd1_hd U714 ( .A(b_m[4]), .Y(n1027) );
  xo2d1_hd U715 ( .A(n1013), .B(n1377), .Y(intadd_4_B_8_) );
  scg2d1_hd U716 ( .A(a_e[6]), .B(n1754), .C(C81_DATA2_6), .D(n1757), .Y(n312)
         );
  xo2d1_hd U717 ( .A(n1013), .B(n1376), .Y(intadd_4_B_7_) );
  xo2d1_hd U718 ( .A(n1013), .B(n1375), .Y(intadd_4_B_6_) );
  scg2d1_hd U719 ( .A(a_e[5]), .B(n1754), .C(C81_DATA2_5), .D(n1757), .Y(n313)
         );
  xo2d1_hd U720 ( .A(n1013), .B(n1374), .Y(intadd_4_B_5_) );
  scg10d1_hd U721 ( .A(n1591), .B(n1551), .C(z[31]), .D(n1010), .Y(n229) );
  scg2d1_hd U722 ( .A(z_m[19]), .B(n1592), .C(n1011), .D(z[19]), .Y(n241) );
  scg2d1_hd U723 ( .A(z_m[18]), .B(n1592), .C(n1011), .D(z[18]), .Y(n242) );
  scg2d1_hd U724 ( .A(z_m[17]), .B(n1592), .C(n1011), .D(z[17]), .Y(n243) );
  scg2d1_hd U725 ( .A(z_m[16]), .B(n1592), .C(n1011), .D(z[16]), .Y(n244) );
  scg2d1_hd U726 ( .A(z_m[15]), .B(n1592), .C(n1011), .D(z[15]), .Y(n245) );
  scg2d1_hd U727 ( .A(z_m[14]), .B(n1592), .C(n1011), .D(z[14]), .Y(n246) );
  scg2d1_hd U728 ( .A(z_m[13]), .B(n1592), .C(n1011), .D(z[13]), .Y(n247) );
  scg2d1_hd U729 ( .A(z_m[12]), .B(n1592), .C(n1011), .D(z[12]), .Y(n248) );
  scg2d1_hd U730 ( .A(z_m[11]), .B(n1592), .C(n1011), .D(z[11]), .Y(n249) );
  scg2d1_hd U731 ( .A(z_m[10]), .B(n1592), .C(n1011), .D(z[10]), .Y(n250) );
  scg2d1_hd U732 ( .A(z_m[9]), .B(n1592), .C(n1011), .D(z[9]), .Y(n251) );
  scg2d1_hd U733 ( .A(a_e[4]), .B(n1754), .C(C81_DATA2_4), .D(n1757), .Y(n314)
         );
  scg2d1_hd U734 ( .A(z_m[21]), .B(n1592), .C(n1011), .D(z[21]), .Y(n239) );
  scg2d1_hd U735 ( .A(z_m[20]), .B(n1592), .C(n1011), .D(z[20]), .Y(n240) );
  xo2d1_hd U736 ( .A(n1016), .B(n1171), .Y(intadd_0_B_5_) );
  scg2d1_hd U737 ( .A(z_m[5]), .B(n1592), .C(n1011), .D(z[5]), .Y(n255) );
  scg2d1_hd U738 ( .A(z_m[6]), .B(n1592), .C(n1011), .D(z[6]), .Y(n254) );
  scg2d1_hd U739 ( .A(z_m[7]), .B(n1592), .C(n1011), .D(z[7]), .Y(n253) );
  scg2d1_hd U740 ( .A(z_m[8]), .B(n1592), .C(n1011), .D(z[8]), .Y(n252) );
  xo2d1_hd U741 ( .A(n1016), .B(n1170), .Y(intadd_0_B_4_) );
  scg9d1_hd U742 ( .A(n1074), .B(n1073), .C(intadd_0_A_0_), .Y(N179) );
  xo2d1_hd U743 ( .A(n1013), .B(n1373), .Y(intadd_4_B_4_) );
  xo2d1_hd U744 ( .A(n1016), .B(n1169), .Y(intadd_0_B_3_) );
  scg2d1_hd U745 ( .A(z_e[8]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n42), .Y(DP_OP_125J3_130_6300_n32) );
  xo2d1_hd U746 ( .A(n1013), .B(n1372), .Y(intadd_4_B_3_) );
  xo2d1_hd U747 ( .A(n1017), .B(n1388), .Y(intadd_5_A_3_) );
  xo2d1_hd U748 ( .A(n1013), .B(n1371), .Y(intadd_4_B_2_) );
  scg2d1_hd U749 ( .A(n1020), .B(b[0]), .C(n7), .D(n1742), .Y(n308) );
  xo2d1_hd U750 ( .A(n1016), .B(n1100), .Y(intadd_0_A_2_) );
  scg9d1_hd U751 ( .A(n1068), .B(n1067), .C(n1069), .Y(N178) );
  scg2d1_hd U752 ( .A(z_e[7]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n41), .Y(DP_OP_125J3_130_6300_n31) );
  xo2d1_hd U753 ( .A(n1017), .B(n1387), .Y(intadd_5_A_2_) );
  scg2d1_hd U754 ( .A(n1020), .B(a[0]), .C(n1829), .D(a_m[0]), .Y(n349) );
  xo2d1_hd U755 ( .A(n1013), .B(n1353), .Y(intadd_4_A_1_) );
  xo2d1_hd U756 ( .A(n1016), .B(n1141), .Y(intadd_0_B_1_) );
  xo2d1_hd U757 ( .A(a_m[11]), .B(n1354), .Y(n1382) );
  scg2d1_hd U758 ( .A(z_e[6]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n40), .Y(DP_OP_125J3_130_6300_n30) );
  xo2d1_hd U759 ( .A(n1017), .B(n1394), .Y(intadd_5_B_0_) );
  xo2d1_hd U760 ( .A(n1017), .B(n1386), .Y(intadd_5_A_1_) );
  xo2d1_hd U761 ( .A(n1869), .B(n1443), .Y(intadd_7_A_1_) );
  or2d1_hd U762 ( .A(n1470), .B(n1469), .Y(n1908) );
  xo2d1_hd U763 ( .A(a_m[8]), .B(n1323), .Y(n1348) );
  xo2d1_hd U764 ( .A(a_m[20]), .B(n1435), .Y(n1462) );
  xo2d1_hd U765 ( .A(n1013), .B(n1359), .Y(intadd_4_B_0_) );
  xo2d1_hd U766 ( .A(a_m[2]), .B(n1072), .Y(n1073) );
  xo2d1_hd U767 ( .A(a_m[2]), .B(n1066), .Y(n1067) );
  xo2d1_hd U768 ( .A(a_m[17]), .B(n1417), .Y(n1455) );
  xo2d1_hd U769 ( .A(n1016), .B(n1101), .Y(intadd_0_B_0_) );
  scg2d1_hd U770 ( .A(n1020), .B(b[29]), .C(b_e[6]), .D(n1850), .Y(n775) );
  scg2d1_hd U771 ( .A(z_e[1]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n35), .Y(DP_OP_125J3_130_6300_n25) );
  xo2d1_hd U772 ( .A(n1869), .B(n1451), .Y(intadd_7_B_0_) );
  scg2d1_hd U773 ( .A(z_e[2]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n36), .Y(DP_OP_125J3_130_6300_n26) );
  xn2d1_hd U774 ( .A(n1064), .B(n1063), .Y(N177) );
  scg2d1_hd U775 ( .A(n1020), .B(a[29]), .C(n1833), .D(a_e[6]), .Y(C1_Z_6) );
  scg2d1_hd U776 ( .A(z_e[3]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n37), .Y(DP_OP_125J3_130_6300_n27) );
  scg2d1_hd U777 ( .A(z_e[4]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n38), .Y(DP_OP_125J3_130_6300_n28) );
  scg2d1_hd U778 ( .A(n1020), .B(b[28]), .C(b_e[5]), .D(n1850), .Y(n774) );
  scg2d1_hd U779 ( .A(z_e[5]), .B(n1844), .C(n1004), .D(
        DP_OP_125J3_130_6300_n39), .Y(DP_OP_125J3_130_6300_n29) );
  xo2d1_hd U780 ( .A(a_m[14]), .B(n1410), .Y(n1440) );
  scg2d1_hd U781 ( .A(n1020), .B(a[28]), .C(n1833), .D(a_e[5]), .Y(C1_Z_5) );
  scg2d1_hd U782 ( .A(n1467), .B(n1887), .C(n1022), .D(n1878), .Y(n1416) );
  nr2d2_hd U783 ( .A(n1312), .B(n1311), .Y(n1933) );
  scg2d1_hd U784 ( .A(n1818), .B(z_m[0]), .C(n2865), .D(round_bit), .Y(n1493)
         );
  scg2d1_hd U785 ( .A(n1467), .B(n1902), .C(n1022), .D(n1905), .Y(n1468) );
  nr2d2_hd U786 ( .A(n1088), .B(n1087), .Y(n1365) );
  nr2d2_hd U787 ( .A(n1291), .B(n1290), .Y(n1866) );
  nr2d2_hd U788 ( .A(n1415), .B(n1234), .Y(n1919) );
  nr2d2_hd U789 ( .A(n1240), .B(n1239), .Y(n1878) );
  scg12d2_hd U790 ( .A(n1290), .B(n1291), .C(n1285), .Y(n1876) );
  ad2d1_hd U791 ( .A(n1112), .B(a_m[23]), .Y(n1077) );
  or2d1_hd U792 ( .A(n1535), .B(n1060), .Y(n1111) );
  xo2d1_hd U793 ( .A(a_m[17]), .B(n1265), .Y(intadd_13_B_1_) );
  xo2d1_hd U794 ( .A(n1891), .B(n1272), .Y(intadd_15_A_2_) );
  or2d1_hd U795 ( .A(n1535), .B(n1548), .Y(n1712) );
  nr2d2_hd U796 ( .A(n1409), .B(n1238), .Y(n1879) );
  or2d1_hd U797 ( .A(n1809), .B(state[1]), .Y(n1497) );
  scg12d2_hd U798 ( .A(n1434), .B(n1216), .C(n1217), .Y(n1904) );
  nr2d2_hd U799 ( .A(n1216), .B(n1434), .Y(n1905) );
  nr2bd2_hd U800 ( .AN(n1517), .B(n1016), .Y(n1207) );
  nr2d2_hd U801 ( .A(a_m[0]), .B(n1804), .Y(n1198) );
  or4d1_hd U802 ( .A(n1771), .B(n1763), .C(n1842), .D(b_e[4]), .Y(n1523) );
  ivd3_hd U803 ( .A(a_m[23]), .Y(n1059) );
  or4d1_hd U804 ( .A(product[3]), .B(product[10]), .C(product[11]), .D(
        product[6]), .Y(n1698) );
  clknd2d1_hd U805 ( .A(n1586), .B(n1566), .Y(n231) );
  clknd2d1_hd U806 ( .A(n1586), .B(n1573), .Y(n233) );
  scg2d1_hd U807 ( .A(b_e[6]), .B(n1768), .C(n1838), .D(C82_DATA2_6), .Y(n321)
         );
  scg2d1_hd U808 ( .A(b_e[5]), .B(n1768), .C(n1838), .D(C82_DATA2_5), .Y(n322)
         );
  scg2d1_hd U809 ( .A(b_e[4]), .B(n1768), .C(n1838), .D(C82_DATA2_4), .Y(n323)
         );
  scg2d1_hd U810 ( .A(b_e[3]), .B(n1768), .C(n1838), .D(C82_DATA2_3), .Y(n324)
         );
  scg2d1_hd U811 ( .A(b_e[2]), .B(n1768), .C(n1838), .D(C82_DATA2_2), .Y(n325)
         );
  nr2ad1_hd U812 ( .A(n1535), .B(n1820), .Y(n2865) );
  oa211d2_hd U813 ( .A(n1719), .B(n1501), .C(n1500), .D(n1111), .Y(n110) );
  scg2d1_hd U814 ( .A(n1467), .B(n1918), .C(n1022), .D(n1921), .Y(n1419) );
  nr2d2_hd U815 ( .A(n1235), .B(n1233), .Y(n1921) );
  nr2d2_hd U816 ( .A(n1061), .B(n1806), .Y(n1209) );
  scg2d1_hd U817 ( .A(z_m[0]), .B(n1592), .C(n1011), .D(z[0]), .Y(n260) );
  scg2d1_hd U818 ( .A(z_m[1]), .B(n1592), .C(n1011), .D(z[1]), .Y(n259) );
  scg2d1_hd U819 ( .A(z_m[2]), .B(n1592), .C(n1011), .D(z[2]), .Y(n258) );
  scg2d1_hd U820 ( .A(z_m[3]), .B(n1592), .C(n1011), .D(z[3]), .Y(n257) );
  scg2d1_hd U821 ( .A(z_m[4]), .B(n1592), .C(n1011), .D(z[4]), .Y(n256) );
  nr2d4_hd U822 ( .A(n1589), .B(n1588), .Y(n1592) );
  oa21d2_hd U823 ( .A(n1754), .B(n1810), .C(n1118), .Y(n1757) );
  scg2d1_hd U824 ( .A(n1757), .B(n1755), .C(a_e[0]), .D(n1754), .Y(n318) );
  scg2d1_hd U825 ( .A(a_e[2]), .B(n1754), .C(C81_DATA2_2), .D(n1757), .Y(n316)
         );
  scg2d1_hd U826 ( .A(a_e[3]), .B(n1754), .C(C81_DATA2_3), .D(n1757), .Y(n315)
         );
  ao21d2_hd U827 ( .A(n1836), .B(n1745), .C(n1783), .Y(n1754) );
  nr2ad1_hd U828 ( .A(n1707), .B(n1815), .Y(n1713) );
  scg2d1_hd U829 ( .A(n1020), .B(b[24]), .C(b_e[1]), .D(n1850), .Y(n770) );
  scg2d1_hd U830 ( .A(n1020), .B(b[23]), .C(b_e[0]), .D(n1850), .Y(n769) );
  scg2d1_hd U831 ( .A(n1019), .B(b[25]), .C(b_e[2]), .D(n1850), .Y(n771) );
  scg2d1_hd U832 ( .A(n1019), .B(b[26]), .C(b_e[3]), .D(n1850), .Y(n772) );
  scg2d1_hd U833 ( .A(n1019), .B(b[27]), .C(b_e[4]), .D(n1850), .Y(n773) );
  nr2ad1_hd U834 ( .A(n1535), .B(n1812), .Y(n1850) );
  scg2d1_hd U835 ( .A(n1020), .B(a[24]), .C(n1833), .D(a_e[1]), .Y(C1_Z_1) );
  scg2d1_hd U836 ( .A(n1019), .B(a[25]), .C(n1833), .D(a_e[2]), .Y(C1_Z_2) );
  scg2d1_hd U837 ( .A(n1019), .B(a[26]), .C(n1833), .D(a_e[3]), .Y(C1_Z_3) );
  scg2d1_hd U838 ( .A(n1019), .B(a[27]), .C(n1833), .D(a_e[4]), .Y(C1_Z_4) );
  nr2ad1_hd U839 ( .A(n1820), .B(n1807), .Y(n1833) );
  nr2ad1_hd U840 ( .A(n1593), .B(n105), .Y(n1707) );
  ao21d2_hd U841 ( .A(n1055), .B(n1116), .C(n1057), .Y(n1928) );
  nid2_hd U842 ( .A(b_m[5]), .Y(n1028) );
  xo3d1_hd U843 ( .A(n1079), .B(intadd_1_n1), .C(n1078), .Y(N223) );
  scg4d1_hd U844 ( .A(n1052), .B(n1905), .C(n1050), .D(n1903), .E(n1048), .F(
        n1904), .G(n1902), .H(intadd_3_SUM_17_), .Y(n1276) );
  scg14d1_hd U845 ( .A(n1054), .B(n1904), .C(n1858), .Y(n1859) );
  scg17d1_hd U846 ( .A(n1819), .B(n1818), .C(n2017), .D(n1828), .Y(n1845) );
  ad3d1_hd U847 ( .A(n1808), .B(o_AB_ACK), .C(i_AB_STB), .Y(n2017) );
  nid2_hd U848 ( .A(n359), .Y(n1021) );
  ivd1_hd U849 ( .A(n1850), .Y(n1765) );
  ivd1_hd U850 ( .A(n1713), .Y(n1710) );
  ivd1_hd U851 ( .A(n1711), .Y(n1686) );
  ivd1_hd U852 ( .A(n1677), .Y(n1594) );
  ivd1_hd U853 ( .A(n2865), .Y(n1815) );
  ivd1_hd U854 ( .A(n1821), .Y(n1535) );
  ivd1_hd U855 ( .A(n1874), .Y(n2029) );
  nid2_hd U856 ( .A(n1913), .Y(n1016) );
  ivd1_hd U857 ( .A(n1886), .Y(n2027) );
  ivd1_hd U858 ( .A(intadd_11_n1), .Y(n1182) );
  nid2_hd U859 ( .A(n1938), .Y(n1017) );
  ivd1_hd U860 ( .A(n1233), .Y(n1415) );
  nid2_hd U861 ( .A(n1881), .Y(n1015) );
  ivd1_hd U862 ( .A(n1864), .Y(n2031) );
  ivd1_hd U863 ( .A(n1057), .Y(n1056) );
  clknd2d2_hd U864 ( .A(n1850), .B(n1720), .Y(n1744) );
  ivd2_hd U865 ( .A(n1783), .Y(n1829) );
  ivd2_hd U866 ( .A(n1118), .Y(n1019) );
  ivd1_hd U867 ( .A(n1558), .Y(n1588) );
  ivd2_hd U868 ( .A(n1010), .Y(n1011) );
  nr2d1_hd U869 ( .A(n1809), .B(n1548), .Y(n1558) );
  ivd1_hd U870 ( .A(n1833), .Y(n1810) );
  ivd1_hd U871 ( .A(n1754), .Y(n1762) );
  clknd2d2_hd U872 ( .A(n1833), .B(n1059), .Y(n1832) );
  ao21d1_hd U873 ( .A(n1118), .B(n1765), .C(n1768), .Y(n1838) );
  ivd1_hd U874 ( .A(n1768), .Y(n1843) );
  ao21d1_hd U875 ( .A(n1747), .B(n1745), .C(n1720), .Y(n1768) );
  oa21d1_hd U876 ( .A(n1765), .B(b_m[23]), .C(n1118), .Y(n1720) );
  nr2d1_hd U877 ( .A(n1549), .B(n1546), .Y(n1745) );
  ivd1_hd U878 ( .A(n1553), .Y(n1546) );
  nr2d1_hd U879 ( .A(n1548), .B(n1807), .Y(n1553) );
  nd3d1_hd U880 ( .A(n1552), .B(n1540), .C(n1538), .Y(n1549) );
  nr2d1_hd U881 ( .A(n1505), .B(n1504), .Y(n1836) );
  nr2d1_hd U882 ( .A(n1523), .B(n1522), .Y(n1747) );
  ivd2_hd U883 ( .A(n1704), .Y(n1705) );
  ivd2_hd U884 ( .A(n1712), .Y(n1012) );
  nr2ad1_hd U885 ( .A(n1707), .B(n1594), .Y(n1711) );
  nr2bd1_hd U886 ( .AN(n1818), .B(n1819), .Y(n1699) );
  nr2d1_hd U887 ( .A(n1497), .B(n1534), .Y(n1677) );
  ivd1_hd U888 ( .A(n1604), .Y(n1603) );
  ivd1_hd U889 ( .A(n1613), .Y(n1612) );
  ivd1_hd U890 ( .A(n1622), .Y(n1621) );
  ivd1_hd U891 ( .A(n1631), .Y(n1630) );
  ivd1_hd U892 ( .A(n1640), .Y(n1639) );
  ivd1_hd U893 ( .A(state[2]), .Y(n1822) );
  nid2_hd U894 ( .A(n1797), .Y(n1014) );
  ad2d2_hd U895 ( .A(n1095), .B(n1168), .Y(n1490) );
  ivd1_hd U896 ( .A(n1324), .Y(n1311) );
  ivd1_hd U897 ( .A(intadd_17_SUM_2_), .Y(n1179) );
  ivd1_hd U898 ( .A(n1882), .Y(n2028) );
  ivd1_hd U899 ( .A(n1355), .Y(n1290) );
  nid2_hd U900 ( .A(b_m[6]), .Y(n1029) );
  ivd1_hd U901 ( .A(a_m[8]), .Y(n1791) );
  ivd1_hd U902 ( .A(intadd_16_SUM_2_), .Y(n1177) );
  ivd1_hd U903 ( .A(n1895), .Y(n2025) );
  ivd1_hd U904 ( .A(intadd_11_SUM_5_), .Y(n1183) );
  nid2_hd U905 ( .A(b_m[9]), .Y(n1034) );
  nid2_hd U906 ( .A(b_m[11]), .Y(n1037) );
  ivd1_hd U907 ( .A(n1898), .Y(n2024) );
  ivd1_hd U908 ( .A(a_m[18]), .Y(n1775) );
  ivd1_hd U909 ( .A(a_m[19]), .Y(n1773) );
  ivd1_hd U910 ( .A(intadd_15_n1), .Y(n1184) );
  nid2_hd U911 ( .A(b_m[18]), .Y(n1047) );
  ivd1_hd U912 ( .A(n1860), .Y(n2032) );
  ivd1_hd U913 ( .A(n1303), .Y(n1076) );
  ivd2_hd U914 ( .A(n1720), .Y(n1742) );
  ivd1_hd U915 ( .A(n1745), .Y(n1835) );
  scg17d1_hd U916 ( .A(z_m[10]), .B(n1713), .C(n1647), .D(n1646), .Y(n272) );
  scg17d1_hd U917 ( .A(z_m[2]), .B(n1713), .C(n1684), .D(n1683), .Y(n280) );
  scg17d1_hd U918 ( .A(z_m[6]), .B(n1713), .C(n1665), .D(n1664), .Y(n276) );
  ivd1_hd U919 ( .A(n1580), .Y(n1587) );
  ao21d1_hd U920 ( .A(n1560), .B(n1559), .C(n1588), .Y(n1580) );
  ao22d1_hd U921 ( .A(n1554), .B(n1553), .C(n1589), .D(n1558), .Y(n1586) );
  scg20d1_hd U922 ( .A(z_e[7]), .B(z_e[8]), .C(z_e[9]), .Y(n1589) );
  scg17d1_hd U923 ( .A(z_m[14]), .B(n1713), .C(n1629), .D(n1628), .Y(n268) );
  scg2d1_hd U924 ( .A(state[0]), .B(n1828), .C(n1827), .D(n1826), .Y(n353) );
  nr2d1_hd U925 ( .A(n1809), .B(n1820), .Y(n359) );
  scg17d1_hd U926 ( .A(z_m[18]), .B(n1713), .C(n1611), .D(n1610), .Y(n264) );
  ivd1_hd U927 ( .A(n1838), .Y(n1770) );
  ivd1_hd U928 ( .A(state[3]), .Y(n1846) );
  ivd1_hd U929 ( .A(b_e[8]), .Y(n1763) );
  ivd1_hd U930 ( .A(b_e[0]), .Y(n1771) );
  scg17d1_hd U931 ( .A(z_m[20]), .B(n1713), .C(n1602), .D(n1601), .Y(n262) );
  ivd1_hd U932 ( .A(z_m[23]), .Y(n1814) );
  ivd1_hd U933 ( .A(state[0]), .Y(n1534) );
  ivd1_hd U934 ( .A(a_e[9]), .Y(n1761) );
  ivd1_hd U935 ( .A(b_e[9]), .Y(n1842) );
  ivd1_hd U936 ( .A(state[1]), .Y(n1824) );
  nr2d1_hd U937 ( .A(n1822), .B(state[3]), .Y(n1821) );
  ivd1_hd U938 ( .A(a_m[0]), .Y(n1806) );
  ivd1_hd U939 ( .A(a_m[1]), .Y(n1804) );
  ivd1_hd U940 ( .A(a_m[3]), .Y(n1801) );
  ivd1_hd U941 ( .A(a_m[4]), .Y(n1799) );
  ivd1_hd U942 ( .A(n1467), .Y(n1404) );
  ivd1_hd U943 ( .A(a_m[7]), .Y(n1793) );
  ivd1_hd U944 ( .A(n1096), .Y(n1168) );
  ivd1_hd U945 ( .A(a_m[6]), .Y(n1795) );
  ivd1_hd U946 ( .A(a_m[5]), .Y(n1797) );
  fad1_hd U947 ( .A(n1873), .B(n1872), .CI(n1871), .CO(n1874), .S(n1870) );
  ivd1_hd U948 ( .A(a_m[10]), .Y(n1787) );
  ivd1_hd U949 ( .A(a_m[9]), .Y(n1789) );
  ivd1_hd U950 ( .A(a_m[2]), .Y(n1913) );
  fad1_hd U951 ( .A(n1885), .B(n1884), .CI(n1883), .CO(n1886), .S(n1882) );
  ivd1_hd U952 ( .A(a_m[13]), .Y(n1782) );
  ivd1_hd U953 ( .A(a_m[12]), .Y(n1784) );
  ivd1_hd U954 ( .A(a_m[15]), .Y(n1779) );
  ivd1_hd U955 ( .A(a_m[16]), .Y(n1777) );
  fad1_hd U956 ( .A(intadd_15_SUM_1_), .B(n1900), .CI(n1899), .CO(n1901), .S(
        n1898) );
  fad1_hd U957 ( .A(n1863), .B(n1862), .CI(n1861), .CO(n1864), .S(n1860) );
  ivd1_hd U958 ( .A(a_m[21]), .Y(n1831) );
  ivd2_hd U959 ( .A(n1118), .Y(n1020) );
  nr2d1_hd U960 ( .A(n1497), .B(state[0]), .Y(n1818) );
  nr2d1_hd U961 ( .A(n1806), .B(n1009), .Y(N176) );
  ivd2_hd U962 ( .A(n1488), .Y(n1363) );
  ivd2_hd U963 ( .A(n1356), .Y(n1934) );
  ivd2_hd U964 ( .A(n1402), .Y(n1867) );
  ivd2_hd U965 ( .A(n1281), .Y(n1888) );
  ad3d2_hd U966 ( .A(n1235), .B(n1234), .C(n1233), .Y(n1920) );
  nr2d1_hd U967 ( .A(n1807), .B(n1812), .Y(n1808) );
  ad2d2_hd U968 ( .A(n1240), .B(n1409), .Y(n1887) );
  oa21d1_hd U969 ( .A(n1009), .B(n1022), .C(n1070), .Y(n1467) );
  ao22d1_hd U970 ( .A(a_m[2]), .B(a_m[1]), .C(n1804), .D(n1913), .Y(n1061) );
  ao22d1_hd U971 ( .A(n7), .B(n1198), .C(n1022), .D(n1209), .Y(n1062) );
  oa21d1_hd U972 ( .A(n1404), .B(n1158), .C(n1062), .Y(n1064) );
  nr3d1_hd U973 ( .A(N176), .B(n1064), .C(n1016), .Y(n1068) );
  nr2d1_hd U974 ( .A(a_m[0]), .B(a_m[1]), .Y(n1517) );
  ivd1_hd U975 ( .A(n1070), .Y(n1065) );
  ao22d1_hd U976 ( .A(n1007), .B(n1065), .C(n1070), .D(n1024), .Y(n1465) );
  scg4d1_hd U977 ( .A(n7), .B(n1207), .C(n1022), .D(n1198), .E(n1465), .F(
        n1175), .G(n1209), .H(n1007), .Y(n1066) );
  nr2d1_hd U978 ( .A(a_m[3]), .B(a_m[2]), .Y(n1512) );
  ao21d1_hd U979 ( .A(a_m[2]), .B(a_m[3]), .C(n1512), .Y(n1086) );
  oa211d1_hd U980 ( .A(n1023), .B(n1024), .C(n1525), .D(n1070), .Y(n1071) );
  scg4d1_hd U981 ( .A(n1025), .B(n1209), .C(n1022), .D(n1207), .E(n1198), .F(
        n1007), .G(n1475), .H(n1175), .Y(n1072) );
  oa22d1_hd U982 ( .A(n1891), .B(n1831), .C(a_m[21]), .D(a_m[20]), .Y(n1434)
         );
  nr2d1_hd U983 ( .A(a_m[21]), .B(a_m[22]), .Y(n1511) );
  ao21d1_hd U984 ( .A(a_m[22]), .B(a_m[21]), .C(n1511), .Y(n1217) );
  ao22d1_hd U985 ( .A(b_m[23]), .B(n1904), .C(n1902), .D(n1928), .Y(n1303) );
  oa22d1_hd U986 ( .A(n1077), .B(n1076), .C(n1059), .D(n1075), .Y(n1079) );
  nr2d1_hd U987 ( .A(n1059), .B(n1053), .Y(n1862) );
  oa22ad1_hd U988 ( .A(n1059), .B(n1526), .C(n1056), .D(n1862), .Y(n1078) );
  ao22d1_hd U989 ( .A(a_e[9]), .B(b_e[9]), .C(n1842), .D(n1761), .Y(n1081) );
  nr2d1_hd U990 ( .A(DP_OP_125J3_130_6300_n12), .B(n1081), .Y(n1080) );
  ao211d1_hd U991 ( .A(DP_OP_125J3_130_6300_n12), .B(n1081), .C(n1111), .D(
        n1080), .Y(n1082) );
  ao21d1_hd U992 ( .A(z_e[9]), .B(n1844), .C(n1082), .Y(n1083) );
  ivd1_hd U993 ( .A(n1086), .Y(n1087) );
  oa22d1_hd U994 ( .A(n1799), .B(n1801), .C(a_m[3]), .D(a_m[4]), .Y(n1085) );
  nr2d1_hd U995 ( .A(a_m[5]), .B(a_m[4]), .Y(n1513) );
  ao21d1_hd U996 ( .A(a_m[4]), .B(a_m[5]), .C(n1513), .Y(n1088) );
  nd3d1_hd U997 ( .A(n1087), .B(n1085), .C(n1088), .Y(n1488) );
  scg4d1_hd U998 ( .A(n7), .B(n1363), .C(n1022), .D(n1366), .E(n1465), .F(
        n1364), .G(n1007), .H(n1365), .Y(n1166) );
  ao21d1_hd U999 ( .A(n7), .B(n1366), .C(n1089), .Y(n1215) );
  nd3d1_hd U1000 ( .A(n1215), .B(a_m[5]), .C(n1213), .Y(n1165) );
  oa211d1_hd U1001 ( .A(n1052), .B(intadd_3_n1), .C(n1054), .D(n1057), .Y(
        n1091) );
  ao22d1_hd U1002 ( .A(n1056), .B(n1366), .C(n1364), .D(n1857), .Y(n1092) );
  oa21d1_hd U1003 ( .A(n1488), .B(n1055), .C(n1092), .Y(n1093) );
  oa22d1_hd U1004 ( .A(n1791), .B(n1793), .C(a_m[7]), .D(a_m[8]), .Y(n1095) );
  oa22d1_hd U1005 ( .A(n1797), .B(n1795), .C(a_m[6]), .D(a_m[5]), .Y(n1096) );
  nr2d1_hd U1006 ( .A(a_m[7]), .B(a_m[6]), .Y(n1514) );
  ao21d1_hd U1007 ( .A(a_m[6]), .B(a_m[7]), .C(n1514), .Y(n1094) );
  nr3d1_hd U1008 ( .A(n1168), .B(n1094), .C(n1095), .Y(n1930) );
  scg4d1_hd U1009 ( .A(n1052), .B(n1490), .C(n1050), .D(n1491), .E(n1048), .F(
        n1005), .G(n1929), .H(intadd_3_SUM_17_), .Y(n1097) );
  fad1_hd U1010 ( .A(intadd_5_SUM_14_), .B(n1099), .CI(n1098), .CO(
        intadd_0_A_24_), .S(intadd_0_A_23_) );
  scg4d1_hd U1011 ( .A(n1028), .B(n1198), .C(n1029), .D(n1209), .E(n1207), .F(
        n1006), .G(n1175), .H(intadd_3_SUM_2_), .Y(n1100) );
  scg4d1_hd U1012 ( .A(n1006), .B(n1209), .C(n1007), .D(n1207), .E(n1198), .F(
        n1025), .G(n1175), .H(intadd_3_SUM_0_), .Y(n1101) );
  scg4d1_hd U1013 ( .A(n1041), .B(n1209), .C(n1038), .D(n1207), .E(n1198), .F(
        n1039), .G(n1175), .H(intadd_3_SUM_10_), .Y(n1102) );
  scg4d1_hd U1014 ( .A(n1042), .B(n1209), .C(n1039), .D(n1207), .E(n1198), .F(
        n1041), .G(n1175), .H(intadd_3_SUM_11_), .Y(n1104) );
  scg4d1_hd U1015 ( .A(n1008), .B(n1209), .C(n1041), .D(n1207), .E(n1198), .F(
        n1042), .G(n1175), .H(intadd_3_SUM_12_), .Y(n1105) );
  scg4d1_hd U1016 ( .A(n1045), .B(n1209), .C(n1042), .D(n1207), .E(n1198), .F(
        n1008), .G(n1175), .H(intadd_3_SUM_13_), .Y(n1106) );
  scg4d1_hd U1017 ( .A(n1045), .B(n1198), .C(n1047), .D(n1209), .E(n1207), .F(
        n1008), .G(n1175), .H(intadd_3_SUM_14_), .Y(n1107) );
  scg4d1_hd U1018 ( .A(n1045), .B(n1207), .C(n1047), .D(n1198), .E(n1048), .F(
        n1209), .G(n1175), .H(intadd_3_SUM_15_), .Y(n1108) );
  scg4d1_hd U1019 ( .A(n1048), .B(n1198), .C(n1047), .D(n1207), .E(n1050), .F(
        n1209), .G(n1175), .H(intadd_3_SUM_16_), .Y(n1109) );
  scg4d1_hd U1020 ( .A(n1052), .B(n1209), .C(n1050), .D(n1198), .E(n1207), .F(
        n1048), .G(n1175), .H(intadd_3_SUM_17_), .Y(n1110) );
  scg4d1_hd U1021 ( .A(n1936), .B(n1175), .C(n1052), .D(n1198), .E(n1209), .F(
        n1054), .G(n1207), .H(n1050), .Y(n1114) );
  oa21d1_hd U1022 ( .A(intadd_3_n1), .B(n1052), .C(n1054), .Y(n1115) );
  scg4d1_hd U1023 ( .A(n1054), .B(n1198), .C(n1056), .D(n1209), .E(n1207), .F(
        n1052), .G(n1175), .H(n1429), .Y(n1136) );
  scg4d1_hd U1024 ( .A(n1028), .B(n1209), .C(n1025), .D(n1207), .E(n1198), .F(
        n1006), .G(n1175), .H(intadd_3_SUM_1_), .Y(n1141) );
  ao21d1_hd U1025 ( .A(n1517), .B(n1054), .C(n1016), .Y(n1154) );
  mx2id1_hd U1026 ( .D0(n1154), .D1(n1016), .S(n1150), .YN(intadd_0_B_20_) );
  ao22d1_hd U1027 ( .A(n1056), .B(n1207), .C(n1175), .D(n1928), .Y(n1164) );
  ivd1_hd U1028 ( .A(n1928), .Y(n1486) );
  nr2d1_hd U1029 ( .A(n1158), .B(n1486), .Y(n1162) );
  ao22d1_hd U1030 ( .A(a_m[2]), .B(n1164), .C(n1162), .D(n1016), .Y(
        intadd_0_B_21_) );
  nr2d1_hd U1031 ( .A(n1166), .B(n1165), .Y(n1318) );
  scg4d1_hd U1032 ( .A(n1025), .B(n1365), .C(n1022), .D(n1363), .E(n1366), .F(
        n1007), .G(n1475), .H(n1364), .Y(n1167) );
  xo3d1_hd U1033 ( .A(n1318), .B(n1317), .C(n1344), .Y(intadd_0_B_2_) );
  scg4d1_hd U1034 ( .A(n1028), .B(n1207), .C(n1029), .D(n1198), .E(n1030), .F(
        n1209), .G(n1175), .H(intadd_3_SUM_3_), .Y(n1169) );
  scg4d1_hd U1035 ( .A(n1032), .B(n1209), .C(n1029), .D(n1207), .E(n1198), .F(
        n1030), .G(n1175), .H(intadd_3_SUM_4_), .Y(n1170) );
  scg4d1_hd U1036 ( .A(n1032), .B(n1198), .C(n1034), .D(n1209), .E(n1207), .F(
        n1030), .G(n1175), .H(intadd_3_SUM_5_), .Y(n1171) );
  scg4d1_hd U1037 ( .A(n1032), .B(n1207), .C(n1035), .D(n1209), .E(n1034), .F(
        n1198), .G(n1175), .H(intadd_3_SUM_6_), .Y(n1172) );
  scg4d1_hd U1038 ( .A(n1037), .B(n1209), .C(n1035), .D(n1198), .E(n1207), .F(
        n1034), .G(n1175), .H(intadd_3_SUM_7_), .Y(n1173) );
  scg4d1_hd U1039 ( .A(n1038), .B(n1209), .C(n1035), .D(n1207), .E(n1198), .F(
        n1037), .G(n1175), .H(intadd_3_SUM_8_), .Y(n1174) );
  scg4d1_hd U1040 ( .A(n1039), .B(n1209), .C(n1037), .D(n1207), .E(n1198), .F(
        n1038), .G(n1175), .H(intadd_3_SUM_9_), .Y(n1212) );
  nr2d1_hd U1041 ( .A(n1014), .B(n1213), .Y(n1214) );
  nr2d1_hd U1042 ( .A(n1059), .B(n1031), .Y(intadd_10_A_2_) );
  scg4d1_hd U1043 ( .A(n1037), .B(n1905), .C(n1035), .D(n1903), .E(n1034), .F(
        n1904), .G(n1902), .H(intadd_3_SUM_7_), .Y(n1218) );
  ao21d1_hd U1044 ( .A(a_m[8]), .B(n1223), .C(n1219), .Y(n1229) );
  scg4d1_hd U1045 ( .A(n1038), .B(n1905), .C(n1035), .D(n1904), .E(n1903), .F(
        b_m[11]), .G(n1902), .H(intadd_3_SUM_8_), .Y(n1226) );
  ivd1_hd U1046 ( .A(n1227), .Y(intadd_10_A_4_) );
  fad1_hd U1047 ( .A(n2034), .B(n1229), .CI(n1228), .CO(n1230), .S(n1227) );
  ivd1_hd U1048 ( .A(n1230), .Y(intadd_10_A_5_) );
  scg4d1_hd U1049 ( .A(n1032), .B(n1903), .C(n1034), .D(n1905), .E(n1030), .F(
        n1904), .G(n1902), .H(intadd_3_SUM_5_), .Y(n1231) );
  oa211d1_hd U1050 ( .A(n1033), .B(n1031), .C(n1058), .D(n1524), .Y(n1232) );
  oa22d1_hd U1051 ( .A(n1773), .B(a_m[20]), .C(n1891), .D(a_m[19]), .Y(n1235)
         );
  oa22d1_hd U1052 ( .A(n1881), .B(n1775), .C(a_m[18]), .D(a_m[17]), .Y(n1233)
         );
  oa22d1_hd U1053 ( .A(n1773), .B(n1775), .C(a_m[18]), .D(a_m[19]), .Y(n1234)
         );
  scg4d1_hd U1054 ( .A(n1042), .B(n1921), .C(n1039), .D(n1920), .E(n1041), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_11_), .Y(n1236) );
  scg4d1_hd U1055 ( .A(n1045), .B(n1921), .C(n1042), .D(n1920), .E(n1008), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_13_), .Y(n1237) );
  oa22d1_hd U1056 ( .A(n1777), .B(a_m[17]), .C(n1881), .D(a_m[16]), .Y(n1240)
         );
  nr2d1_hd U1057 ( .A(a_m[15]), .B(a_m[14]), .Y(n1515) );
  ao21d1_hd U1058 ( .A(a_m[14]), .B(a_m[15]), .C(n1515), .Y(n1409) );
  ivd1_hd U1059 ( .A(n1409), .Y(n1239) );
  oa22d1_hd U1060 ( .A(n1777), .B(n1779), .C(a_m[15]), .D(a_m[16]), .Y(n1238)
         );
  nd3d1_hd U1061 ( .A(n1239), .B(n1238), .C(n1240), .Y(n1281) );
  scg4d1_hd U1062 ( .A(n1052), .B(n1878), .C(n1050), .D(n1879), .E(n1888), .F(
        n1048), .G(n1887), .H(intadd_3_SUM_17_), .Y(n1241) );
  nr2d1_hd U1063 ( .A(n1059), .B(n1040), .Y(intadd_11_A_1_) );
  scg4d1_hd U1064 ( .A(n1045), .B(n1905), .C(n1042), .D(n1904), .E(n1903), .F(
        n1008), .G(n1902), .H(intadd_3_SUM_13_), .Y(n1242) );
  nr2d1_hd U1065 ( .A(n1059), .B(n1043), .Y(n1274) );
  ivd1_hd U1066 ( .A(n1274), .Y(intadd_13_A_0_) );
  nr2d1_hd U1067 ( .A(n1041), .B(n1039), .Y(n1243) );
  nr2d1_hd U1068 ( .A(n1243), .B(n1059), .Y(n1252) );
  ivd1_hd U1069 ( .A(n1252), .Y(n1244) );
  ao21d1_hd U1070 ( .A(a_m[14]), .B(n1253), .C(n1244), .Y(n1248) );
  scg4d1_hd U1071 ( .A(n1045), .B(n1903), .C(n1047), .D(n1905), .E(n1008), .F(
        n1904), .G(n1902), .H(intadd_3_SUM_14_), .Y(n1245) );
  ivd1_hd U1072 ( .A(n1246), .Y(intadd_11_A_3_) );
  fad1_hd U1073 ( .A(intadd_13_A_0_), .B(n1248), .CI(n1247), .CO(n1249), .S(
        n1246) );
  ivd1_hd U1074 ( .A(n1249), .Y(intadd_11_A_4_) );
  ivd1_hd U1075 ( .A(n2034), .Y(n1251) );
  nr2d1_hd U1076 ( .A(a_m[11]), .B(n1259), .Y(n1250) );
  oa22d1_hd U1077 ( .A(n1037), .B(n1017), .C(n1251), .D(n1250), .Y(
        intadd_11_B_0_) );
  scg4d1_hd U1078 ( .A(n1052), .B(n1921), .C(n1050), .D(n1919), .E(n1048), .F(
        n1920), .G(n1918), .H(intadd_3_SUM_17_), .Y(n1255) );
  scg4d1_hd U1079 ( .A(n1054), .B(n1919), .C(n1056), .D(n1921), .E(n1918), .F(
        n1429), .G(n1052), .H(n1920), .Y(n1256) );
  scg4d1_hd U1080 ( .A(n1042), .B(n1905), .C(n1039), .D(n1904), .E(n1903), .F(
        n1041), .G(n1902), .H(intadd_3_SUM_11_), .Y(n1257) );
  scg4d1_hd U1081 ( .A(n1041), .B(n1905), .C(n1038), .D(n1904), .E(n1903), .F(
        n1039), .G(n1902), .H(intadd_3_SUM_10_), .Y(n1258) );
  nr2d1_hd U1082 ( .A(n1059), .B(n1036), .Y(intadd_12_B_0_) );
  oa22d1_hd U1083 ( .A(n1034), .B(n1259), .C(n1037), .D(n2034), .Y(n1260) );
  scg4d1_hd U1084 ( .A(n1045), .B(n1919), .C(n1047), .D(n1921), .E(n1918), .F(
        intadd_3_SUM_14_), .G(n1008), .H(n1920), .Y(n1261) );
  scg4d1_hd U1085 ( .A(n1054), .B(n1879), .C(n1056), .D(n1878), .E(n1888), .F(
        n1052), .G(n1887), .H(n1429), .Y(n1262) );
  scg4d1_hd U1086 ( .A(n1039), .B(n1905), .C(b_m[11]), .D(n1904), .E(n1903), 
        .F(n1038), .G(n1902), .H(intadd_3_SUM_9_), .Y(n1263) );
  scg4d1_hd U1087 ( .A(n1048), .B(n1903), .C(n1047), .D(n1904), .E(n1050), .F(
        n1905), .G(n1902), .H(intadd_3_SUM_16_), .Y(n1264) );
  nr2d1_hd U1088 ( .A(n1059), .B(n1044), .Y(intadd_13_B_0_) );
  oa211d1_hd U1089 ( .A(n1046), .B(n1043), .C(n1058), .D(n1532), .Y(n1265) );
  ao22d1_hd U1090 ( .A(n1054), .B(n1920), .C(n1918), .D(n1857), .Y(n1266) );
  scg14d1_hd U1091 ( .A(n1056), .B(n1919), .C(n1266), .Y(n1267) );
  scg4d1_hd U1092 ( .A(n1045), .B(n1904), .C(n1047), .D(n1903), .E(n1905), .F(
        n1048), .G(n1902), .H(intadd_3_SUM_15_), .Y(n1268) );
  scg4d1_hd U1093 ( .A(n1032), .B(n1905), .C(n1029), .D(n1904), .E(n1903), .F(
        n1030), .G(n1902), .H(intadd_3_SUM_4_), .Y(n1269) );
  nr2d1_hd U1094 ( .A(n1059), .B(n1027), .Y(intadd_14_B_0_) );
  scg4d1_hd U1095 ( .A(n1038), .B(n1921), .C(n1035), .D(n1920), .E(n1037), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_8_), .Y(n1270) );
  scg4d1_hd U1096 ( .A(n1028), .B(n1904), .C(n1029), .D(n1903), .E(n1905), .F(
        n1030), .G(n1902), .H(intadd_3_SUM_3_), .Y(n1271) );
  nr2d1_hd U1097 ( .A(n1059), .B(n1049), .Y(intadd_15_A_1_) );
  oa211d1_hd U1098 ( .A(n1049), .B(n1051), .C(n1058), .D(n1855), .Y(n1272) );
  nr3d1_hd U1099 ( .A(a_m[17]), .B(n1059), .C(n1046), .Y(n1273) );
  oa22d1_hd U1100 ( .A(n1045), .B(n1015), .C(n1274), .D(n1273), .Y(
        intadd_15_B_0_) );
  scg4d1_hd U1101 ( .A(n1054), .B(n1903), .C(n1056), .D(n1905), .E(n1052), .F(
        n1904), .G(n1902), .H(n1429), .Y(n1275) );
  scg4d1_hd U1102 ( .A(n1008), .B(n1905), .C(n1041), .D(n1904), .E(n1903), .F(
        n1042), .G(n1902), .H(intadd_3_SUM_12_), .Y(n1277) );
  scg4d1_hd U1103 ( .A(n1045), .B(n1920), .C(n1047), .D(n1919), .E(n1921), .F(
        n1048), .G(n1918), .H(intadd_3_SUM_15_), .Y(n1278) );
  scg4d1_hd U1104 ( .A(n1048), .B(n1919), .C(n1047), .D(n1920), .E(n1921), .F(
        n1050), .G(n1918), .H(intadd_3_SUM_16_), .Y(n1279) );
  ao22d1_hd U1105 ( .A(b_m[23]), .B(n1879), .C(n1887), .D(n1857), .Y(n1280) );
  oa21d1_hd U1106 ( .A(n1281), .B(n1055), .C(n1280), .Y(n1282) );
  scg4d1_hd U1107 ( .A(n1008), .B(n1921), .C(n1041), .D(n1920), .E(n1042), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_12_), .Y(n1283) );
  scg4d1_hd U1108 ( .A(n1048), .B(n1879), .C(n1047), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_16_), .G(n1050), .H(n1878), .Y(n1284) );
  oa22d1_hd U1109 ( .A(n1938), .B(a_m[12]), .C(n1784), .D(a_m[11]), .Y(n1355)
         );
  nr2d1_hd U1110 ( .A(a_m[13]), .B(a_m[12]), .Y(n1516) );
  ao21d1_hd U1111 ( .A(a_m[12]), .B(a_m[13]), .C(n1516), .Y(n1285) );
  oa22d1_hd U1112 ( .A(n1782), .B(a_m[14]), .C(n1869), .D(a_m[13]), .Y(n1291)
         );
  ao22d1_hd U1113 ( .A(n1054), .B(n1876), .C(n1875), .D(n1857), .Y(n1286) );
  oa21d1_hd U1114 ( .A(n1057), .B(n1402), .C(n1286), .Y(n1287) );
  scg4d1_hd U1115 ( .A(n1045), .B(n1888), .C(n1047), .D(n1879), .E(n1048), .F(
        n1878), .G(n1887), .H(intadd_3_SUM_15_), .Y(n1288) );
  scg4d1_hd U1116 ( .A(n1008), .B(n1878), .C(n1041), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_12_), .G(n1879), .H(n1042), .Y(n1289) );
  scg4d1_hd U1117 ( .A(n1048), .B(n1867), .C(n1047), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_16_), .G(n1866), .H(n1050), .Y(n1292) );
  oa22d1_hd U1118 ( .A(n1013), .B(a_m[9]), .C(n1789), .D(a_m[8]), .Y(n1324) );
  nr2d1_hd U1119 ( .A(a_m[9]), .B(a_m[10]), .Y(n1510) );
  ao21d1_hd U1120 ( .A(a_m[10]), .B(a_m[9]), .C(n1510), .Y(n1293) );
  ao22d1_hd U1121 ( .A(a_m[11]), .B(a_m[10]), .C(n1787), .D(n1938), .Y(n1312)
         );
  ao22d1_hd U1122 ( .A(n1054), .B(n1932), .C(n1935), .D(n1857), .Y(n1294) );
  oa21d1_hd U1123 ( .A(n1057), .B(n1356), .C(n1294), .Y(n1295) );
  scg4d1_hd U1124 ( .A(n1045), .B(n1876), .C(n1047), .D(n1867), .E(n1875), .F(
        intadd_3_SUM_15_), .G(n1048), .H(n1866), .Y(n1296) );
  scg4d1_hd U1125 ( .A(n1032), .B(n1904), .C(n1035), .D(n1905), .E(n1903), .F(
        n1034), .G(n1902), .H(intadd_3_SUM_6_), .Y(n1297) );
  scg4d1_hd U1126 ( .A(n1041), .B(n1921), .C(n1038), .D(n1920), .E(n1039), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_10_), .Y(n1298) );
  scg4d1_hd U1127 ( .A(n1045), .B(n1879), .C(n1047), .D(n1878), .E(n1888), .F(
        n1008), .G(n1887), .H(intadd_3_SUM_14_), .Y(n1299) );
  scg4d1_hd U1128 ( .A(n1039), .B(n1921), .C(n1037), .D(n1920), .E(n1038), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_9_), .Y(n1300) );
  nr2d1_hd U1129 ( .A(n1059), .B(n1026), .Y(intadd_1_B_0_) );
  nr2d1_hd U1130 ( .A(n1059), .B(n1301), .Y(n1302) );
  scg4d1_hd U1131 ( .A(n1037), .B(n1921), .C(n1035), .D(n1919), .E(n1034), .F(
        n1920), .G(n1918), .H(intadd_3_SUM_7_), .Y(n1304) );
  scg4d1_hd U1132 ( .A(n1042), .B(n1878), .C(n1039), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_11_), .G(n1879), .H(n1041), .Y(n1305) );
  scg4d1_hd U1133 ( .A(n1045), .B(n1878), .C(n1042), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_13_), .G(n1879), .H(n1008), .Y(n1306) );
  scg4d1_hd U1134 ( .A(n1052), .B(n1866), .C(n1050), .D(n1867), .E(n1875), .F(
        intadd_3_SUM_17_), .G(n1876), .H(n1048), .Y(n1307) );
  scg4d1_hd U1135 ( .A(n1054), .B(n1867), .C(n1056), .D(n1866), .E(n1875), .F(
        n1429), .G(n1876), .H(n1052), .Y(n1308) );
  scg4d1_hd U1136 ( .A(n1028), .B(n1903), .C(n1029), .D(n1905), .E(n1006), .F(
        n1904), .G(n1902), .H(intadd_3_SUM_2_), .Y(n1309) );
  scg4d1_hd U1137 ( .A(n1008), .B(n1866), .C(n1041), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_12_), .G(n1042), .H(n1867), .Y(n1310) );
  scg4d1_hd U1138 ( .A(n1048), .B(n1934), .C(n1047), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_16_), .G(n1933), .H(n1050), .Y(n1313) );
  ao22d1_hd U1139 ( .A(b_m[23]), .B(n1491), .C(n1929), .D(n1857), .Y(n1314) );
  scg14d1_hd U1140 ( .A(n1005), .B(n1054), .C(n1314), .Y(n1315) );
  scg4d1_hd U1141 ( .A(n1045), .B(n1932), .C(n1047), .D(n1934), .E(n1935), .F(
        intadd_3_SUM_15_), .G(n1048), .H(n1933), .Y(n1316) );
  scg16d1_hd U1142 ( .A(n1344), .B(n1318), .C(n1317), .Y(intadd_2_A_0_) );
  scg4d1_hd U1143 ( .A(n1041), .B(n1365), .C(n1038), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_10_), .G(n1039), .H(n1366), .Y(n1319) );
  scg4d1_hd U1144 ( .A(n1045), .B(n1365), .C(n1042), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_13_), .G(n1008), .H(n1366), .Y(n1320) );
  scg4d1_hd U1145 ( .A(n1936), .B(n1364), .C(n1052), .D(n1366), .E(n1365), .F(
        n1054), .G(n1363), .H(n1050), .Y(n1321) );
  scg4d1_hd U1146 ( .A(n1028), .B(n1365), .C(n1025), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_1_), .G(n1006), .H(n1366), .Y(n1322) );
  scg4d1_hd U1147 ( .A(n1025), .B(n1490), .C(n1022), .D(n1005), .E(n1475), .F(
        n1929), .G(n1491), .H(n1007), .Y(n1323) );
  scg4d1_hd U1148 ( .A(n7), .B(n1005), .C(n1022), .D(n1491), .E(n1007), .F(
        n1490), .G(n1465), .H(n1929), .Y(n1335) );
  ao21d1_hd U1149 ( .A(n7), .B(n1491), .C(n1325), .Y(n1346) );
  nd3d1_hd U1150 ( .A(a_m[8]), .B(n1346), .C(n1344), .Y(n1333) );
  nr2d1_hd U1151 ( .A(n1335), .B(n1333), .Y(n1349) );
  xo3d1_hd U1152 ( .A(n1348), .B(n1379), .C(n1349), .Y(intadd_2_A_2_) );
  scg4d1_hd U1153 ( .A(n1006), .B(n1365), .C(n1007), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_0_), .G(n1025), .H(n1366), .Y(n1326) );
  scg4d1_hd U1154 ( .A(n1042), .B(n1365), .C(n1039), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_11_), .G(n1041), .H(n1366), .Y(n1327) );
  scg4d1_hd U1155 ( .A(n1008), .B(n1365), .C(n1041), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_12_), .G(n1042), .H(n1366), .Y(n1328) );
  scg4d1_hd U1156 ( .A(n1045), .B(n1366), .C(n1047), .D(n1365), .E(n1364), .F(
        intadd_3_SUM_14_), .G(n1008), .H(n1363), .Y(n1329) );
  scg4d1_hd U1157 ( .A(n1045), .B(n1363), .C(n1047), .D(n1366), .E(n1364), .F(
        intadd_3_SUM_15_), .G(n1365), .H(n1048), .Y(n1330) );
  scg4d1_hd U1158 ( .A(n1048), .B(n1366), .C(n1047), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_16_), .G(n1365), .H(n1050), .Y(n1331) );
  scg4d1_hd U1159 ( .A(n1052), .B(n1365), .C(n1050), .D(n1366), .E(n1364), .F(
        intadd_3_SUM_17_), .G(n1048), .H(n1363), .Y(n1332) );
  scg4d1_hd U1160 ( .A(n1028), .B(n1366), .C(n1029), .D(n1365), .E(n1364), .F(
        intadd_3_SUM_2_), .G(n1006), .H(n1363), .Y(n1336) );
  scg4d1_hd U1161 ( .A(n1028), .B(n1363), .C(n1029), .D(n1366), .E(n1364), .F(
        intadd_3_SUM_3_), .G(n1365), .H(n1030), .Y(n1337) );
  scg4d1_hd U1162 ( .A(n1032), .B(n1365), .C(n1029), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_4_), .G(n1030), .H(n1366), .Y(n1338) );
  scg4d1_hd U1163 ( .A(n1032), .B(n1366), .C(n1034), .D(n1365), .E(n1364), .F(
        intadd_3_SUM_5_), .G(n1030), .H(n1363), .Y(n1339) );
  scg4d1_hd U1164 ( .A(n1032), .B(n1363), .C(n1035), .D(n1365), .E(n1364), .F(
        intadd_3_SUM_6_), .G(n1366), .H(n1034), .Y(n1340) );
  scg4d1_hd U1165 ( .A(n1037), .B(n1365), .C(n1035), .D(n1366), .E(n1364), .F(
        intadd_3_SUM_7_), .G(n1034), .H(n1363), .Y(n1341) );
  scg4d1_hd U1166 ( .A(n1038), .B(n1365), .C(n1035), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_8_), .G(n1037), .H(n1366), .Y(n1342) );
  scg4d1_hd U1167 ( .A(n1039), .B(n1365), .C(n1037), .D(n1363), .E(n1364), .F(
        intadd_3_SUM_9_), .G(n1038), .H(n1366), .Y(n1343) );
  nr2d1_hd U1168 ( .A(n1013), .B(n1344), .Y(n1345) );
  oa22d1_hd U1169 ( .A(n1347), .B(n1026), .C(n1024), .D(n1023), .Y(intadd_3_CI) );
  scg16d1_hd U1170 ( .A(n1379), .B(n1349), .C(n1348), .Y(intadd_4_A_0_) );
  scg4d1_hd U1171 ( .A(n1041), .B(n1490), .C(n1038), .D(n1005), .E(n1039), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_10_), .Y(n1350) );
  scg4d1_hd U1172 ( .A(n1045), .B(n1490), .C(n1042), .D(n1005), .E(n1008), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_13_), .Y(n1351) );
  scg4d1_hd U1173 ( .A(n1045), .B(n1005), .C(n1047), .D(n1491), .E(n1490), .F(
        n1048), .G(n1929), .H(intadd_3_SUM_15_), .Y(n1352) );
  scg4d1_hd U1174 ( .A(n1028), .B(n1490), .C(n1025), .D(n1005), .E(n1006), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_1_), .Y(n1353) );
  scg4d1_hd U1175 ( .A(n1025), .B(n1933), .C(n1022), .D(n1932), .E(n1007), .F(
        n1934), .G(n1935), .H(n1475), .Y(n1354) );
  scg4d1_hd U1176 ( .A(n7), .B(n1932), .C(n1022), .D(n1934), .E(n1933), .F(
        n1007), .G(n1465), .H(n1935), .Y(n1370) );
  oa22d1_hd U1177 ( .A(n1404), .B(n1357), .C(n1009), .D(n1356), .Y(n1358) );
  ao21d1_hd U1178 ( .A(n1022), .B(n1933), .C(n1358), .Y(n1381) );
  nd3d1_hd U1179 ( .A(a_m[11]), .B(n1381), .C(n1379), .Y(n1368) );
  nr2d1_hd U1180 ( .A(n1370), .B(n1368), .Y(n1383) );
  xo3d1_hd U1181 ( .A(n1382), .B(n1412), .C(n1383), .Y(intadd_4_A_2_) );
  scg4d1_hd U1182 ( .A(n1006), .B(n1490), .C(n1007), .D(n1005), .E(n1025), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_0_), .Y(n1359) );
  scg4d1_hd U1183 ( .A(n1042), .B(n1490), .C(n1039), .D(n1005), .E(n1041), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_11_), .Y(n1360) );
  scg4d1_hd U1184 ( .A(n1008), .B(n1490), .C(n1041), .D(n1005), .E(n1042), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_12_), .Y(n1361) );
  scg4d1_hd U1185 ( .A(n1045), .B(n1491), .C(n1047), .D(n1490), .E(n1005), .F(
        n1008), .G(n1929), .H(intadd_3_SUM_14_), .Y(n1362) );
  scg4d1_hd U1186 ( .A(n1054), .B(n1366), .C(n1056), .D(n1365), .E(n1364), .F(
        n1429), .G(n1052), .H(n1363), .Y(n1367) );
  scg4d1_hd U1187 ( .A(n1028), .B(n1491), .C(n1029), .D(n1490), .E(n1005), .F(
        n1006), .G(n1929), .H(intadd_3_SUM_2_), .Y(n1371) );
  scg4d1_hd U1188 ( .A(n1028), .B(n1005), .C(n1029), .D(n1491), .E(n1490), .F(
        n1030), .G(n1929), .H(intadd_3_SUM_3_), .Y(n1372) );
  scg4d1_hd U1189 ( .A(n1032), .B(n1490), .C(n1029), .D(n1005), .E(n1030), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_4_), .Y(n1373) );
  scg4d1_hd U1190 ( .A(n1032), .B(n1491), .C(n1034), .D(n1490), .E(n1005), .F(
        n1030), .G(n1929), .H(intadd_3_SUM_5_), .Y(n1374) );
  scg4d1_hd U1191 ( .A(n1032), .B(n1005), .C(n1035), .D(n1490), .E(n1034), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_6_), .Y(n1375) );
  scg4d1_hd U1192 ( .A(n1037), .B(n1490), .C(n1035), .D(n1491), .E(n1034), .F(
        n1005), .G(n1929), .H(intadd_3_SUM_7_), .Y(n1376) );
  scg4d1_hd U1193 ( .A(n1038), .B(n1490), .C(n1035), .D(n1005), .E(n1037), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_8_), .Y(n1377) );
  scg4d1_hd U1194 ( .A(n1039), .B(n1490), .C(n1037), .D(n1005), .E(n1038), .F(
        n1491), .G(n1929), .H(intadd_3_SUM_9_), .Y(n1378) );
  nr2d1_hd U1195 ( .A(n1017), .B(n1379), .Y(n1380) );
  scg16d1_hd U1196 ( .A(n1412), .B(n1383), .C(n1382), .Y(intadd_5_A_0_) );
  scg4d1_hd U1197 ( .A(n1042), .B(n1933), .C(n1039), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_11_), .G(n1041), .H(n1934), .Y(n1384) );
  scg4d1_hd U1198 ( .A(n1048), .B(n1491), .C(n1047), .D(n1005), .E(n1490), .F(
        n1050), .G(n1929), .H(intadd_3_SUM_16_), .Y(n1385) );
  scg4d1_hd U1199 ( .A(n1028), .B(n1933), .C(n1025), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_1_), .G(n1006), .H(n1934), .Y(n1386) );
  scg4d1_hd U1200 ( .A(n1028), .B(n1934), .C(n1029), .D(n1933), .E(n1935), .F(
        intadd_3_SUM_2_), .G(n1932), .H(n1006), .Y(n1387) );
  scg4d1_hd U1201 ( .A(n1028), .B(n1932), .C(n1029), .D(n1934), .E(n1935), .F(
        intadd_3_SUM_3_), .G(n1030), .H(n1933), .Y(n1388) );
  scg4d1_hd U1202 ( .A(n1032), .B(n1933), .C(n1029), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_4_), .G(n1030), .H(n1934), .Y(n1389) );
  scg4d1_hd U1203 ( .A(n1032), .B(n1934), .C(n1034), .D(n1933), .E(n1935), .F(
        intadd_3_SUM_5_), .G(n1932), .H(n1030), .Y(n1390) );
  scg4d1_hd U1204 ( .A(n1032), .B(n1932), .C(n1035), .D(n1933), .E(n1935), .F(
        intadd_3_SUM_6_), .G(n1034), .H(n1934), .Y(n1391) );
  scg4d1_hd U1205 ( .A(n1037), .B(n1933), .C(n1035), .D(n1934), .E(n1935), .F(
        intadd_3_SUM_7_), .G(n1932), .H(n1034), .Y(n1392) );
  scg4d1_hd U1206 ( .A(n1039), .B(n1933), .C(n1037), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_9_), .G(n1038), .H(n1934), .Y(n1393) );
  scg4d1_hd U1207 ( .A(n1006), .B(n1933), .C(n1007), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_0_), .G(n1025), .H(n1934), .Y(n1394) );
  scg4d1_hd U1208 ( .A(n1041), .B(n1933), .C(n1038), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_10_), .G(n1039), .H(n1934), .Y(n1395) );
  scg4d1_hd U1209 ( .A(n1008), .B(n1933), .C(n1041), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_12_), .G(n1042), .H(n1934), .Y(n1396) );
  scg4d1_hd U1210 ( .A(n1045), .B(n1934), .C(n1047), .D(n1933), .E(n1935), .F(
        intadd_3_SUM_14_), .G(n1932), .H(n1008), .Y(n1397) );
  scg4d1_hd U1211 ( .A(n1042), .B(n1866), .C(n1039), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_11_), .G(n1041), .H(n1867), .Y(n1398) );
  fad1_hd U1212 ( .A(intadd_6_SUM_8_), .B(n1400), .CI(n1399), .CO(
        intadd_5_B_15_), .S(intadd_5_B_14_) );
  scg4d1_hd U1213 ( .A(n1054), .B(n1491), .C(n1056), .D(n1490), .E(n1005), .F(
        n1052), .G(n1929), .H(n1429), .Y(n1401) );
  scg4d1_hd U1214 ( .A(n7), .B(n1876), .C(n1022), .D(n1867), .E(n1866), .F(
        n1007), .G(n1465), .H(n1875), .Y(n1408) );
  oa22d1_hd U1215 ( .A(n1404), .B(n1403), .C(n1009), .D(n1402), .Y(n1405) );
  ao21d1_hd U1216 ( .A(n1022), .B(n1866), .C(n1405), .Y(n1414) );
  nd3d1_hd U1217 ( .A(a_m[14]), .B(n1414), .C(n1412), .Y(n1407) );
  nr2d1_hd U1218 ( .A(n1408), .B(n1407), .Y(n1441) );
  scg4d1_hd U1219 ( .A(n1025), .B(n1866), .C(n1022), .D(n1876), .E(n1007), .F(
        n1867), .G(n1875), .H(n1475), .Y(n1410) );
  xo3d1_hd U1220 ( .A(n1441), .B(n1459), .C(n1440), .Y(intadd_5_B_2_) );
  scg4d1_hd U1221 ( .A(n1038), .B(n1933), .C(n1035), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_8_), .G(n1037), .H(n1934), .Y(n1411) );
  nr2d1_hd U1222 ( .A(n1869), .B(n1412), .Y(n1413) );
  scg4d1_hd U1223 ( .A(n7), .B(n1888), .C(n1022), .D(n1879), .E(n1887), .F(
        n1465), .G(n1878), .H(n1007), .Y(n1454) );
  ao21d1_hd U1224 ( .A(n7), .B(n1879), .C(n1416), .Y(n1461) );
  nd3d1_hd U1225 ( .A(a_m[17]), .B(n1461), .C(n1459), .Y(n1452) );
  nr2d1_hd U1226 ( .A(n1454), .B(n1452), .Y(n1457) );
  scg4d1_hd U1227 ( .A(n1025), .B(n1878), .C(n1022), .D(n1888), .E(n1887), .F(
        n1475), .G(n1007), .H(n1879), .Y(n1417) );
  scg16d1_hd U1228 ( .A(n1456), .B(n1457), .C(n1455), .Y(intadd_6_A_0_) );
  scg4d1_hd U1229 ( .A(n1045), .B(n1866), .C(n1042), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_13_), .G(n1008), .H(n1867), .Y(n1418) );
  scg4d1_hd U1230 ( .A(n7), .B(n1920), .C(n1022), .D(n1919), .E(n1918), .F(
        n1465), .G(n1007), .H(n1921), .Y(n1433) );
  ao21d1_hd U1231 ( .A(n7), .B(n1919), .C(n1419), .Y(n1439) );
  nd3d1_hd U1232 ( .A(a_m[20]), .B(n1439), .C(n1456), .Y(n1432) );
  scg4d1_hd U1233 ( .A(n1028), .B(n1879), .C(n1029), .D(n1878), .E(n1888), .F(
        n1006), .G(n1887), .H(intadd_3_SUM_2_), .Y(n1421) );
  scg4d1_hd U1234 ( .A(n1028), .B(n1888), .C(n1029), .D(n1879), .E(n1030), .F(
        n1878), .G(n1887), .H(intadd_3_SUM_3_), .Y(n1422) );
  scg4d1_hd U1235 ( .A(n1032), .B(n1878), .C(n1029), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_4_), .G(n1879), .H(n1030), .Y(n1423) );
  scg4d1_hd U1236 ( .A(n1032), .B(n1879), .C(n1034), .D(n1878), .E(n1888), .F(
        n1030), .G(n1887), .H(intadd_3_SUM_5_), .Y(n1424) );
  scg4d1_hd U1237 ( .A(n1041), .B(n1866), .C(n1038), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_10_), .G(n1039), .H(n1867), .Y(n1425) );
  scg4d1_hd U1238 ( .A(n1038), .B(n1878), .C(n1035), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_8_), .G(n1879), .H(n1037), .Y(n1426) );
  scg4d1_hd U1239 ( .A(n1006), .B(n1878), .C(n1007), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_0_), .G(n1879), .H(n1025), .Y(n1427) );
  scg4d1_hd U1240 ( .A(n1052), .B(n1933), .C(n1050), .D(n1934), .E(n1935), .F(
        intadd_3_SUM_17_), .G(n1932), .H(n1048), .Y(n1428) );
  scg4d1_hd U1241 ( .A(n1054), .B(n1934), .C(n1056), .D(n1933), .E(n1935), .F(
        n1429), .G(n1932), .H(n1052), .Y(n1430) );
  scg4d1_hd U1242 ( .A(n1028), .B(n1878), .C(n1025), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_1_), .G(n1879), .H(n1006), .Y(n1431) );
  nr2d1_hd U1243 ( .A(n1433), .B(n1432), .Y(n1463) );
  nr2d1_hd U1244 ( .A(n1009), .B(n1434), .Y(n1464) );
  ivd1_hd U1245 ( .A(n1464), .Y(n1483) );
  scg4d1_hd U1246 ( .A(n1025), .B(n1921), .C(n1022), .D(n1920), .E(n1918), .F(
        n1475), .G(n1007), .H(n1919), .Y(n1435) );
  xo3d1_hd U1247 ( .A(n1463), .B(n1483), .C(n1462), .Y(intadd_6_B_2_) );
  scg4d1_hd U1248 ( .A(n1032), .B(n1888), .C(n1035), .D(n1878), .E(n1034), .F(
        n1879), .G(n1887), .H(intadd_3_SUM_6_), .Y(n1436) );
  scg4d1_hd U1249 ( .A(n1039), .B(n1878), .C(n1037), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_9_), .G(n1879), .H(n1038), .Y(n1437) );
  nr2d1_hd U1250 ( .A(n1891), .B(n1456), .Y(n1438) );
  scg16d1_hd U1251 ( .A(n1459), .B(n1441), .C(n1440), .Y(intadd_7_A_0_) );
  scg4d1_hd U1252 ( .A(n1045), .B(n1933), .C(n1042), .D(n1932), .E(n1935), .F(
        intadd_3_SUM_13_), .G(n1008), .H(n1934), .Y(n1442) );
  scg4d1_hd U1253 ( .A(n1028), .B(n1866), .C(n1025), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_1_), .G(n1006), .H(n1867), .Y(n1443) );
  scg4d1_hd U1254 ( .A(n1028), .B(n1867), .C(n1029), .D(n1866), .E(n1875), .F(
        intadd_3_SUM_2_), .G(n1876), .H(n1006), .Y(n1444) );
  scg4d1_hd U1255 ( .A(n1028), .B(n1876), .C(n1029), .D(n1867), .E(n1875), .F(
        intadd_3_SUM_3_), .G(n1030), .H(n1866), .Y(n1445) );
  scg4d1_hd U1256 ( .A(n1032), .B(n1866), .C(n1029), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_4_), .G(n1030), .H(n1867), .Y(n1446) );
  scg4d1_hd U1257 ( .A(n1032), .B(n1867), .C(n1034), .D(n1866), .E(n1875), .F(
        intadd_3_SUM_5_), .G(n1876), .H(n1030), .Y(n1447) );
  scg4d1_hd U1258 ( .A(n1032), .B(n1876), .C(n1035), .D(n1866), .E(n1875), .F(
        intadd_3_SUM_6_), .G(n1034), .H(n1867), .Y(n1448) );
  scg4d1_hd U1259 ( .A(n1037), .B(n1866), .C(n1035), .D(n1867), .E(n1875), .F(
        intadd_3_SUM_7_), .G(n1876), .H(n1034), .Y(n1449) );
  scg4d1_hd U1260 ( .A(n1038), .B(n1866), .C(n1035), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_8_), .G(n1037), .H(n1867), .Y(n1450) );
  scg4d1_hd U1261 ( .A(n1006), .B(n1866), .C(n1007), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_0_), .G(n1025), .H(n1867), .Y(n1451) );
  xo3d1_hd U1262 ( .A(n1457), .B(n1456), .C(n1455), .Y(intadd_7_B_2_) );
  scg4d1_hd U1263 ( .A(n1039), .B(n1866), .C(n1037), .D(n1876), .E(n1875), .F(
        intadd_3_SUM_9_), .G(n1038), .H(n1867), .Y(n1458) );
  nr2d1_hd U1264 ( .A(n1015), .B(n1459), .Y(n1460) );
  oa21d1_hd U1265 ( .A(n1464), .B(n1463), .C(n1462), .Y(intadd_8_A_0_) );
  scg4d1_hd U1266 ( .A(n7), .B(n1904), .C(n1022), .D(n1903), .E(n1905), .F(
        n1007), .G(n1465), .H(n1902), .Y(n1466) );
  ao21d1_hd U1267 ( .A(n7), .B(n1903), .C(n1468), .Y(n1485) );
  nd3d1_hd U1268 ( .A(n1058), .B(n1485), .C(n1483), .Y(n1469) );
  scg14d1_hd U1269 ( .A(n1470), .B(n1469), .C(n1908), .Y(intadd_8_A_1_) );
  scg4d1_hd U1270 ( .A(n1028), .B(n1919), .C(n1029), .D(n1921), .E(n1918), .F(
        intadd_3_SUM_2_), .G(n1006), .H(n1920), .Y(n1471) );
  scg4d1_hd U1271 ( .A(n1037), .B(n1878), .C(n1035), .D(n1879), .E(n1888), .F(
        n1034), .G(n1887), .H(intadd_3_SUM_7_), .Y(n1472) );
  scg4d1_hd U1272 ( .A(n1006), .B(n1921), .C(n1007), .D(n1920), .E(n1025), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_0_), .Y(n1473) );
  scg4d1_hd U1273 ( .A(n1028), .B(n1921), .C(n1025), .D(n1920), .E(n1006), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_1_), .Y(n1474) );
  scg4d1_hd U1274 ( .A(n1025), .B(n1905), .C(n1022), .D(n1904), .E(n1903), .F(
        n1007), .G(n1902), .H(n1475), .Y(n1476) );
  xo3d1_hd U1275 ( .A(n1908), .B(n1909), .C(n1907), .Y(intadd_8_B_2_) );
  scg4d1_hd U1276 ( .A(n1028), .B(n1920), .C(n1029), .D(n1919), .E(n1921), .F(
        n1030), .G(n1918), .H(intadd_3_SUM_3_), .Y(n1477) );
  ivd1_hd U1277 ( .A(intadd_1_SUM_0_), .Y(n1853) );
  scg4d1_hd U1278 ( .A(n1028), .B(n1905), .C(n1025), .D(n1904), .E(n1903), .F(
        n1006), .G(n1902), .H(intadd_3_SUM_1_), .Y(n1478) );
  scg4d1_hd U1279 ( .A(n1032), .B(n1919), .C(n1034), .D(n1921), .E(n1918), .F(
        intadd_3_SUM_5_), .G(n1030), .H(n1920), .Y(n1479) );
  scg4d1_hd U1280 ( .A(n1032), .B(n1920), .C(n1035), .D(n1921), .E(n1918), .F(
        intadd_3_SUM_6_), .G(n1919), .H(n1034), .Y(n1480) );
  scg4d1_hd U1281 ( .A(n1041), .B(n1878), .C(n1038), .D(n1888), .E(n1887), .F(
        intadd_3_SUM_10_), .G(n1879), .H(n1039), .Y(n1481) );
  scg4d1_hd U1282 ( .A(n1045), .B(n1867), .C(n1047), .D(n1866), .E(n1875), .F(
        intadd_3_SUM_14_), .G(n1876), .H(n1008), .Y(n1482) );
  nr2d1_hd U1283 ( .A(n1059), .B(n1483), .Y(n1484) );
  oa22d1_hd U1284 ( .A(n1057), .B(n1488), .C(n1487), .D(n1486), .Y(n1489) );
  scg4d1_hd U1285 ( .A(n1936), .B(n1929), .C(n1052), .D(n1491), .E(n1490), .F(
        n1054), .G(n1005), .H(n1050), .Y(n1492) );
  ao21d1_hd U1286 ( .A(n1012), .B(product[25]), .C(n1493), .Y(n104) );
  nr2d1_hd U1287 ( .A(z_e[4]), .B(z_e[3]), .Y(n1495) );
  nr2d1_hd U1288 ( .A(z_e[6]), .B(z_e[5]), .Y(n1494) );
  nr3d1_hd U1289 ( .A(z_e[2]), .B(z_e[1]), .C(n1556), .Y(n1496) );
  oa21d1_hd U1290 ( .A(n1496), .B(n1555), .C(z_e[9]), .Y(n1819) );
  ao21d1_hd U1291 ( .A(n2865), .B(n1814), .C(n1699), .Y(n1500) );
  nd3d1_hd U1292 ( .A(z_m[0]), .B(z_m[1]), .C(z_m[2]), .Y(n1676) );
  ivd1_hd U1293 ( .A(n1676), .Y(n1675) );
  nd3d1_hd U1294 ( .A(n1675), .B(z_m[3]), .C(z_m[4]), .Y(n1667) );
  ivd1_hd U1295 ( .A(n1667), .Y(n1666) );
  nd3d1_hd U1296 ( .A(n1666), .B(z_m[5]), .C(z_m[6]), .Y(n1658) );
  ivd1_hd U1297 ( .A(n1658), .Y(n1657) );
  nd3d1_hd U1298 ( .A(n1657), .B(z_m[7]), .C(z_m[8]), .Y(n1649) );
  ivd1_hd U1299 ( .A(n1649), .Y(n1648) );
  nd3d1_hd U1300 ( .A(n1648), .B(z_m[9]), .C(z_m[10]), .Y(n1640) );
  nd3d1_hd U1301 ( .A(n1639), .B(z_m[11]), .C(z_m[12]), .Y(n1631) );
  nd3d1_hd U1302 ( .A(n1630), .B(z_m[13]), .C(z_m[14]), .Y(n1622) );
  nd3d1_hd U1303 ( .A(n1621), .B(z_m[15]), .C(z_m[16]), .Y(n1613) );
  nd3d1_hd U1304 ( .A(n1612), .B(z_m[17]), .C(z_m[18]), .Y(n1604) );
  nd3d1_hd U1305 ( .A(n1603), .B(z_m[19]), .C(z_m[20]), .Y(n1597) );
  ivd1_hd U1306 ( .A(n1597), .Y(n1595) );
  nd3d1_hd U1307 ( .A(z_m[22]), .B(z_m[21]), .C(n1595), .Y(n1719) );
  nr2d1_hd U1308 ( .A(round_bit), .B(sticky), .Y(n1499) );
  ivd1_hd U1309 ( .A(z_m[0]), .Y(n1498) );
  ao211d1_hd U1310 ( .A(n1499), .B(n1498), .C(net922), .D(n1594), .Y(n1593) );
  nr4d1_hd U1311 ( .A(a_e[4]), .B(n10), .C(a_e[6]), .D(a_e[1]), .Y(n1502) );
  scg13d1_hd U1312 ( .A(a_e[3]), .B(a_e[2]), .C(n1502), .Y(n1505) );
  ivd1_hd U1313 ( .A(a_e[5]), .Y(n1503) );
  nd4d1_hd U1314 ( .A(a_e[9]), .B(a_e[8]), .C(a_e[0]), .D(n1503), .Y(n1504) );
  nd2bd1_hd U1315 ( .AN(n1505), .B(n1761), .Y(n1506) );
  nr4d1_hd U1316 ( .A(a_e[8]), .B(a_e[5]), .C(a_e[0]), .D(n1506), .Y(n1545) );
  nr4d1_hd U1317 ( .A(b_e[5]), .B(b_e[2]), .C(b_e[1]), .D(n14), .Y(n1508) );
  nr2d1_hd U1318 ( .A(b_e[6]), .B(b_e[3]), .Y(n1507) );
  nr4d1_hd U1319 ( .A(b_e[4]), .B(b_e[0]), .C(n1522), .D(n1509), .Y(n1543) );
  nr2d1_hd U1320 ( .A(n1545), .B(n1543), .Y(n1552) );
  nd4d1_hd U1321 ( .A(n1059), .B(n1017), .C(n1777), .D(n1773), .Y(n1521) );
  nd4d1_hd U1322 ( .A(n1015), .B(n1775), .C(n1013), .D(n1891), .Y(n1520) );
  nd4d1_hd U1323 ( .A(n1513), .B(n1512), .C(n1511), .D(n1510), .Y(n1519) );
  nd4d1_hd U1324 ( .A(n1517), .B(n1516), .C(n1515), .D(n1514), .Y(n1518) );
  nr4d1_hd U1325 ( .A(n1521), .B(n1520), .C(n1519), .D(n1518), .Y(n1539) );
  nr4d1_hd U1326 ( .A(n1054), .B(n1006), .C(n1025), .D(n7), .Y(n1530) );
  nr4d1_hd U1327 ( .A(n1526), .B(n1855), .C(n1525), .D(n1524), .Y(n1529) );
  nr4d1_hd U1328 ( .A(n1029), .B(n1037), .C(n1034), .D(n1035), .Y(n1528) );
  nr4d1_hd U1329 ( .A(n1041), .B(n1039), .C(n1047), .D(n1038), .Y(n1527) );
  nd4d1_hd U1330 ( .A(n1530), .B(n1529), .C(n1528), .D(n1527), .Y(n1531) );
  nr4d1_hd U1331 ( .A(n1008), .B(n1028), .C(n1532), .D(n1531), .Y(n1541) );
  nr2d1_hd U1332 ( .A(n1810), .B(n10), .Y(n1750) );
  ivd1_hd U1333 ( .A(n1750), .Y(n1748) );
  ivd1_hd U1334 ( .A(DP_OP_113J3_124_6892_n3), .Y(n1749) );
  ao22d1_hd U1335 ( .A(DP_OP_113J3_124_6892_n3), .B(n1748), .C(n1750), .D(
        n1749), .Y(n1533) );
  ao22d1_hd U1336 ( .A(n1754), .B(a_e[7]), .C(n1757), .D(n1533), .Y(n141) );
  oa22ad1_hd U1337 ( .A(n1765), .B(n14), .C(n1020), .D(b[30]), .Y(n1537) );
  nr2d1_hd U1338 ( .A(DP_OP_116J3_127_7148_n3), .B(n1537), .Y(n1764) );
  oa22ad1_hd U1339 ( .A(n14), .B(n1843), .C(n1838), .D(n1764), .Y(n1536) );
  ao21d1_hd U1340 ( .A(DP_OP_116J3_127_7148_n3), .B(n1537), .C(n1536), .Y(n151) );
  ao22d1_hd U1341 ( .A(n1545), .B(n1544), .C(n1543), .D(n1542), .Y(n1547) );
  nr2d1_hd U1342 ( .A(n1547), .B(n1546), .Y(n1591) );
  ao22d1_hd U1343 ( .A(n1553), .B(b_s), .C(n1558), .D(z_s), .Y(n1550) );
  ivd1_hd U1344 ( .A(n1552), .Y(n1554) );
  nr2d1_hd U1345 ( .A(z_e[1]), .B(z_e[0]), .Y(n1582) );
  ivd1_hd U1346 ( .A(z_e[2]), .Y(n1578) );
  nr2d1_hd U1347 ( .A(z_e[3]), .B(n1577), .Y(n1574) );
  ivd1_hd U1348 ( .A(z_e[4]), .Y(n1571) );
  nr2d1_hd U1349 ( .A(z_e[5]), .B(n1570), .Y(n1567) );
  ivd1_hd U1350 ( .A(z_e[6]), .Y(n1564) );
  nr2d1_hd U1351 ( .A(z_m[23]), .B(z_e[0]), .Y(n1560) );
  ivd1_hd U1352 ( .A(z_e[1]), .Y(n1557) );
  nr4d1_hd U1353 ( .A(z_e[2]), .B(n1557), .C(n1556), .D(n1555), .Y(n1559) );
  oa211d1_hd U1354 ( .A(z_e[7]), .B(n1563), .C(n1580), .D(n1561), .Y(n1562) );
  scg15d1_hd U1355 ( .A(n1011), .B(z[30]), .C(n1586), .D(n1562), .Y(n230) );
  oa21d1_hd U1356 ( .A(n1567), .B(n1564), .C(n1563), .Y(n1565) );
  ao22d1_hd U1357 ( .A(n1011), .B(z[29]), .C(n1580), .D(n1565), .Y(n1566) );
  ao21d1_hd U1358 ( .A(z_e[5]), .B(n1570), .C(n1567), .Y(n1569) );
  oa211d1_hd U1359 ( .A(n1569), .B(n1587), .C(n1586), .D(n1568), .Y(n232) );
  oa21d1_hd U1360 ( .A(n1574), .B(n1571), .C(n1570), .Y(n1572) );
  ao22d1_hd U1361 ( .A(n1011), .B(z[27]), .C(n1580), .D(n1572), .Y(n1573) );
  ao21d1_hd U1362 ( .A(z_e[3]), .B(n1577), .C(n1574), .Y(n1576) );
  oa211d1_hd U1363 ( .A(n1576), .B(n1587), .C(n1586), .D(n1575), .Y(n234) );
  oa21d1_hd U1364 ( .A(n1582), .B(n1578), .C(n1577), .Y(n1579) );
  ao22d1_hd U1365 ( .A(n1011), .B(z[25]), .C(n1580), .D(n1579), .Y(n1581) );
  ao21d1_hd U1366 ( .A(z_e[0]), .B(z_e[1]), .C(n1582), .Y(n1584) );
  oa211d1_hd U1367 ( .A(n1584), .B(n1587), .C(n1586), .D(n1583), .Y(n236) );
  oa211d1_hd U1368 ( .A(z_e[0]), .B(n1587), .C(n1586), .D(n1585), .Y(n237) );
  scg17d1_hd U1369 ( .A(z_m[22]), .B(n1592), .C(n1591), .D(n1590), .Y(n238) );
  ao21d1_hd U1370 ( .A(n1711), .B(n1597), .C(n1707), .Y(n1600) );
  ivd1_hd U1371 ( .A(z_m[21]), .Y(n1599) );
  nr2d1_hd U1372 ( .A(z_m[22]), .B(n1686), .Y(n1715) );
  scg14d1_hd U1373 ( .A(n1595), .B(n1715), .C(n1710), .Y(n1596) );
  scg4d1_hd U1374 ( .A(n1714), .B(z_m[22]), .C(n1596), .D(z_m[21]), .E(n1012), 
        .F(product[48]), .G(z_m[23]), .H(n1705), .Y(n261) );
  oa22d1_hd U1375 ( .A(n1600), .B(n1599), .C(n1598), .D(n1597), .Y(n1602) );
  ao22d1_hd U1376 ( .A(z_m[22]), .B(n1705), .C(n1012), .D(product[47]), .Y(
        n1601) );
  oa21d1_hd U1377 ( .A(z_m[20]), .B(n1608), .C(n1710), .Y(n1606) );
  ivd1_hd U1378 ( .A(n105), .Y(n1702) );
  ao21d1_hd U1379 ( .A(n1702), .B(n1604), .C(n1707), .Y(n1609) );
  oa21d1_hd U1380 ( .A(z_m[19]), .B(n1686), .C(n1609), .Y(n1605) );
  scg4d1_hd U1381 ( .A(n1606), .B(z_m[19]), .C(n1605), .D(z_m[20]), .E(z_m[21]), .F(n1705), .G(n1012), .H(product[46]), .Y(n263) );
  ivd1_hd U1382 ( .A(z_m[19]), .Y(n1607) );
  ao22d1_hd U1383 ( .A(z_m[19]), .B(n1609), .C(n1608), .D(n1607), .Y(n1611) );
  ao22d1_hd U1384 ( .A(n1012), .B(product[45]), .C(z_m[20]), .D(n1705), .Y(
        n1610) );
  oa21d1_hd U1385 ( .A(z_m[18]), .B(n1620), .C(n1710), .Y(n1615) );
  ao21d1_hd U1386 ( .A(n1677), .B(n1613), .C(n1707), .Y(n1616) );
  oa21d1_hd U1387 ( .A(z_m[17]), .B(n1686), .C(n1616), .Y(n1614) );
  scg4d1_hd U1388 ( .A(n1615), .B(z_m[17]), .C(n1614), .D(z_m[18]), .E(z_m[19]), .F(n1705), .G(n1012), .H(product[44]), .Y(n265) );
  ao22d1_hd U1389 ( .A(n1012), .B(product[43]), .C(z_m[18]), .D(n1705), .Y(
        n1619) );
  ivd1_hd U1390 ( .A(n1616), .Y(n1617) );
  ao22d1_hd U1391 ( .A(z_m[16]), .B(n1713), .C(z_m[17]), .D(n1617), .Y(n1618)
         );
  oa211d1_hd U1392 ( .A(z_m[17]), .B(n1620), .C(n1619), .D(n1618), .Y(n266) );
  oa21d1_hd U1393 ( .A(z_m[16]), .B(n1626), .C(n1710), .Y(n1624) );
  ao21d1_hd U1394 ( .A(n1702), .B(n1622), .C(n1707), .Y(n1627) );
  oa21d1_hd U1395 ( .A(z_m[15]), .B(n1686), .C(n1627), .Y(n1623) );
  scg4d1_hd U1396 ( .A(n1624), .B(z_m[15]), .C(n1623), .D(z_m[16]), .E(z_m[17]), .F(n1705), .G(n1012), .H(product[42]), .Y(n267) );
  ivd1_hd U1397 ( .A(z_m[15]), .Y(n1625) );
  ao22d1_hd U1398 ( .A(z_m[15]), .B(n1627), .C(n1626), .D(n1625), .Y(n1629) );
  ao22d1_hd U1399 ( .A(n1012), .B(product[41]), .C(z_m[16]), .D(n1705), .Y(
        n1628) );
  oa21d1_hd U1400 ( .A(z_m[14]), .B(n1638), .C(n1710), .Y(n1633) );
  ao21d1_hd U1401 ( .A(n1677), .B(n1631), .C(n1707), .Y(n1634) );
  oa21d1_hd U1402 ( .A(z_m[13]), .B(n1686), .C(n1634), .Y(n1632) );
  scg4d1_hd U1403 ( .A(n1633), .B(z_m[13]), .C(n1632), .D(z_m[14]), .E(z_m[15]), .F(n1705), .G(n1012), .H(product[40]), .Y(n269) );
  ao22d1_hd U1404 ( .A(n1012), .B(product[39]), .C(z_m[14]), .D(n1705), .Y(
        n1637) );
  ivd1_hd U1405 ( .A(n1634), .Y(n1635) );
  ao22d1_hd U1406 ( .A(z_m[12]), .B(n1713), .C(z_m[13]), .D(n1635), .Y(n1636)
         );
  oa211d1_hd U1407 ( .A(z_m[13]), .B(n1638), .C(n1637), .D(n1636), .Y(n270) );
  oa21d1_hd U1408 ( .A(z_m[12]), .B(n1644), .C(n1710), .Y(n1642) );
  ao21d1_hd U1409 ( .A(n1677), .B(n1640), .C(n1707), .Y(n1645) );
  oa21d1_hd U1410 ( .A(z_m[11]), .B(n1686), .C(n1645), .Y(n1641) );
  scg4d1_hd U1411 ( .A(n1642), .B(z_m[11]), .C(n1641), .D(z_m[12]), .E(z_m[13]), .F(n1705), .G(n1012), .H(product[38]), .Y(n271) );
  ivd1_hd U1412 ( .A(z_m[11]), .Y(n1643) );
  ao22d1_hd U1413 ( .A(z_m[11]), .B(n1645), .C(n1644), .D(n1643), .Y(n1647) );
  ao22d1_hd U1414 ( .A(n1012), .B(product[37]), .C(z_m[12]), .D(n1705), .Y(
        n1646) );
  oa21d1_hd U1415 ( .A(z_m[10]), .B(n1656), .C(n1710), .Y(n1651) );
  ao21d1_hd U1416 ( .A(n1702), .B(n1649), .C(n1707), .Y(n1652) );
  oa21d1_hd U1417 ( .A(z_m[9]), .B(n1686), .C(n1652), .Y(n1650) );
  scg4d1_hd U1418 ( .A(n1651), .B(z_m[9]), .C(n1650), .D(z_m[10]), .E(z_m[11]), 
        .F(n1705), .G(n1012), .H(product[36]), .Y(n273) );
  ao22d1_hd U1419 ( .A(n1012), .B(product[35]), .C(z_m[10]), .D(n1705), .Y(
        n1655) );
  ivd1_hd U1420 ( .A(n1652), .Y(n1653) );
  ao22d1_hd U1421 ( .A(z_m[8]), .B(n1713), .C(z_m[9]), .D(n1653), .Y(n1654) );
  oa211d1_hd U1422 ( .A(z_m[9]), .B(n1656), .C(n1655), .D(n1654), .Y(n274) );
  oa21d1_hd U1423 ( .A(z_m[8]), .B(n1662), .C(n1710), .Y(n1660) );
  ao21d1_hd U1424 ( .A(n1677), .B(n1658), .C(n1707), .Y(n1663) );
  oa21d1_hd U1425 ( .A(z_m[7]), .B(n1686), .C(n1663), .Y(n1659) );
  scg4d1_hd U1426 ( .A(n1660), .B(z_m[7]), .C(n1659), .D(z_m[8]), .E(z_m[9]), 
        .F(n1705), .G(n1012), .H(product[34]), .Y(n275) );
  ivd1_hd U1427 ( .A(z_m[7]), .Y(n1661) );
  ao22d1_hd U1428 ( .A(z_m[7]), .B(n1663), .C(n1662), .D(n1661), .Y(n1665) );
  ao22d1_hd U1429 ( .A(n1012), .B(product[33]), .C(z_m[8]), .D(n1705), .Y(
        n1664) );
  oa21d1_hd U1430 ( .A(z_m[6]), .B(n1674), .C(n1710), .Y(n1669) );
  ao21d1_hd U1431 ( .A(n1702), .B(n1667), .C(n1707), .Y(n1670) );
  oa21d1_hd U1432 ( .A(z_m[5]), .B(n1686), .C(n1670), .Y(n1668) );
  scg4d1_hd U1433 ( .A(n1669), .B(z_m[5]), .C(n1668), .D(z_m[6]), .E(z_m[7]), 
        .F(n1705), .G(n1012), .H(product[32]), .Y(n277) );
  ao22d1_hd U1434 ( .A(n1012), .B(product[31]), .C(z_m[6]), .D(n1705), .Y(
        n1673) );
  ivd1_hd U1435 ( .A(n1670), .Y(n1671) );
  ao22d1_hd U1436 ( .A(z_m[4]), .B(n1713), .C(z_m[5]), .D(n1671), .Y(n1672) );
  oa211d1_hd U1437 ( .A(z_m[5]), .B(n1674), .C(n1673), .D(n1672), .Y(n278) );
  oa21d1_hd U1438 ( .A(z_m[4]), .B(n1681), .C(n1710), .Y(n1679) );
  ao21d1_hd U1439 ( .A(n1677), .B(n1676), .C(n1707), .Y(n1682) );
  oa21d1_hd U1440 ( .A(z_m[3]), .B(n1686), .C(n1682), .Y(n1678) );
  scg4d1_hd U1441 ( .A(n1679), .B(z_m[3]), .C(n1678), .D(z_m[4]), .E(z_m[5]), 
        .F(n1705), .G(n1012), .H(product[30]), .Y(n279) );
  ivd1_hd U1442 ( .A(z_m[3]), .Y(n1680) );
  ao22d1_hd U1443 ( .A(z_m[3]), .B(n1682), .C(n1681), .D(n1680), .Y(n1684) );
  ao22d1_hd U1444 ( .A(n1012), .B(product[29]), .C(z_m[4]), .D(n1705), .Y(
        n1683) );
  oa21d1_hd U1445 ( .A(z_m[2]), .B(n1685), .C(n1710), .Y(n1688) );
  nr2d1_hd U1446 ( .A(z_m[0]), .B(n1686), .Y(n1706) );
  nr2d1_hd U1447 ( .A(n1707), .B(n1706), .Y(n1690) );
  nd2bd1_hd U1448 ( .AN(z_m[1]), .B(n1711), .Y(n1689) );
  scg4d1_hd U1449 ( .A(n1688), .B(z_m[1]), .C(n1687), .D(z_m[2]), .E(z_m[3]), 
        .F(n1705), .G(n1012), .H(product[28]), .Y(n281) );
  ivd1_hd U1450 ( .A(n1690), .Y(n1691) );
  scg4d1_hd U1451 ( .A(n1692), .B(z_m[0]), .C(n1691), .D(z_m[1]), .E(z_m[2]), 
        .F(n1705), .G(n1012), .H(product[27]), .Y(n282) );
  nr4d1_hd U1452 ( .A(product[14]), .B(product[12]), .C(product[19]), .D(
        product[17]), .Y(n1696) );
  nr4d1_hd U1453 ( .A(product[15]), .B(product[8]), .C(product[20]), .D(
        product[4]), .Y(n1695) );
  nr4d1_hd U1454 ( .A(product[21]), .B(product[2]), .C(product[13]), .D(
        product[16]), .Y(n1694) );
  nr4d1_hd U1455 ( .A(product[23]), .B(product[5]), .C(product[22]), .D(
        product[18]), .Y(n1693) );
  nd4d1_hd U1456 ( .A(n1696), .B(n1695), .C(n1694), .D(n1693), .Y(n1697) );
  nr4d1_hd U1457 ( .A(product[9]), .B(product[7]), .C(n1698), .D(n1697), .Y(
        n1701) );
  ao22d1_hd U1458 ( .A(round_bit), .B(n1699), .C(sticky), .D(n1712), .Y(n1700)
         );
  oa21d1_hd U1459 ( .A(n1701), .B(n1712), .C(n1700), .Y(n283) );
  ao22d1_hd U1460 ( .A(n1012), .B(product[24]), .C(n1702), .D(round_bit), .Y(
        n1703) );
  oa21d1_hd U1461 ( .A(net922), .B(n1704), .C(n1703), .Y(n284) );
  ao22d1_hd U1462 ( .A(n1012), .B(product[26]), .C(z_m[1]), .D(n1705), .Y(
        n1709) );
  ao21d1_hd U1463 ( .A(n1707), .B(z_m[0]), .C(n1706), .Y(n1708) );
  oa211d1_hd U1464 ( .A(net922), .B(n1710), .C(n1709), .D(n1708), .Y(n285) );
  ao22d1_hd U1465 ( .A(z_m[22]), .B(n1713), .C(n1012), .D(product[49]), .Y(
        n1717) );
  oa21d1_hd U1466 ( .A(n1715), .B(n1714), .C(z_m[23]), .Y(n1716) );
  oa211d1_hd U1467 ( .A(n1719), .B(n1718), .C(n1717), .D(n1716), .Y(n286) );
  ao22d1_hd U1468 ( .A(n1004), .B(DP_OP_125J3_130_6300_n34), .C(z_e[0]), .D(
        n1844), .Y(n2863) );
  ao22d1_hd U1469 ( .A(n1019), .B(b[22]), .C(n1054), .D(n1742), .Y(n1721) );
  oa21d1_hd U1470 ( .A(n1053), .B(n1744), .C(n1721), .Y(n287) );
  ao22d1_hd U1471 ( .A(n1020), .B(b[20]), .C(n1050), .D(n1742), .Y(n1722) );
  oa21d1_hd U1472 ( .A(n1049), .B(n1744), .C(n1722), .Y(n288) );
  ao22d1_hd U1473 ( .A(n1019), .B(b[19]), .C(n1048), .D(n1742), .Y(n1723) );
  scg16d1_hd U1474 ( .A(n1047), .B(n1744), .C(n1723), .Y(n289) );
  ao22d1_hd U1475 ( .A(n1019), .B(b[18]), .C(n1047), .D(n1742), .Y(n1724) );
  oa21d1_hd U1476 ( .A(n1046), .B(n1744), .C(n1724), .Y(n290) );
  ao22d1_hd U1477 ( .A(n1019), .B(b[17]), .C(n1045), .D(n1742), .Y(n1725) );
  oa21d1_hd U1478 ( .A(n1044), .B(n1744), .C(n1725), .Y(n291) );
  ao22d1_hd U1479 ( .A(n1019), .B(b[16]), .C(n1008), .D(n1742), .Y(n1726) );
  oa21d1_hd U1480 ( .A(n1043), .B(n1744), .C(n1726), .Y(n292) );
  ao22d1_hd U1481 ( .A(n1019), .B(b[15]), .C(n1042), .D(n1742), .Y(n1727) );
  scg16d1_hd U1482 ( .A(n1041), .B(n1744), .C(n1727), .Y(n293) );
  ao22d1_hd U1483 ( .A(n1019), .B(b[14]), .C(n1041), .D(n1742), .Y(n1728) );
  oa21d1_hd U1484 ( .A(n1040), .B(n1744), .C(n1728), .Y(n294) );
  ao22d1_hd U1485 ( .A(n1019), .B(b[13]), .C(n1039), .D(n1742), .Y(n1729) );
  scg16d1_hd U1486 ( .A(n1038), .B(n1744), .C(n1729), .Y(n295) );
  ao22d1_hd U1487 ( .A(n1019), .B(b[12]), .C(n1038), .D(n1742), .Y(n1730) );
  scg16d1_hd U1488 ( .A(n1037), .B(n1744), .C(n1730), .Y(n296) );
  ao22d1_hd U1489 ( .A(n1019), .B(b[11]), .C(n1037), .D(n1742), .Y(n1731) );
  oa21d1_hd U1490 ( .A(n1036), .B(n1744), .C(n1731), .Y(n297) );
  ao22d1_hd U1491 ( .A(n1019), .B(b[10]), .C(n1035), .D(n1742), .Y(n1732) );
  scg16d1_hd U1492 ( .A(n1034), .B(n1744), .C(n1732), .Y(n298) );
  ao22d1_hd U1493 ( .A(n1019), .B(b[9]), .C(n1034), .D(n1742), .Y(n1733) );
  oa21d1_hd U1494 ( .A(n1033), .B(n1744), .C(n1733), .Y(n299) );
  ao22d1_hd U1495 ( .A(n1019), .B(b[8]), .C(n1032), .D(n1742), .Y(n1734) );
  oa21d1_hd U1496 ( .A(n1031), .B(n1744), .C(n1734), .Y(n300) );
  ao22d1_hd U1497 ( .A(n1019), .B(b[7]), .C(n1030), .D(n1742), .Y(n1735) );
  scg16d1_hd U1498 ( .A(n1029), .B(n1744), .C(n1735), .Y(n301) );
  ao22d1_hd U1499 ( .A(n1020), .B(b[6]), .C(n1029), .D(n1742), .Y(n1736) );
  scg16d1_hd U1500 ( .A(n1028), .B(n1744), .C(n1736), .Y(n302) );
  ao22d1_hd U1501 ( .A(n1020), .B(b[5]), .C(n1028), .D(n1742), .Y(n1737) );
  oa21d1_hd U1502 ( .A(n1027), .B(n1744), .C(n1737), .Y(n303) );
  ao22d1_hd U1503 ( .A(n1020), .B(b[4]), .C(n1006), .D(n1742), .Y(n1738) );
  oa21d1_hd U1504 ( .A(n1026), .B(n1744), .C(n1738), .Y(n304) );
  ao22d1_hd U1505 ( .A(n1020), .B(b[3]), .C(n1025), .D(n1742), .Y(n1739) );
  oa21d1_hd U1506 ( .A(n1024), .B(n1744), .C(n1739), .Y(n305) );
  ao22d1_hd U1507 ( .A(n1020), .B(b[2]), .C(n1007), .D(n1742), .Y(n1740) );
  oa21d1_hd U1508 ( .A(n1023), .B(n1744), .C(n1740), .Y(n306) );
  ao22d1_hd U1509 ( .A(n1020), .B(b[1]), .C(n1022), .D(n1742), .Y(n1741) );
  oa21d1_hd U1510 ( .A(n1009), .B(n1744), .C(n1741), .Y(n307) );
  ao22d1_hd U1511 ( .A(n1020), .B(b[21]), .C(n1052), .D(n1742), .Y(n1743) );
  oa21d1_hd U1512 ( .A(n1051), .B(n1744), .C(n1743), .Y(n309) );
  ao22d1_hd U1513 ( .A(n1850), .B(n1054), .C(b_m[23]), .D(n1118), .Y(n1746) );
  oa21d1_hd U1514 ( .A(n1747), .B(n1835), .C(n1746), .Y(n310) );
  oa211d1_hd U1515 ( .A(n1810), .B(n1749), .C(n1762), .D(n1748), .Y(n1751) );
  ao211d1_hd U1516 ( .A(a_e[8]), .B(n1833), .C(DP_OP_113J3_124_6892_n3), .D(
        n1750), .Y(n1759) );
  ao22d1_hd U1517 ( .A(a_e[8]), .B(n1751), .C(n1759), .D(n1757), .Y(n1752) );
  ao22d1_hd U1518 ( .A(a_e[1]), .B(n1754), .C(C81_DATA2_1), .D(n1757), .Y(
        n1753) );
  ao22d1_hd U1519 ( .A(n1020), .B(a[23]), .C(n1833), .D(a_e[0]), .Y(n1755) );
  ivd1_hd U1520 ( .A(n1755), .Y(n768) );
  nr2d1_hd U1521 ( .A(n1810), .B(n1761), .Y(n1758) );
  oa211d1_hd U1522 ( .A(n1759), .B(n1758), .C(n1757), .D(n1756), .Y(n1760) );
  oa211d1_hd U1523 ( .A(n1762), .B(n1761), .C(n138), .D(n1760), .Y(n319) );
  oa21d1_hd U1524 ( .A(n1763), .B(n1765), .C(n1764), .Y(n1840) );
  oa21d1_hd U1525 ( .A(n1765), .B(n1764), .C(n1843), .Y(n1766) );
  oa211d1_hd U1526 ( .A(n1840), .B(n1770), .C(n148), .D(n1767), .Y(n320) );
  ao22d1_hd U1527 ( .A(b_e[1]), .B(n1768), .C(n1838), .D(C82_DATA2_1), .Y(
        n1769) );
  oa22d1_hd U1528 ( .A(n1771), .B(n1843), .C(n1770), .D(n769), .Y(n327) );
  oa22d1_hd U1529 ( .A(n1832), .B(n1891), .C(n1783), .D(n1831), .Y(n328) );
  ao22d1_hd U1530 ( .A(n1020), .B(a[20]), .C(n1829), .D(a_m[20]), .Y(n1772) );
  oa21d1_hd U1531 ( .A(n1832), .B(n1773), .C(n1772), .Y(n329) );
  ao22d1_hd U1532 ( .A(n1020), .B(a[19]), .C(n1829), .D(a_m[19]), .Y(n1774) );
  oa21d1_hd U1533 ( .A(n1832), .B(n1775), .C(n1774), .Y(n330) );
  oa22d1_hd U1534 ( .A(n1832), .B(n1015), .C(n1783), .D(n1775), .Y(n331) );
  ao22d1_hd U1535 ( .A(n1020), .B(a[17]), .C(n1829), .D(a_m[17]), .Y(n1776) );
  oa21d1_hd U1536 ( .A(n1832), .B(n1777), .C(n1776), .Y(n332) );
  ao22d1_hd U1537 ( .A(n1020), .B(a[16]), .C(n1829), .D(a_m[16]), .Y(n1778) );
  oa21d1_hd U1538 ( .A(n1832), .B(n1779), .C(n1778), .Y(n333) );
  ao22d1_hd U1539 ( .A(n1020), .B(a[15]), .C(n1829), .D(a_m[15]), .Y(n1780) );
  oa21d1_hd U1540 ( .A(n1832), .B(n1869), .C(n1780), .Y(n334) );
  ao22d1_hd U1541 ( .A(n1019), .B(a[14]), .C(n1829), .D(a_m[14]), .Y(n1781) );
  oa21d1_hd U1542 ( .A(n1832), .B(n1782), .C(n1781), .Y(n335) );
  oa22d1_hd U1543 ( .A(n1832), .B(n1784), .C(n1783), .D(n1782), .Y(n336) );
  ao22d1_hd U1544 ( .A(n1019), .B(a[12]), .C(n1829), .D(a_m[12]), .Y(n1785) );
  oa21d1_hd U1545 ( .A(n1832), .B(n1017), .C(n1785), .Y(n337) );
  ao22d1_hd U1546 ( .A(n1019), .B(a[11]), .C(n1829), .D(a_m[11]), .Y(n1786) );
  oa21d1_hd U1547 ( .A(n1832), .B(n1787), .C(n1786), .Y(n338) );
  ao22d1_hd U1548 ( .A(n1019), .B(a[10]), .C(n1829), .D(a_m[10]), .Y(n1788) );
  oa21d1_hd U1549 ( .A(n1832), .B(n1789), .C(n1788), .Y(n339) );
  ao22d1_hd U1550 ( .A(n1019), .B(a[9]), .C(n1829), .D(a_m[9]), .Y(n1790) );
  oa21d1_hd U1551 ( .A(n1832), .B(n1013), .C(n1790), .Y(n340) );
  ao22d1_hd U1552 ( .A(n1019), .B(a[8]), .C(n1829), .D(a_m[8]), .Y(n1792) );
  oa21d1_hd U1553 ( .A(n1832), .B(n1793), .C(n1792), .Y(n341) );
  ao22d1_hd U1554 ( .A(n1019), .B(a[7]), .C(n1829), .D(a_m[7]), .Y(n1794) );
  oa21d1_hd U1555 ( .A(n1832), .B(n1795), .C(n1794), .Y(n342) );
  ao22d1_hd U1556 ( .A(n1020), .B(a[6]), .C(n1829), .D(a_m[6]), .Y(n1796) );
  oa21d1_hd U1557 ( .A(n1832), .B(n1014), .C(n1796), .Y(n343) );
  ao22d1_hd U1558 ( .A(n1019), .B(a[5]), .C(n1829), .D(a_m[5]), .Y(n1798) );
  oa21d1_hd U1559 ( .A(n1832), .B(n1799), .C(n1798), .Y(n344) );
  ao22d1_hd U1560 ( .A(n1019), .B(a[4]), .C(n1829), .D(a_m[4]), .Y(n1800) );
  oa21d1_hd U1561 ( .A(n1832), .B(n1801), .C(n1800), .Y(n345) );
  ao22d1_hd U1562 ( .A(n1019), .B(a[3]), .C(n1829), .D(a_m[3]), .Y(n1802) );
  oa21d1_hd U1563 ( .A(n1832), .B(n1016), .C(n1802), .Y(n346) );
  ao22d1_hd U1564 ( .A(n1019), .B(a[2]), .C(n1829), .D(a_m[2]), .Y(n1803) );
  oa21d1_hd U1565 ( .A(n1832), .B(n1804), .C(n1803), .Y(n347) );
  ao22d1_hd U1566 ( .A(n1019), .B(a[1]), .C(n1829), .D(a_m[1]), .Y(n1805) );
  oa21d1_hd U1567 ( .A(n1832), .B(n1806), .C(n1805), .Y(n348) );
  scg21d1_hd U1568 ( .A(n1808), .B(o_AB_ACK), .C(i_RST), .D(n1018), .Y(n350)
         );
  nr2d1_hd U1569 ( .A(n1810), .B(n1059), .Y(n1817) );
  nd3d1_hd U1570 ( .A(o_Z_STB), .B(i_Z_ACK), .C(n1021), .Y(n1811) );
  nd2bd1_hd U1571 ( .AN(i_RST), .B(n1811), .Y(n1849) );
  ao21d1_hd U1572 ( .A(b_m[23]), .B(n1850), .C(n1849), .Y(n1813) );
  oa211d1_hd U1573 ( .A(n1846), .B(n1822), .C(n1820), .D(n1812), .Y(n1825) );
  oa211d1_hd U1574 ( .A(n1815), .B(n1814), .C(n1813), .D(n1825), .Y(n1816) );
  nr2d1_hd U1575 ( .A(n1817), .B(n1816), .Y(n1828) );
  ao22d1_hd U1576 ( .A(n1821), .B(n1820), .C(n1833), .D(n1845), .Y(n1823) );
  oa22d1_hd U1577 ( .A(n1220), .B(n1823), .C(n1822), .D(n1845), .Y(n351) );
  oa22d1_hd U1578 ( .A(n1220), .B(n1825), .C(n1824), .D(n1845), .Y(n352) );
  nr2d1_hd U1579 ( .A(state[0]), .B(n1847), .Y(n1827) );
  ao22d1_hd U1580 ( .A(n1019), .B(a[22]), .C(n1829), .D(a_m[22]), .Y(n1830) );
  oa21d1_hd U1581 ( .A(n1832), .B(n1831), .C(n1830), .Y(n354) );
  ao22d1_hd U1582 ( .A(a_m[22]), .B(n1833), .C(n1058), .D(n1118), .Y(n1834) );
  oa21d1_hd U1583 ( .A(n1836), .B(n1835), .C(n1834), .Y(n355) );
  oa211d1_hd U1584 ( .A(n1840), .B(n1839), .C(n1838), .D(n1837), .Y(n1841) );
  oa211d1_hd U1585 ( .A(n1843), .B(n1842), .C(n148), .D(n1841), .Y(n356) );
  nr2d1_hd U1586 ( .A(n1010), .B(n1844), .Y(n1848) );
  oa22d1_hd U1587 ( .A(n1848), .B(n1847), .C(n1846), .D(n1845), .Y(n357) );
  scg20d1_hd U1588 ( .A(o_Z_STB), .B(n1021), .C(n1849), .Y(n358) );
  fad1_hd U1589 ( .A(n1853), .B(n1852), .CI(n1851), .CO(n1854), .S(
        intadd_8_B_5_) );
  ivd1_hd U1590 ( .A(n1854), .Y(n2033) );
  scg17d1_hd U1591 ( .A(n1856), .B(a_m[20]), .C(n1059), .D(n1855), .Y(n1863)
         );
  ao22d1_hd U1592 ( .A(b_m[23]), .B(n1903), .C(n1902), .D(n1857), .Y(n1858) );
  ivd1_hd U1593 ( .A(intadd_1_SUM_7_), .Y(n1873) );
  ao22d1_hd U1594 ( .A(b_m[23]), .B(n1932), .C(n1935), .D(n1928), .Y(n1865) );
  scg4d1_hd U1595 ( .A(n1936), .B(n1875), .C(n1052), .D(n1867), .E(n1866), .F(
        n1054), .G(n1050), .H(n1876), .Y(n1868) );
  ivd1_hd U1596 ( .A(n1870), .Y(n2030) );
  ivd1_hd U1597 ( .A(intadd_12_SUM_3_), .Y(n1885) );
  ao22d1_hd U1598 ( .A(b_m[23]), .B(n1876), .C(n1875), .D(n1928), .Y(n1877) );
  scg4d1_hd U1599 ( .A(n1936), .B(n1887), .C(n1052), .D(n1879), .E(n1878), .F(
        n1054), .G(n1888), .H(n1050), .Y(n1880) );
  ao22d1_hd U1600 ( .A(b_m[23]), .B(n1888), .C(n1887), .D(n1928), .Y(n1889) );
  scg4d1_hd U1601 ( .A(n1936), .B(n1918), .C(n1052), .D(n1919), .E(n1921), .F(
        n1054), .G(n1920), .H(n1050), .Y(n1890) );
  ivd1_hd U1602 ( .A(n1892), .Y(n2026) );
  fad1_hd U1603 ( .A(intadd_11_SUM_4_), .B(n1894), .CI(n1893), .CO(n1895), .S(
        n1892) );
  ao22d1_hd U1604 ( .A(b_m[23]), .B(n1920), .C(n1918), .D(n1928), .Y(n1896) );
  scg4d1_hd U1605 ( .A(n1936), .B(n1902), .C(n1052), .D(n1903), .E(n1905), .F(
        n1054), .G(n1050), .H(n1904), .Y(n1897) );
  ivd1_hd U1606 ( .A(n1901), .Y(n2023) );
  scg4d1_hd U1607 ( .A(n1006), .B(n1905), .C(n1007), .D(n1904), .E(n1903), .F(
        n1025), .G(n1902), .H(intadd_3_SUM_0_), .Y(n1906) );
  ao21d1_hd U1608 ( .A(n1909), .B(n1908), .C(n1907), .Y(n1916) );
  nr2d1_hd U1609 ( .A(n1059), .B(n1023), .Y(n1915) );
  ivd1_hd U1610 ( .A(n1910), .Y(n2022) );
  fad1_hd U1611 ( .A(n1016), .B(n1912), .CI(n1911), .CO(n1852), .S(n1914) );
  ivd1_hd U1612 ( .A(n1914), .Y(n1926) );
  fad1_hd U1613 ( .A(n1917), .B(n1916), .CI(n1915), .CO(n1925), .S(n1910) );
  scg4d1_hd U1614 ( .A(n1032), .B(n1921), .C(n1029), .D(n1920), .E(n1030), .F(
        n1919), .G(n1918), .H(intadd_3_SUM_4_), .Y(n1922) );
  ivd1_hd U1615 ( .A(n1923), .Y(n2021) );
  fad1_hd U1616 ( .A(n1926), .B(n1925), .CI(n1924), .CO(n1927), .S(n1923) );
  ivd1_hd U1617 ( .A(n1927), .Y(n2020) );
  ao22d1_hd U1618 ( .A(b_m[23]), .B(n1005), .C(n1929), .D(n1928), .Y(n1931) );
  scg4d1_hd U1619 ( .A(n1936), .B(n1935), .C(n1052), .D(n1934), .E(n1933), .F(
        n1054), .G(n1050), .H(n1932), .Y(n1937) );
  ivd1_hd U1620 ( .A(n1939), .Y(n2019) );
  fad1_hd U1621 ( .A(intadd_6_SUM_12_), .B(n1941), .CI(n1940), .CO(n1942), .S(
        n1939) );
  ivd1_hd U1622 ( .A(n1942), .Y(n2018) );
  ivd1_hd U1623 ( .A(intadd_10_B_2_), .Y(n1225) );
  ivd1_hd U1624 ( .A(intadd_10_SUM_0_), .Y(n1224) );
  ivd1_hd U1625 ( .A(intadd_11_B_1_), .Y(n1222) );
  ivd1_hd U1626 ( .A(intadd_15_B_1_), .Y(n1221) );
  ivd1_hd U1627 ( .A(intadd_10_SUM_1_), .Y(n1211) );
  ivd1_hd U1628 ( .A(intadd_1_SUM_1_), .Y(n1210) );
  ivd1_hd U1629 ( .A(intadd_1_SUM_2_), .Y(n1208) );
  ivd1_hd U1630 ( .A(intadd_12_SUM_0_), .Y(n1206) );
  ivd1_hd U1631 ( .A(intadd_19_SUM_0_), .Y(n1205) );
  ivd1_hd U1632 ( .A(intadd_12_SUM_1_), .Y(n1204) );
  ivd1_hd U1633 ( .A(intadd_19_SUM_1_), .Y(n1203) );
  ivd1_hd U1634 ( .A(intadd_11_SUM_0_), .Y(n1202) );
  ivd1_hd U1635 ( .A(intadd_1_SUM_3_), .Y(n1201) );
  ivd1_hd U1636 ( .A(intadd_1_SUM_4_), .Y(n1200) );
  ivd1_hd U1637 ( .A(intadd_1_SUM_5_), .Y(n1199) );
  ivd1_hd U1638 ( .A(intadd_12_SUM_2_), .Y(n1197) );
  ivd1_hd U1639 ( .A(intadd_19_SUM_2_), .Y(n1196) );
  ivd1_hd U1640 ( .A(intadd_19_n1), .Y(n1195) );
  ivd1_hd U1641 ( .A(intadd_13_SUM_0_), .Y(n1194) );
  ivd1_hd U1642 ( .A(intadd_16_SUM_0_), .Y(n1193) );
  ivd1_hd U1643 ( .A(intadd_17_SUM_0_), .Y(n1192) );
  ivd1_hd U1644 ( .A(intadd_13_SUM_1_), .Y(n1191) );
  ivd1_hd U1645 ( .A(intadd_16_SUM_1_), .Y(n1190) );
  ivd1_hd U1646 ( .A(intadd_17_SUM_1_), .Y(n1189) );
  ivd1_hd U1647 ( .A(intadd_10_n1), .Y(n1188) );
  ivd1_hd U1648 ( .A(intadd_15_SUM_0_), .Y(n1187) );
  ivd1_hd U1649 ( .A(intadd_1_SUM_6_), .Y(n1186) );
  ivd1_hd U1650 ( .A(intadd_15_SUM_2_), .Y(n1185) );
  ivd1_hd U1651 ( .A(intadd_18_SUM_2_), .Y(n1181) );
  ivd1_hd U1652 ( .A(intadd_18_n1), .Y(n1180) );
  ivd1_hd U1653 ( .A(intadd_17_n1), .Y(n1178) );
  ivd1_hd U1654 ( .A(intadd_16_n1), .Y(n1176) );
  ivd1_hd U1655 ( .A(intadd_0_SUM_0_), .Y(n1163) );
  ivd1_hd U1656 ( .A(intadd_0_SUM_1_), .Y(n1161) );
  ivd1_hd U1657 ( .A(intadd_0_SUM_2_), .Y(n1160) );
  ivd1_hd U1658 ( .A(intadd_0_SUM_3_), .Y(n1159) );
  ivd1_hd U1659 ( .A(intadd_0_SUM_4_), .Y(n1157) );
  ivd1_hd U1660 ( .A(intadd_0_SUM_5_), .Y(n1156) );
  ivd1_hd U1661 ( .A(intadd_0_SUM_6_), .Y(n1155) );
  ivd1_hd U1662 ( .A(intadd_0_SUM_7_), .Y(n1153) );
  ivd1_hd U1663 ( .A(intadd_0_SUM_8_), .Y(n1152) );
  ivd1_hd U1664 ( .A(intadd_0_SUM_9_), .Y(n1151) );
  ivd1_hd U1665 ( .A(intadd_0_SUM_10_), .Y(n1149) );
  ivd1_hd U1666 ( .A(intadd_0_SUM_11_), .Y(n1147) );
  ivd1_hd U1667 ( .A(intadd_0_SUM_12_), .Y(n1146) );
  ivd1_hd U1668 ( .A(intadd_0_SUM_13_), .Y(n1144) );
  ivd1_hd U1669 ( .A(intadd_0_SUM_14_), .Y(n1143) );
  ivd1_hd U1670 ( .A(intadd_0_SUM_15_), .Y(n1142) );
  ivd1_hd U1671 ( .A(intadd_0_SUM_16_), .Y(n1140) );
  ivd1_hd U1672 ( .A(intadd_0_SUM_17_), .Y(n1139) );
  ivd1_hd U1673 ( .A(intadd_0_SUM_18_), .Y(n1138) );
  ivd1_hd U1674 ( .A(intadd_0_SUM_19_), .Y(n1137) );
  ivd1_hd U1675 ( .A(intadd_0_SUM_20_), .Y(n1135) );
  ivd1_hd U1676 ( .A(intadd_0_SUM_21_), .Y(n1134) );
  ivd1_hd U1677 ( .A(intadd_0_SUM_22_), .Y(n1133) );
  ivd1_hd U1678 ( .A(intadd_0_SUM_23_), .Y(n1131) );
  ivd1_hd U1679 ( .A(intadd_5_SUM_15_), .Y(n1130) );
  ivd1_hd U1680 ( .A(intadd_9_SUM_0_), .Y(n1129) );
  ivd1_hd U1681 ( .A(intadd_0_SUM_24_), .Y(n1128) );
  ivd1_hd U1682 ( .A(intadd_5_SUM_16_), .Y(n1126) );
  ivd1_hd U1683 ( .A(intadd_5_n1), .Y(n1125) );
  ivd1_hd U1684 ( .A(intadd_20_SUM_2_), .Y(n1124) );
  ivd1_hd U1685 ( .A(intadd_20_n1), .Y(n1123) );
  ivd1_hd U1686 ( .A(intadd_6_SUM_13_), .Y(n1122) );
  ivd1_hd U1687 ( .A(intadd_6_n1), .Y(n1121) );
  ivd1_hd U1688 ( .A(n2863), .Y(n1103) );
endmodule


module float_multiplier_0 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, 
        i_Z_ACK, i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N34, a_s, b_s, N35, round_bit, sticky, z_s, N176, N177, N178, N179,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, C82_DATA2_1, C82_DATA2_2,
         C82_DATA2_3, C82_DATA2_4, C82_DATA2_5, C82_DATA2_6, C81_DATA2_1,
         C81_DATA2_2, C81_DATA2_3, C81_DATA2_4, C81_DATA2_5, C81_DATA2_6,
         net922, n10, n14, n104, n105, n110, n138, n141, n148, n151, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359,
         DP_OP_116J3_127_7148_n3, DP_OP_116J3_127_7148_n4,
         DP_OP_116J3_127_7148_n5, DP_OP_116J3_127_7148_n6,
         DP_OP_116J3_127_7148_n7, DP_OP_116J3_127_7148_n8,
         DP_OP_113J3_124_6892_n3, DP_OP_113J3_124_6892_n4,
         DP_OP_113J3_124_6892_n5, DP_OP_113J3_124_6892_n6,
         DP_OP_113J3_124_6892_n7, DP_OP_113J3_124_6892_n8, C1_Z_6, C1_Z_5,
         C1_Z_4, C1_Z_3, C1_Z_2, C1_Z_1, DP_OP_125J3_130_6300_n42,
         DP_OP_125J3_130_6300_n41, DP_OP_125J3_130_6300_n40,
         DP_OP_125J3_130_6300_n39, DP_OP_125J3_130_6300_n38,
         DP_OP_125J3_130_6300_n37, DP_OP_125J3_130_6300_n36,
         DP_OP_125J3_130_6300_n35, DP_OP_125J3_130_6300_n34,
         DP_OP_125J3_130_6300_n32, DP_OP_125J3_130_6300_n31,
         DP_OP_125J3_130_6300_n30, DP_OP_125J3_130_6300_n29,
         DP_OP_125J3_130_6300_n28, DP_OP_125J3_130_6300_n27,
         DP_OP_125J3_130_6300_n26, DP_OP_125J3_130_6300_n25,
         DP_OP_125J3_130_6300_n20, DP_OP_125J3_130_6300_n19,
         DP_OP_125J3_130_6300_n18, DP_OP_125J3_130_6300_n17,
         DP_OP_125J3_130_6300_n16, DP_OP_125J3_130_6300_n15,
         DP_OP_125J3_130_6300_n14, DP_OP_125J3_130_6300_n13,
         DP_OP_125J3_130_6300_n12, DP_OP_125J3_130_6300_n9,
         DP_OP_125J3_130_6300_n8, DP_OP_125J3_130_6300_n7,
         DP_OP_125J3_130_6300_n6, DP_OP_125J3_130_6300_n5,
         DP_OP_125J3_130_6300_n4, DP_OP_125J3_130_6300_n3,
         DP_OP_125J3_130_6300_n2, n768, n769, n770, n771, n772, n773, n774,
         n775, intadd_24_CI, intadd_24_SUM_17_, intadd_24_SUM_16_,
         intadd_24_SUM_15_, intadd_24_SUM_14_, intadd_24_SUM_13_,
         intadd_24_SUM_12_, intadd_24_SUM_11_, intadd_24_SUM_10_,
         intadd_24_SUM_9_, intadd_24_SUM_8_, intadd_24_SUM_7_,
         intadd_24_SUM_6_, intadd_24_SUM_5_, intadd_24_SUM_4_,
         intadd_24_SUM_3_, intadd_24_SUM_2_, intadd_24_SUM_1_,
         intadd_24_SUM_0_, intadd_24_n18, intadd_24_n17, intadd_24_n16,
         intadd_24_n15, intadd_24_n14, intadd_24_n13, intadd_24_n12,
         intadd_24_n11, intadd_24_n10, intadd_24_n9, intadd_24_n8,
         intadd_24_n7, intadd_24_n6, intadd_24_n5, intadd_24_n4, intadd_24_n3,
         intadd_24_n2, intadd_24_n1, intadd_26_A_16_, intadd_26_A_15_,
         intadd_26_A_13_, intadd_26_A_12_, intadd_26_A_11_, intadd_26_A_10_,
         intadd_26_A_9_, intadd_26_A_8_, intadd_26_A_7_, intadd_26_A_6_,
         intadd_26_A_5_, intadd_26_A_4_, intadd_26_A_3_, intadd_26_A_2_,
         intadd_26_A_1_, intadd_26_A_0_, intadd_26_B_16_, intadd_26_B_15_,
         intadd_26_B_14_, intadd_26_B_13_, intadd_26_B_12_, intadd_26_B_11_,
         intadd_26_B_10_, intadd_26_B_9_, intadd_26_B_8_, intadd_26_B_7_,
         intadd_26_B_6_, intadd_26_B_5_, intadd_26_B_4_, intadd_26_B_3_,
         intadd_26_B_2_, intadd_26_B_1_, intadd_26_B_0_, intadd_26_CI,
         intadd_26_SUM_16_, intadd_26_SUM_15_, intadd_26_SUM_14_,
         intadd_26_SUM_13_, intadd_26_SUM_12_, intadd_26_SUM_11_,
         intadd_26_SUM_10_, intadd_26_SUM_9_, intadd_26_SUM_8_,
         intadd_26_SUM_7_, intadd_26_SUM_6_, intadd_26_SUM_5_,
         intadd_26_SUM_4_, intadd_26_SUM_3_, intadd_26_SUM_2_,
         intadd_26_SUM_1_, intadd_26_SUM_0_, intadd_26_n17, intadd_26_n16,
         intadd_26_n15, intadd_26_n14, intadd_26_n13, intadd_26_n12,
         intadd_26_n11, intadd_26_n10, intadd_26_n9, intadd_26_n8,
         intadd_26_n7, intadd_26_n6, intadd_26_n5, intadd_26_n4, intadd_26_n3,
         intadd_26_n2, intadd_26_n1, intadd_27_A_13_, intadd_27_A_11_,
         intadd_27_A_10_, intadd_27_A_9_, intadd_27_A_8_, intadd_27_A_7_,
         intadd_27_A_6_, intadd_27_A_5_, intadd_27_A_4_, intadd_27_A_3_,
         intadd_27_A_2_, intadd_27_A_1_, intadd_27_A_0_, intadd_27_B_13_,
         intadd_27_B_12_, intadd_27_B_11_, intadd_27_B_10_, intadd_27_B_9_,
         intadd_27_B_8_, intadd_27_B_7_, intadd_27_B_6_, intadd_27_B_5_,
         intadd_27_B_4_, intadd_27_B_3_, intadd_27_B_2_, intadd_27_B_1_,
         intadd_27_B_0_, intadd_27_CI, intadd_27_SUM_13_, intadd_27_SUM_12_,
         intadd_27_SUM_11_, intadd_27_SUM_10_, intadd_27_SUM_9_,
         intadd_27_SUM_8_, intadd_27_SUM_7_, intadd_27_SUM_6_,
         intadd_27_SUM_5_, intadd_27_SUM_4_, intadd_27_SUM_3_,
         intadd_27_SUM_2_, intadd_27_SUM_1_, intadd_27_SUM_0_, intadd_27_n14,
         intadd_27_n13, intadd_27_n12, intadd_27_n11, intadd_27_n10,
         intadd_27_n9, intadd_27_n8, intadd_27_n7, intadd_27_n6, intadd_27_n5,
         intadd_27_n4, intadd_27_n3, intadd_27_n2, intadd_27_n1,
         intadd_28_A_10_, intadd_28_A_8_, intadd_28_A_7_, intadd_28_A_6_,
         intadd_28_A_5_, intadd_28_A_4_, intadd_28_A_3_, intadd_28_A_2_,
         intadd_28_A_1_, intadd_28_A_0_, intadd_28_B_9_, intadd_28_B_2_,
         intadd_28_B_1_, intadd_28_B_0_, intadd_28_CI, intadd_28_n11,
         intadd_28_n10, intadd_28_n9, intadd_28_n8, intadd_28_n7, intadd_28_n6,
         intadd_28_n5, intadd_28_n4, intadd_28_n3, intadd_28_n2, intadd_28_n1,
         intadd_29_A_4_, intadd_29_A_2_, intadd_29_A_1_, intadd_29_A_0_,
         intadd_29_B_8_, intadd_29_B_7_, intadd_29_B_6_, intadd_29_B_5_,
         intadd_29_B_3_, intadd_29_B_2_, intadd_29_B_1_, intadd_29_B_0_,
         intadd_29_CI, intadd_29_n9, intadd_29_n8, intadd_29_n7, intadd_29_n6,
         intadd_29_n5, intadd_29_n4, intadd_29_n3, intadd_29_n2, intadd_29_n1,
         intadd_31_A_5_, intadd_31_A_4_, intadd_31_A_3_, intadd_31_A_2_,
         intadd_31_B_7_, intadd_31_B_6_, intadd_31_B_4_, intadd_31_B_3_,
         intadd_31_B_2_, intadd_31_B_1_, intadd_31_CI, intadd_31_SUM_7_,
         intadd_31_SUM_6_, intadd_31_SUM_5_, intadd_31_SUM_4_,
         intadd_31_SUM_3_, intadd_31_SUM_2_, intadd_31_SUM_1_,
         intadd_31_SUM_0_, intadd_31_n8, intadd_31_n7, intadd_31_n6,
         intadd_31_n5, intadd_31_n4, intadd_31_n3, intadd_31_n2, intadd_31_n1,
         intadd_32_A_4_, intadd_32_A_3_, intadd_32_A_2_, intadd_32_A_1_,
         intadd_32_B_5_, intadd_32_B_3_, intadd_32_B_2_, intadd_32_B_1_,
         intadd_32_B_0_, intadd_32_CI, intadd_32_SUM_5_, intadd_32_SUM_4_,
         intadd_32_SUM_3_, intadd_32_SUM_2_, intadd_32_SUM_1_,
         intadd_32_SUM_0_, intadd_32_n6, intadd_32_n5, intadd_32_n4,
         intadd_32_n3, intadd_32_n2, intadd_32_n1, intadd_33_A_1_,
         intadd_33_B_4_, intadd_33_B_2_, intadd_33_B_1_, intadd_33_B_0_,
         intadd_33_CI, intadd_33_SUM_4_, intadd_33_SUM_3_, intadd_33_SUM_2_,
         intadd_33_SUM_1_, intadd_33_SUM_0_, intadd_33_n5, intadd_33_n4,
         intadd_33_n3, intadd_33_n2, intadd_33_n1, intadd_34_A_1_,
         intadd_34_A_0_, intadd_34_B_2_, intadd_34_B_1_, intadd_34_B_0_,
         intadd_34_CI, intadd_34_SUM_2_, intadd_34_SUM_1_, intadd_34_SUM_0_,
         intadd_34_n3, intadd_34_n2, intadd_34_n1, intadd_35_A_1_,
         intadd_35_B_2_, intadd_35_B_0_, intadd_35_CI, intadd_35_SUM_2_,
         intadd_35_SUM_1_, intadd_35_SUM_0_, intadd_35_n3, intadd_35_n2,
         intadd_35_n1, intadd_36_A_2_, intadd_36_A_1_, intadd_36_B_2_,
         intadd_36_B_1_, intadd_36_B_0_, intadd_36_CI, intadd_36_SUM_2_,
         intadd_36_SUM_1_, intadd_36_SUM_0_, intadd_36_n3, intadd_36_n2,
         intadd_36_n1, intadd_37_A_0_, intadd_37_B_2_, intadd_37_B_1_,
         intadd_37_B_0_, intadd_37_SUM_2_, intadd_37_SUM_1_, intadd_37_SUM_0_,
         intadd_37_n3, intadd_37_n2, intadd_37_n1, intadd_38_B_2_,
         intadd_38_B_1_, intadd_38_B_0_, intadd_38_CI, intadd_38_SUM_2_,
         intadd_38_SUM_1_, intadd_38_SUM_0_, intadd_38_n3, intadd_38_n2,
         intadd_38_n1, intadd_39_B_2_, intadd_39_B_1_, intadd_39_B_0_,
         intadd_39_CI, intadd_39_SUM_2_, intadd_39_n3, intadd_39_n2,
         intadd_39_n1, intadd_40_B_2_, intadd_40_B_1_, intadd_40_B_0_,
         intadd_40_CI, intadd_40_SUM_2_, intadd_40_SUM_1_, intadd_40_SUM_0_,
         intadd_40_n3, intadd_40_n2, intadd_40_n1, intadd_41_A_1_,
         intadd_41_A_0_, intadd_41_B_2_, intadd_41_CI, intadd_41_SUM_2_,
         intadd_41_n3, intadd_41_n2, intadd_41_n1, intadd_21_A_24_,
         intadd_21_A_23_, intadd_21_A_22_, intadd_21_A_21_, intadd_21_A_20_,
         intadd_21_A_19_, intadd_21_A_18_, intadd_21_A_17_, intadd_21_A_16_,
         intadd_21_A_15_, intadd_21_A_14_, intadd_21_A_13_, intadd_21_A_12_,
         intadd_21_A_11_, intadd_21_A_10_, intadd_21_A_9_, intadd_21_A_8_,
         intadd_21_A_7_, intadd_21_A_6_, intadd_21_A_5_, intadd_21_A_4_,
         intadd_21_A_3_, intadd_21_A_2_, intadd_21_A_1_, intadd_21_A_0_,
         intadd_21_B_21_, intadd_21_B_20_, intadd_21_B_19_, intadd_21_B_18_,
         intadd_21_B_17_, intadd_21_B_16_, intadd_21_B_15_, intadd_21_B_14_,
         intadd_21_B_13_, intadd_21_B_12_, intadd_21_B_11_, intadd_21_B_10_,
         intadd_21_B_9_, intadd_21_B_8_, intadd_21_B_7_, intadd_21_B_6_,
         intadd_21_B_5_, intadd_21_B_4_, intadd_21_B_3_, intadd_21_B_2_,
         intadd_21_B_1_, intadd_21_B_0_, intadd_21_CI, intadd_21_SUM_24_,
         intadd_21_SUM_23_, intadd_21_SUM_22_, intadd_21_SUM_21_,
         intadd_21_SUM_20_, intadd_21_SUM_19_, intadd_21_SUM_18_,
         intadd_21_SUM_17_, intadd_21_SUM_16_, intadd_21_SUM_15_,
         intadd_21_SUM_14_, intadd_21_SUM_13_, intadd_21_SUM_12_,
         intadd_21_SUM_11_, intadd_21_SUM_10_, intadd_21_SUM_9_,
         intadd_21_SUM_8_, intadd_21_SUM_7_, intadd_21_SUM_6_,
         intadd_21_SUM_5_, intadd_21_SUM_4_, intadd_21_SUM_3_,
         intadd_21_SUM_2_, intadd_21_SUM_1_, intadd_21_SUM_0_, intadd_21_n25,
         intadd_21_n24, intadd_21_n23, intadd_21_n22, intadd_21_n21,
         intadd_21_n20, intadd_21_n19, intadd_21_n18, intadd_21_n17,
         intadd_21_n16, intadd_21_n15, intadd_21_n14, intadd_21_n13,
         intadd_21_n12, intadd_21_n11, intadd_21_n10, intadd_21_n9,
         intadd_21_n8, intadd_21_n7, intadd_21_n6, intadd_21_n5, intadd_21_n4,
         intadd_21_n3, intadd_21_n2, intadd_21_n1, intadd_22_B_19_,
         intadd_22_B_8_, intadd_22_B_6_, intadd_22_B_5_, intadd_22_B_3_,
         intadd_22_B_2_, intadd_22_B_0_, intadd_22_CI, intadd_22_SUM_8_,
         intadd_22_SUM_7_, intadd_22_SUM_6_, intadd_22_SUM_5_,
         intadd_22_SUM_4_, intadd_22_SUM_3_, intadd_22_SUM_2_,
         intadd_22_SUM_1_, intadd_22_SUM_0_, intadd_22_n20, intadd_22_n19,
         intadd_22_n18, intadd_22_n17, intadd_22_n16, intadd_22_n15,
         intadd_22_n14, intadd_22_n13, intadd_22_n12, intadd_22_n11,
         intadd_22_n10, intadd_22_n9, intadd_22_n8, intadd_22_n7, intadd_22_n6,
         intadd_22_n5, intadd_22_n4, intadd_22_n3, intadd_22_n2, intadd_22_n1,
         intadd_23_A_18_, intadd_23_A_17_, intadd_23_A_16_, intadd_23_A_15_,
         intadd_23_A_14_, intadd_23_A_13_, intadd_23_A_12_, intadd_23_A_11_,
         intadd_23_A_10_, intadd_23_A_9_, intadd_23_A_8_, intadd_23_A_7_,
         intadd_23_A_6_, intadd_23_A_5_, intadd_23_A_4_, intadd_23_A_3_,
         intadd_23_A_2_, intadd_23_A_1_, intadd_23_A_0_, intadd_23_B_18_,
         intadd_23_B_17_, intadd_23_B_16_, intadd_23_B_15_, intadd_23_B_14_,
         intadd_23_B_13_, intadd_23_B_12_, intadd_23_B_11_, intadd_23_B_10_,
         intadd_23_B_9_, intadd_23_B_8_, intadd_23_B_7_, intadd_23_B_6_,
         intadd_23_B_5_, intadd_23_B_4_, intadd_23_B_3_, intadd_23_B_2_,
         intadd_23_B_1_, intadd_23_B_0_, intadd_23_CI, intadd_23_n19,
         intadd_23_n18, intadd_23_n17, intadd_23_n16, intadd_23_n15,
         intadd_23_n14, intadd_23_n13, intadd_23_n12, intadd_23_n11,
         intadd_23_n10, intadd_23_n9, intadd_23_n8, intadd_23_n7, intadd_23_n6,
         intadd_23_n5, intadd_23_n4, intadd_23_n3, intadd_23_n2, intadd_23_n1,
         intadd_25_A_15_, intadd_25_A_13_, intadd_25_A_10_, intadd_25_A_2_,
         intadd_25_A_1_, intadd_25_A_0_, intadd_25_B_16_, intadd_25_B_14_,
         intadd_25_B_12_, intadd_25_B_11_, intadd_25_B_9_, intadd_25_B_8_,
         intadd_25_B_7_, intadd_25_B_6_, intadd_25_B_5_, intadd_25_B_4_,
         intadd_25_B_3_, intadd_25_B_2_, intadd_25_B_1_, intadd_25_B_0_,
         intadd_25_CI, intadd_25_n17, intadd_25_n16, intadd_25_n15,
         intadd_25_n14, intadd_25_n13, intadd_25_n12, intadd_25_n11,
         intadd_25_n10, intadd_25_n9, intadd_25_n8, intadd_25_n7, intadd_25_n6,
         intadd_25_n5, intadd_25_n4, intadd_25_n3, intadd_25_n2, intadd_25_n1,
         intadd_30_B_0_, intadd_30_CI, intadd_30_SUM_0_, intadd_30_n8,
         intadd_30_n7, intadd_30_n6, intadd_30_n5, intadd_30_n4, intadd_30_n3,
         intadd_30_n2, intadd_30_n1, n1004, n1005, n1007, n1106, n1112, n1113,
         n1120, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1137, n1138, n1139, n1141, n1142, n1143, n1145, n1147,
         n1148, n1149, n1151, n1152, n1154, n1156, n1157, n1158, n1160, n1161,
         n1162, n1164, n1165, n1166, n1168, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1212, n1213, n1215, n1221, n1222,
         n1224, n1225, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1107, n1108, n1109,
         n1110, n1111, n1114, n1115, n1116, n1117, n1118, n1119, n1121, n1122,
         n1123, n1124, n1136, n1140, n1144, n1146, n1150, n1153, n1155, n1159,
         n1163, n1167, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1202, n1211, n1214, n1216, n1217, n1218, n1219,
         n1220, n1223, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [23:0] a_m;
  wire   [9:0] b_e;
  wire   [23:1] b_m;
  wire   [49:2] product;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U364 ( .A(i_RST), .Y(N34) );
  fad1_hd DP_OP_116J3_127_7148_U6 ( .A(n1007), .B(n775), .CI(
        DP_OP_116J3_127_7148_n4), .CO(DP_OP_116J3_127_7148_n3), .S(C82_DATA2_6) );
  fad1_hd DP_OP_116J3_127_7148_U7 ( .A(n1007), .B(n774), .CI(
        DP_OP_116J3_127_7148_n5), .CO(DP_OP_116J3_127_7148_n4), .S(C82_DATA2_5) );
  fad1_hd DP_OP_116J3_127_7148_U8 ( .A(n1007), .B(n773), .CI(
        DP_OP_116J3_127_7148_n6), .CO(DP_OP_116J3_127_7148_n5), .S(C82_DATA2_4) );
  fad1_hd DP_OP_116J3_127_7148_U9 ( .A(n1007), .B(n772), .CI(
        DP_OP_116J3_127_7148_n7), .CO(DP_OP_116J3_127_7148_n6), .S(C82_DATA2_3) );
  fad1_hd DP_OP_116J3_127_7148_U10 ( .A(n1007), .B(n771), .CI(
        DP_OP_116J3_127_7148_n8), .CO(DP_OP_116J3_127_7148_n7), .S(C82_DATA2_2) );
  fad1_hd DP_OP_116J3_127_7148_U11 ( .A(n1007), .B(n770), .CI(n769), .CO(
        DP_OP_116J3_127_7148_n8), .S(C82_DATA2_1) );
  fad1_hd DP_OP_113J3_124_6892_U6 ( .A(n1007), .B(C1_Z_6), .CI(
        DP_OP_113J3_124_6892_n4), .CO(DP_OP_113J3_124_6892_n3), .S(C81_DATA2_6) );
  fad1_hd DP_OP_113J3_124_6892_U7 ( .A(n1007), .B(C1_Z_5), .CI(
        DP_OP_113J3_124_6892_n5), .CO(DP_OP_113J3_124_6892_n4), .S(C81_DATA2_5) );
  fad1_hd DP_OP_113J3_124_6892_U8 ( .A(n1007), .B(C1_Z_4), .CI(
        DP_OP_113J3_124_6892_n6), .CO(DP_OP_113J3_124_6892_n5), .S(C81_DATA2_4) );
  fad1_hd DP_OP_113J3_124_6892_U9 ( .A(n1007), .B(C1_Z_3), .CI(
        DP_OP_113J3_124_6892_n7), .CO(DP_OP_113J3_124_6892_n6), .S(C81_DATA2_3) );
  fad1_hd DP_OP_113J3_124_6892_U10 ( .A(n1007), .B(C1_Z_2), .CI(
        DP_OP_113J3_124_6892_n8), .CO(DP_OP_113J3_124_6892_n7), .S(C81_DATA2_2) );
  fad1_hd DP_OP_113J3_124_6892_U11 ( .A(n1007), .B(C1_Z_1), .CI(n768), .CO(
        DP_OP_113J3_124_6892_n8), .S(C81_DATA2_1) );
  had1_hd DP_OP_125J3_130_6300_U32 ( .A(b_e[0]), .B(a_e[0]), .CO(
        DP_OP_125J3_130_6300_n20), .S(DP_OP_125J3_130_6300_n34) );
  fad1_hd DP_OP_125J3_130_6300_U31 ( .A(a_e[1]), .B(b_e[1]), .CI(
        DP_OP_125J3_130_6300_n20), .CO(DP_OP_125J3_130_6300_n19), .S(
        DP_OP_125J3_130_6300_n35) );
  fad1_hd DP_OP_125J3_130_6300_U30 ( .A(a_e[2]), .B(b_e[2]), .CI(
        DP_OP_125J3_130_6300_n19), .CO(DP_OP_125J3_130_6300_n18), .S(
        DP_OP_125J3_130_6300_n36) );
  fad1_hd DP_OP_125J3_130_6300_U29 ( .A(a_e[3]), .B(b_e[3]), .CI(
        DP_OP_125J3_130_6300_n18), .CO(DP_OP_125J3_130_6300_n17), .S(
        DP_OP_125J3_130_6300_n37) );
  fad1_hd DP_OP_125J3_130_6300_U28 ( .A(a_e[4]), .B(b_e[4]), .CI(
        DP_OP_125J3_130_6300_n17), .CO(DP_OP_125J3_130_6300_n16), .S(
        DP_OP_125J3_130_6300_n38) );
  fad1_hd DP_OP_125J3_130_6300_U27 ( .A(a_e[5]), .B(b_e[5]), .CI(
        DP_OP_125J3_130_6300_n16), .CO(DP_OP_125J3_130_6300_n15), .S(
        DP_OP_125J3_130_6300_n39) );
  fad1_hd DP_OP_125J3_130_6300_U26 ( .A(a_e[6]), .B(b_e[6]), .CI(
        DP_OP_125J3_130_6300_n15), .CO(DP_OP_125J3_130_6300_n14), .S(
        DP_OP_125J3_130_6300_n40) );
  fad1_hd DP_OP_125J3_130_6300_U25 ( .A(a_e[7]), .B(b_e[7]), .CI(
        DP_OP_125J3_130_6300_n14), .CO(DP_OP_125J3_130_6300_n13), .S(
        DP_OP_125J3_130_6300_n41) );
  fad1_hd DP_OP_125J3_130_6300_U24 ( .A(a_e[8]), .B(b_e[8]), .CI(
        DP_OP_125J3_130_6300_n13), .CO(DP_OP_125J3_130_6300_n12), .S(
        DP_OP_125J3_130_6300_n42) );
  fds2d1_hd a_e_reg_7_ ( .CRN(n141), .D(n138), .CK(i_CLK), .Q(n10), .QN(a_e[7]) );
  fds2d1_hd b_e_reg_7_ ( .CRN(n151), .D(n148), .CK(i_CLK), .Q(n14), .QN(b_e[7]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n359), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1023), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1023), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n1023), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n1023), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n1023), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n1023), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1023), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1023), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1023), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1023), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1023), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n1023), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n1023), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n359), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n359), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n359), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n359), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n359), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n1023), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1023), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n1023), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n1023), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n1023), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1023), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1023), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1023), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1023), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1023), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1023), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1023), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1023), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd product_reg_27_ ( .D(n1138), .E(n1010), .CK(i_CLK), .Q(
        product[27]) );
  fd1eqd1_hd product_reg_28_ ( .D(n1137), .E(n1010), .CK(i_CLK), .Q(
        product[28]) );
  fd1eqd1_hd product_reg_30_ ( .D(n1132), .E(n1010), .CK(i_CLK), .Q(
        product[30]) );
  fd1eqd1_hd product_reg_32_ ( .D(N206), .E(n1010), .CK(i_CLK), .Q(product[32]) );
  fd1eqd1_hd product_reg_34_ ( .D(N208), .E(n1010), .CK(i_CLK), .Q(product[34]) );
  fd1eqd1_hd product_reg_36_ ( .D(N210), .E(n1010), .CK(i_CLK), .Q(product[36]) );
  fd1eqd1_hd product_reg_38_ ( .D(N212), .E(n1010), .CK(i_CLK), .Q(product[38]) );
  fd1eqd1_hd product_reg_40_ ( .D(N214), .E(n1010), .CK(i_CLK), .Q(product[40]) );
  fd1eqd1_hd product_reg_42_ ( .D(N216), .E(n1010), .CK(i_CLK), .Q(product[42]) );
  fd1eqd1_hd product_reg_44_ ( .D(N218), .E(n1010), .CK(i_CLK), .Q(product[44]) );
  fd1eqd1_hd product_reg_46_ ( .D(N220), .E(n1010), .CK(i_CLK), .Q(product[46]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n2022), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n2022), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n2022), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n2022), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd product_reg_24_ ( .D(n1142), .E(n1010), .CK(i_CLK), .Q(
        product[24]) );
  fd1eqd1_hd product_reg_26_ ( .D(n1139), .E(n1010), .CK(i_CLK), .Q(
        product[26]) );
  fd1eqd1_hd product_reg_29_ ( .D(n1135), .E(n1010), .CK(i_CLK), .Q(
        product[29]) );
  fd1eqd1_hd product_reg_31_ ( .D(N205), .E(n1010), .CK(i_CLK), .Q(product[31]) );
  fd1eqd1_hd product_reg_33_ ( .D(N207), .E(n1010), .CK(i_CLK), .Q(product[33]) );
  fd1eqd1_hd product_reg_35_ ( .D(N209), .E(n1010), .CK(i_CLK), .Q(product[35]) );
  fd1eqd1_hd product_reg_37_ ( .D(N211), .E(n1010), .CK(i_CLK), .Q(product[37]) );
  fd1eqd1_hd product_reg_39_ ( .D(N213), .E(n1010), .CK(i_CLK), .Q(product[39]) );
  fd1eqd1_hd product_reg_41_ ( .D(N215), .E(n1010), .CK(i_CLK), .Q(product[41]) );
  fd1eqd1_hd product_reg_43_ ( .D(N217), .E(n1010), .CK(i_CLK), .Q(product[43]) );
  fd1eqd1_hd product_reg_45_ ( .D(N219), .E(n1010), .CK(i_CLK), .Q(product[45]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n2022), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n2022), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n2022), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n2022), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n2022), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n2022), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n2022), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n2022), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n2022), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n2022), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n2022), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n2022), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n2022), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n2022), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n2022), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n2022), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n2022), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n2022), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n2022), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n2022), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n2022), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n2022), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n2022), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n2022), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n2022), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n2022), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n2022), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n2022), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n2022), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n2022), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n2022), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n2022), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n2022), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n2022), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n2022), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n2022), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n2022), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n2022), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n2022), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n2022), .CK(i_CLK), .Q(b[22]) );
  fd1eqd1_hd product_reg_47_ ( .D(N221), .E(n1010), .CK(i_CLK), .Q(product[47]) );
  fd1eqd1_hd product_reg_48_ ( .D(N222), .E(n1010), .CK(i_CLK), .Q(product[48]) );
  fd1eqd1_hd product_reg_49_ ( .D(N223), .E(n1010), .CK(i_CLK), .Q(product[49]) );
  fd1eqd1_hd z_s_reg ( .D(N35), .E(n1010), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd product_reg_25_ ( .D(n1141), .E(n1010), .CK(i_CLK), .Q(
        product[25]) );
  fd1eqd1_hd product_reg_9_ ( .D(n1164), .E(n1010), .CK(i_CLK), .Q(product[9])
         );
  fd1eqd1_hd product_reg_20_ ( .D(n1148), .E(n1010), .CK(i_CLK), .Q(
        product[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n241), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n242), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_17_ ( .D(n243), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n244), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_15_ ( .D(n245), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n246), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_13_ ( .D(n247), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n248), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_11_ ( .D(n249), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n250), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_9_ ( .D(n251), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_3_ ( .D(n257), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_2_ ( .D(n258), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_1_ ( .D(n259), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_0_ ( .D(n260), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_21_ ( .D(n239), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n240), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_29_ ( .D(n231), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n233), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n235), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1120), .CK(i_CLK), .Q(a_s) );
  fd1eqd1_hd product_reg_5_ ( .D(N179), .E(n1010), .CK(i_CLK), .Q(product[5])
         );
  fd1eqd1_hd product_reg_10_ ( .D(n1162), .E(n1010), .CK(i_CLK), .Q(
        product[10]) );
  fd1eqd1_hd product_reg_18_ ( .D(n1151), .E(n1010), .CK(i_CLK), .Q(
        product[18]) );
  fd1eqd1_hd product_reg_19_ ( .D(n1149), .E(n1010), .CK(i_CLK), .Q(
        product[19]) );
  fd1eqd1_hd product_reg_23_ ( .D(n1143), .E(n1010), .CK(i_CLK), .Q(
        product[23]) );
  fd1eqd1_hd product_reg_4_ ( .D(N178), .E(n1010), .CK(i_CLK), .Q(product[4])
         );
  fd1eqd1_hd product_reg_7_ ( .D(n1166), .E(n1010), .CK(i_CLK), .Q(product[7])
         );
  fd1eqd1_hd product_reg_11_ ( .D(n1161), .E(n1010), .CK(i_CLK), .Q(
        product[11]) );
  fd1eqd1_hd product_reg_21_ ( .D(n1147), .E(n1010), .CK(i_CLK), .Q(
        product[21]) );
  fd1eqd1_hd product_reg_22_ ( .D(n1145), .E(n1010), .CK(i_CLK), .Q(
        product[22]) );
  fd1eqd1_hd product_reg_2_ ( .D(N176), .E(n1010), .CK(i_CLK), .Q(product[2])
         );
  fd1eqd1_hd product_reg_6_ ( .D(n1168), .E(n1010), .CK(i_CLK), .Q(product[6])
         );
  fd1eqd1_hd product_reg_15_ ( .D(n1156), .E(n1010), .CK(i_CLK), .Q(
        product[15]) );
  fd1eqd1_hd product_reg_16_ ( .D(n1154), .E(n1010), .CK(i_CLK), .Q(
        product[16]) );
  fd1eqd1_hd product_reg_17_ ( .D(n1152), .E(n1010), .CK(i_CLK), .Q(
        product[17]) );
  fd1eqd1_hd product_reg_3_ ( .D(N177), .E(n1010), .CK(i_CLK), .Q(product[3])
         );
  fd1eqd1_hd product_reg_8_ ( .D(n1165), .E(n1010), .CK(i_CLK), .Q(product[8])
         );
  fd1eqd1_hd product_reg_12_ ( .D(n1160), .E(n1010), .CK(i_CLK), .Q(
        product[12]) );
  fd1eqd1_hd product_reg_13_ ( .D(n1158), .E(n1010), .CK(i_CLK), .Q(
        product[13]) );
  fd1eqd1_hd product_reg_14_ ( .D(n1157), .E(n1010), .CK(i_CLK), .Q(
        product[14]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1120), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n2022), .CK(i_CLK), .Q(b[30]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n262), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n261), .CK(i_CLK), .Q(z_m[22]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n263), .CK(i_CLK), .Q(z_m[20]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n264), .CK(i_CLK), .Q(z_m[19]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n2022), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n2022), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n2022), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n2022), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n2022), .CK(i_CLK), .Q(b[28]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n2022), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd guard_reg ( .D(n104), .E(n105), .CK(i_CLK), .Q(net922) );
  fd1qd1_hd z_m_reg_16_ ( .D(n267), .CK(i_CLK), .Q(z_m[16]) );
  fd1qd1_hd z_m_reg_14_ ( .D(n269), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n265), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n320), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n311), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n270), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n266), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n268), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n319), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n356), .CK(i_CLK), .Q(b_e[9]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n2022), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n2022), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n2022), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n2022), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n2022), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n2022), .CK(i_CLK), .Q(b[26]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n2022), .CK(i_CLK), .Q(b[23]) );
  fd1eqd1_hd z_e_reg_8_ ( .D(N474), .E(n110), .CK(i_CLK), .Q(z_e[8]) );
  fd1eqd1_hd z_e_reg_9_ ( .D(N475), .E(n110), .CK(i_CLK), .Q(z_e[9]) );
  fd1eqd1_hd z_e_reg_2_ ( .D(N468), .E(n110), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n286), .CK(i_CLK), .Q(z_m[23]) );
  fd1eqd1_hd z_e_reg_7_ ( .D(N473), .E(n110), .CK(i_CLK), .Q(z_e[7]) );
  fd1eqd1_hd z_e_reg_1_ ( .D(N467), .E(n110), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n323), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n314), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n322), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n321), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n313), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n312), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n275), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n271), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n273), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n274), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n276), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n272), .CK(i_CLK), .Q(z_m[11]) );
  fd1eqd1_hd z_e_reg_4_ ( .D(N470), .E(n110), .CK(i_CLK), .Q(z_e[4]) );
  fd1eqd1_hd z_e_reg_6_ ( .D(N472), .E(n110), .CK(i_CLK), .Q(z_e[6]) );
  fd1eqd1_hd z_e_reg_3_ ( .D(N469), .E(n110), .CK(i_CLK), .Q(z_e[3]) );
  fd1eqd1_hd z_e_reg_5_ ( .D(N471), .E(n110), .CK(i_CLK), .Q(z_e[5]) );
  fd1eqd1_hd z_e_reg_0_ ( .D(n1004), .E(n110), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n325), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n281), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n324), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n316), .CK(i_CLK), .Q(a_e[2]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n315), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n282), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n279), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n277), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n326), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n317), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n278), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n280), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n327), .CK(i_CLK), .Q(b_e[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n318), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd state_reg_3_ ( .D(n357), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd state_reg_0_ ( .D(n353), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd state_reg_2_ ( .D(n351), .CK(i_CLK), .Q(state[2]) );
  fad1_hd DP_OP_125J3_130_6300_U10 ( .A(n1106), .B(n1112), .CI(
        DP_OP_125J3_130_6300_n25), .CO(DP_OP_125J3_130_6300_n9), .S(N467) );
  ivd1_hd U511 ( .A(N34), .Y(n1005) );
  fad1_hd intadd_26_U18 ( .A(intadd_26_A_0_), .B(intadd_26_B_0_), .CI(
        intadd_26_CI), .CO(intadd_26_n17), .S(intadd_26_SUM_0_) );
  fad1_hd intadd_26_U17 ( .A(intadd_26_A_1_), .B(intadd_26_B_1_), .CI(
        intadd_26_n17), .CO(intadd_26_n16), .S(intadd_26_SUM_1_) );
  fad1_hd intadd_26_U16 ( .A(intadd_26_A_2_), .B(intadd_26_B_2_), .CI(
        intadd_26_n16), .CO(intadd_26_n15), .S(intadd_26_SUM_2_) );
  fad1_hd intadd_26_U15 ( .A(intadd_26_A_3_), .B(intadd_26_B_3_), .CI(
        intadd_26_n15), .CO(intadd_26_n14), .S(intadd_26_SUM_3_) );
  fad1_hd intadd_26_U14 ( .A(intadd_26_A_4_), .B(intadd_26_B_4_), .CI(
        intadd_26_n14), .CO(intadd_26_n13), .S(intadd_26_SUM_4_) );
  fad1_hd intadd_26_U13 ( .A(intadd_26_A_5_), .B(intadd_26_B_5_), .CI(
        intadd_26_n13), .CO(intadd_26_n12), .S(intadd_26_SUM_5_) );
  fad1_hd intadd_26_U12 ( .A(intadd_26_A_6_), .B(intadd_26_B_6_), .CI(
        intadd_26_n12), .CO(intadd_26_n11), .S(intadd_26_SUM_6_) );
  fad1_hd intadd_26_U11 ( .A(intadd_26_A_7_), .B(intadd_26_B_7_), .CI(
        intadd_26_n11), .CO(intadd_26_n10), .S(intadd_26_SUM_7_) );
  fad1_hd intadd_26_U10 ( .A(intadd_26_A_8_), .B(intadd_26_B_8_), .CI(
        intadd_26_n10), .CO(intadd_26_n9), .S(intadd_26_SUM_8_) );
  fad1_hd intadd_26_U9 ( .A(intadd_26_A_9_), .B(intadd_26_B_9_), .CI(
        intadd_26_n9), .CO(intadd_26_n8), .S(intadd_26_SUM_9_) );
  fad1_hd intadd_26_U8 ( .A(intadd_26_A_10_), .B(intadd_26_B_10_), .CI(
        intadd_26_n8), .CO(intadd_26_n7), .S(intadd_26_SUM_10_) );
  fad1_hd intadd_26_U7 ( .A(intadd_26_A_11_), .B(intadd_26_B_11_), .CI(
        intadd_26_n7), .CO(intadd_26_n6), .S(intadd_26_SUM_11_) );
  fad1_hd intadd_26_U6 ( .A(intadd_26_A_12_), .B(intadd_26_B_12_), .CI(
        intadd_26_n6), .CO(intadd_26_n5), .S(intadd_26_SUM_12_) );
  fad1_hd intadd_26_U5 ( .A(intadd_26_A_13_), .B(intadd_26_B_13_), .CI(
        intadd_26_n5), .CO(intadd_26_n4), .S(intadd_26_SUM_13_) );
  fad1_hd intadd_26_U4 ( .A(intadd_28_n1), .B(intadd_26_B_14_), .CI(
        intadd_26_n4), .CO(intadd_26_n3), .S(intadd_26_SUM_14_) );
  fad1_hd intadd_27_U15 ( .A(intadd_27_A_0_), .B(intadd_27_B_0_), .CI(
        intadd_27_CI), .CO(intadd_27_n14), .S(intadd_27_SUM_0_) );
  fad1_hd intadd_27_U14 ( .A(intadd_27_A_1_), .B(intadd_27_B_1_), .CI(
        intadd_27_n14), .CO(intadd_27_n13), .S(intadd_27_SUM_1_) );
  fad1_hd intadd_27_U13 ( .A(intadd_27_A_2_), .B(intadd_27_B_2_), .CI(
        intadd_27_n13), .CO(intadd_27_n12), .S(intadd_27_SUM_2_) );
  fad1_hd intadd_27_U12 ( .A(intadd_27_A_3_), .B(intadd_27_B_3_), .CI(
        intadd_27_n12), .CO(intadd_27_n11), .S(intadd_27_SUM_3_) );
  fad1_hd intadd_27_U11 ( .A(intadd_27_A_4_), .B(intadd_27_B_4_), .CI(
        intadd_27_n11), .CO(intadd_27_n10), .S(intadd_27_SUM_4_) );
  fad1_hd intadd_27_U10 ( .A(intadd_27_A_5_), .B(intadd_27_B_5_), .CI(
        intadd_27_n10), .CO(intadd_27_n9), .S(intadd_27_SUM_5_) );
  fad1_hd intadd_27_U9 ( .A(intadd_27_A_6_), .B(intadd_27_B_6_), .CI(
        intadd_27_n9), .CO(intadd_27_n8), .S(intadd_27_SUM_6_) );
  fad1_hd intadd_27_U8 ( .A(intadd_27_A_7_), .B(intadd_27_B_7_), .CI(
        intadd_27_n8), .CO(intadd_27_n7), .S(intadd_27_SUM_7_) );
  fad1_hd intadd_27_U7 ( .A(intadd_27_A_8_), .B(intadd_27_B_8_), .CI(
        intadd_27_n7), .CO(intadd_27_n6), .S(intadd_27_SUM_8_) );
  fad1_hd intadd_27_U6 ( .A(intadd_27_A_9_), .B(intadd_27_B_9_), .CI(
        intadd_27_n6), .CO(intadd_27_n5), .S(intadd_27_SUM_9_) );
  fad1_hd intadd_27_U5 ( .A(intadd_27_A_10_), .B(intadd_27_B_10_), .CI(
        intadd_27_n5), .CO(intadd_27_n4), .S(intadd_27_SUM_10_) );
  fad1_hd intadd_27_U4 ( .A(intadd_27_A_11_), .B(intadd_27_B_11_), .CI(
        intadd_27_n4), .CO(intadd_27_n3), .S(intadd_27_SUM_11_) );
  fad1_hd intadd_27_U3 ( .A(intadd_29_n1), .B(intadd_27_B_12_), .CI(
        intadd_27_n3), .CO(intadd_27_n2), .S(intadd_27_SUM_12_) );
  fad1_hd intadd_27_U2 ( .A(intadd_27_A_13_), .B(intadd_27_B_13_), .CI(
        intadd_27_n2), .CO(intadd_27_n1), .S(intadd_27_SUM_13_) );
  fad1_hd intadd_28_U12 ( .A(intadd_28_A_0_), .B(intadd_28_B_0_), .CI(
        intadd_28_CI), .CO(intadd_28_n11), .S(intadd_26_B_3_) );
  fad1_hd intadd_28_U11 ( .A(intadd_28_A_1_), .B(intadd_28_B_1_), .CI(
        intadd_28_n11), .CO(intadd_28_n10), .S(intadd_26_B_4_) );
  fad1_hd intadd_28_U10 ( .A(intadd_28_A_2_), .B(intadd_28_B_2_), .CI(
        intadd_28_n10), .CO(intadd_28_n9), .S(intadd_26_B_5_) );
  fad1_hd intadd_28_U9 ( .A(intadd_28_A_3_), .B(intadd_27_SUM_0_), .CI(
        intadd_28_n9), .CO(intadd_28_n8), .S(intadd_26_B_6_) );
  fad1_hd intadd_28_U8 ( .A(intadd_28_A_4_), .B(intadd_27_SUM_1_), .CI(
        intadd_28_n8), .CO(intadd_28_n7), .S(intadd_26_B_7_) );
  fad1_hd intadd_28_U7 ( .A(intadd_28_A_5_), .B(intadd_27_SUM_2_), .CI(
        intadd_28_n7), .CO(intadd_28_n6), .S(intadd_26_A_8_) );
  fad1_hd intadd_28_U6 ( .A(intadd_28_A_6_), .B(intadd_27_SUM_3_), .CI(
        intadd_28_n6), .CO(intadd_28_n5), .S(intadd_26_B_9_) );
  fad1_hd intadd_28_U5 ( .A(intadd_28_A_7_), .B(intadd_27_SUM_4_), .CI(
        intadd_28_n5), .CO(intadd_28_n4), .S(intadd_26_A_10_) );
  fad1_hd intadd_28_U4 ( .A(intadd_28_A_8_), .B(intadd_27_SUM_5_), .CI(
        intadd_28_n4), .CO(intadd_28_n3), .S(intadd_26_B_11_) );
  fad1_hd intadd_28_U3 ( .A(intadd_27_SUM_6_), .B(intadd_28_B_9_), .CI(
        intadd_28_n3), .CO(intadd_28_n2), .S(intadd_26_A_12_) );
  fad1_hd intadd_28_U2 ( .A(intadd_28_A_10_), .B(intadd_27_SUM_7_), .CI(
        intadd_28_n2), .CO(intadd_28_n1), .S(intadd_26_B_13_) );
  fad1_hd intadd_29_U10 ( .A(intadd_29_A_0_), .B(intadd_29_B_0_), .CI(
        intadd_29_CI), .CO(intadd_29_n9), .S(intadd_27_B_3_) );
  fad1_hd intadd_29_U9 ( .A(intadd_29_A_1_), .B(intadd_29_B_1_), .CI(
        intadd_29_n9), .CO(intadd_29_n8), .S(intadd_27_B_4_) );
  fad1_hd intadd_29_U8 ( .A(intadd_29_A_2_), .B(intadd_29_B_2_), .CI(
        intadd_29_n8), .CO(intadd_29_n7), .S(intadd_27_B_5_) );
  fad1_hd intadd_29_U7 ( .A(n2027), .B(intadd_29_B_3_), .CI(intadd_29_n7), 
        .CO(intadd_29_n6), .S(intadd_27_A_6_) );
  fad1_hd intadd_29_U6 ( .A(intadd_29_A_4_), .B(n2026), .CI(intadd_29_n6), 
        .CO(intadd_29_n5), .S(intadd_27_B_7_) );
  fad1_hd intadd_29_U5 ( .A(n2025), .B(intadd_29_B_5_), .CI(intadd_29_n5), 
        .CO(intadd_29_n4), .S(intadd_27_B_8_) );
  fad1_hd intadd_29_U4 ( .A(n1215), .B(intadd_29_B_6_), .CI(intadd_29_n4), 
        .CO(intadd_29_n3), .S(intadd_27_A_9_) );
  fad1_hd intadd_29_U3 ( .A(n1212), .B(intadd_29_B_7_), .CI(intadd_29_n3), 
        .CO(intadd_29_n2), .S(intadd_27_B_10_) );
  fad1_hd intadd_29_U2 ( .A(n1206), .B(intadd_29_B_8_), .CI(intadd_29_n2), 
        .CO(intadd_29_n1), .S(intadd_27_A_11_) );
  fad1_hd intadd_31_U9 ( .A(a_m[5]), .B(a_m[2]), .CI(intadd_31_CI), .CO(
        intadd_31_n8), .S(intadd_31_SUM_0_) );
  fad1_hd intadd_31_U8 ( .A(n1225), .B(intadd_31_B_1_), .CI(intadd_31_n8), 
        .CO(intadd_31_n7), .S(intadd_31_SUM_1_) );
  fad1_hd intadd_31_U7 ( .A(intadd_31_A_2_), .B(intadd_31_B_2_), .CI(
        intadd_31_n7), .CO(intadd_31_n6), .S(intadd_31_SUM_2_) );
  fad1_hd intadd_31_U6 ( .A(intadd_31_A_3_), .B(intadd_31_B_3_), .CI(
        intadd_31_n6), .CO(intadd_31_n5), .S(intadd_31_SUM_3_) );
  fad1_hd intadd_31_U5 ( .A(intadd_31_A_4_), .B(intadd_31_B_4_), .CI(
        intadd_31_n5), .CO(intadd_31_n4), .S(intadd_31_SUM_4_) );
  fad1_hd intadd_31_U4 ( .A(intadd_31_A_5_), .B(n1210), .CI(intadd_31_n4), 
        .CO(intadd_31_n3), .S(intadd_31_SUM_5_) );
  fad1_hd intadd_31_U3 ( .A(n1208), .B(intadd_31_B_6_), .CI(intadd_31_n3), 
        .CO(intadd_31_n2), .S(intadd_31_SUM_6_) );
  fad1_hd intadd_31_U2 ( .A(n1201), .B(intadd_31_B_7_), .CI(intadd_31_n2), 
        .CO(intadd_31_n1), .S(intadd_31_SUM_7_) );
  fad1_hd intadd_32_U7 ( .A(n1222), .B(intadd_32_B_0_), .CI(intadd_32_CI), 
        .CO(intadd_32_n6), .S(intadd_32_SUM_0_) );
  fad1_hd intadd_32_U6 ( .A(intadd_32_A_1_), .B(intadd_32_B_1_), .CI(
        intadd_32_n6), .CO(intadd_32_n5), .S(intadd_32_SUM_1_) );
  fad1_hd intadd_32_U5 ( .A(intadd_32_A_2_), .B(intadd_32_B_2_), .CI(
        intadd_32_n5), .CO(intadd_32_n4), .S(intadd_32_SUM_2_) );
  fad1_hd intadd_32_U4 ( .A(intadd_32_A_3_), .B(intadd_32_B_3_), .CI(
        intadd_32_n4), .CO(intadd_32_n3), .S(intadd_32_SUM_3_) );
  fad1_hd intadd_32_U3 ( .A(intadd_32_A_4_), .B(n1198), .CI(intadd_32_n3), 
        .CO(intadd_32_n2), .S(intadd_32_SUM_4_) );
  fad1_hd intadd_33_U6 ( .A(n2039), .B(intadd_33_B_0_), .CI(intadd_33_CI), 
        .CO(intadd_33_n5), .S(intadd_33_SUM_0_) );
  fad1_hd intadd_33_U5 ( .A(intadd_33_A_1_), .B(intadd_33_B_1_), .CI(
        intadd_33_n5), .CO(intadd_33_n4), .S(intadd_33_SUM_1_) );
  fad1_hd intadd_33_U4 ( .A(n1204), .B(intadd_33_B_2_), .CI(intadd_33_n4), 
        .CO(intadd_33_n3), .S(intadd_33_SUM_2_) );
  fad1_hd intadd_33_U3 ( .A(n1191), .B(n1197), .CI(intadd_33_n3), .CO(
        intadd_33_n2), .S(intadd_33_SUM_3_) );
  fad1_hd intadd_34_U4 ( .A(intadd_34_A_0_), .B(intadd_34_B_0_), .CI(
        intadd_34_CI), .CO(intadd_34_n3), .S(intadd_34_SUM_0_) );
  fad1_hd intadd_34_U3 ( .A(intadd_34_A_1_), .B(intadd_34_B_1_), .CI(
        intadd_34_n3), .CO(intadd_34_n2), .S(intadd_34_SUM_1_) );
  fad1_hd intadd_35_U4 ( .A(a_m[2]), .B(intadd_35_B_0_), .CI(intadd_35_CI), 
        .CO(intadd_35_n3), .S(intadd_35_SUM_0_) );
  fad1_hd intadd_35_U3 ( .A(intadd_35_A_1_), .B(n1224), .CI(intadd_35_n3), 
        .CO(intadd_35_n2), .S(intadd_35_SUM_1_) );
  fad1_hd intadd_35_U2 ( .A(n1213), .B(intadd_35_B_2_), .CI(intadd_35_n2), 
        .CO(intadd_35_n1), .S(intadd_35_SUM_2_) );
  fad1_hd intadd_36_U3 ( .A(intadd_36_A_1_), .B(intadd_36_B_1_), .CI(
        intadd_36_n3), .CO(intadd_36_n2), .S(intadd_36_SUM_1_) );
  fad1_hd intadd_36_U2 ( .A(intadd_36_A_2_), .B(intadd_36_B_2_), .CI(
        intadd_36_n2), .CO(intadd_36_n1), .S(intadd_36_SUM_2_) );
  fad1_hd intadd_37_U4 ( .A(intadd_37_A_0_), .B(intadd_37_B_0_), .CI(
        intadd_32_SUM_1_), .CO(intadd_37_n3), .S(intadd_37_SUM_0_) );
  fad1_hd intadd_37_U3 ( .A(intadd_32_SUM_2_), .B(intadd_37_B_1_), .CI(
        intadd_37_n3), .CO(intadd_37_n2), .S(intadd_37_SUM_1_) );
  fad1_hd intadd_38_U4 ( .A(intadd_31_SUM_5_), .B(intadd_38_B_0_), .CI(
        intadd_38_CI), .CO(intadd_38_n3), .S(intadd_38_SUM_0_) );
  fad1_hd intadd_38_U3 ( .A(intadd_31_SUM_6_), .B(intadd_38_B_1_), .CI(
        intadd_38_n3), .CO(intadd_38_n2), .S(intadd_38_SUM_1_) );
  fad1_hd intadd_39_U4 ( .A(n1205), .B(intadd_39_B_0_), .CI(intadd_39_CI), 
        .CO(intadd_39_n3), .S(intadd_27_B_12_) );
  fad1_hd intadd_39_U3 ( .A(n1203), .B(intadd_39_B_1_), .CI(intadd_39_n3), 
        .CO(intadd_39_n2), .S(intadd_27_A_13_) );
  fad1_hd intadd_40_U4 ( .A(intadd_31_SUM_2_), .B(intadd_40_B_0_), .CI(
        intadd_40_CI), .CO(intadd_40_n3), .S(intadd_40_SUM_0_) );
  fad1_hd intadd_40_U3 ( .A(intadd_31_SUM_3_), .B(intadd_40_B_1_), .CI(
        intadd_40_n3), .CO(intadd_40_n2), .S(intadd_40_SUM_1_) );
  fad1_hd intadd_40_U2 ( .A(intadd_31_SUM_4_), .B(intadd_40_B_2_), .CI(
        intadd_40_n2), .CO(intadd_40_n1), .S(intadd_40_SUM_2_) );
  fad1_hd intadd_41_U4 ( .A(intadd_41_A_0_), .B(intadd_27_SUM_9_), .CI(
        intadd_41_CI), .CO(intadd_41_n3), .S(intadd_26_A_15_) );
  fad1_hd intadd_41_U3 ( .A(intadd_41_A_1_), .B(intadd_27_SUM_10_), .CI(
        intadd_41_n3), .CO(intadd_41_n2), .S(intadd_26_A_16_) );
  fad1_hd intadd_21_U26 ( .A(intadd_21_A_0_), .B(intadd_21_B_0_), .CI(
        intadd_21_CI), .CO(intadd_21_n25), .S(intadd_21_SUM_0_) );
  fad1_hd intadd_21_U25 ( .A(intadd_21_A_1_), .B(intadd_21_B_1_), .CI(
        intadd_21_n25), .CO(intadd_21_n24), .S(intadd_21_SUM_1_) );
  fad1_hd intadd_21_U24 ( .A(intadd_21_A_2_), .B(intadd_21_B_2_), .CI(
        intadd_21_n24), .CO(intadd_21_n23), .S(intadd_21_SUM_2_) );
  fad1_hd intadd_21_U23 ( .A(intadd_21_A_3_), .B(intadd_21_B_3_), .CI(
        intadd_21_n23), .CO(intadd_21_n22), .S(intadd_21_SUM_3_) );
  fad1_hd intadd_21_U22 ( .A(intadd_21_A_4_), .B(intadd_21_B_4_), .CI(
        intadd_21_n22), .CO(intadd_21_n21), .S(intadd_21_SUM_4_) );
  fad1_hd intadd_21_U21 ( .A(intadd_21_A_5_), .B(intadd_21_B_5_), .CI(
        intadd_21_n21), .CO(intadd_21_n20), .S(intadd_21_SUM_5_) );
  fad1_hd intadd_21_U20 ( .A(intadd_21_A_6_), .B(intadd_21_B_6_), .CI(
        intadd_21_n20), .CO(intadd_21_n19), .S(intadd_21_SUM_6_) );
  fad1_hd intadd_21_U19 ( .A(intadd_21_A_7_), .B(intadd_21_B_7_), .CI(
        intadd_21_n19), .CO(intadd_21_n18), .S(intadd_21_SUM_7_) );
  fad1_hd intadd_21_U18 ( .A(intadd_21_A_8_), .B(intadd_21_B_8_), .CI(
        intadd_21_n18), .CO(intadd_21_n17), .S(intadd_21_SUM_8_) );
  fad1_hd intadd_21_U17 ( .A(intadd_21_A_9_), .B(intadd_21_B_9_), .CI(
        intadd_21_n17), .CO(intadd_21_n16), .S(intadd_21_SUM_9_) );
  fad1_hd intadd_21_U16 ( .A(intadd_21_A_10_), .B(intadd_21_B_10_), .CI(
        intadd_21_n16), .CO(intadd_21_n15), .S(intadd_21_SUM_10_) );
  fad1_hd intadd_21_U15 ( .A(intadd_21_A_11_), .B(intadd_21_B_11_), .CI(
        intadd_21_n15), .CO(intadd_21_n14), .S(intadd_21_SUM_11_) );
  fad1_hd intadd_21_U14 ( .A(intadd_21_A_12_), .B(intadd_21_B_12_), .CI(
        intadd_21_n14), .CO(intadd_21_n13), .S(intadd_21_SUM_12_) );
  fad1_hd intadd_21_U13 ( .A(intadd_21_A_13_), .B(intadd_21_B_13_), .CI(
        intadd_21_n13), .CO(intadd_21_n12), .S(intadd_21_SUM_13_) );
  fad1_hd intadd_21_U12 ( .A(intadd_21_A_14_), .B(intadd_21_B_14_), .CI(
        intadd_21_n12), .CO(intadd_21_n11), .S(intadd_21_SUM_14_) );
  fad1_hd intadd_21_U11 ( .A(intadd_21_A_15_), .B(intadd_21_B_15_), .CI(
        intadd_21_n11), .CO(intadd_21_n10), .S(intadd_21_SUM_15_) );
  fad1_hd intadd_21_U10 ( .A(intadd_21_A_16_), .B(intadd_21_B_16_), .CI(
        intadd_21_n10), .CO(intadd_21_n9), .S(intadd_21_SUM_16_) );
  fad1_hd intadd_21_U9 ( .A(intadd_21_A_17_), .B(intadd_21_B_17_), .CI(
        intadd_21_n9), .CO(intadd_21_n8), .S(intadd_21_SUM_17_) );
  fad1_hd intadd_21_U8 ( .A(intadd_21_A_18_), .B(intadd_21_B_18_), .CI(
        intadd_21_n8), .CO(intadd_21_n7), .S(intadd_21_SUM_18_) );
  fad1_hd intadd_21_U7 ( .A(intadd_21_A_19_), .B(intadd_21_B_19_), .CI(
        intadd_21_n7), .CO(intadd_21_n6), .S(intadd_21_SUM_19_) );
  fad1_hd intadd_22_U21 ( .A(a_m[2]), .B(intadd_22_B_0_), .CI(intadd_22_CI), 
        .CO(intadd_22_n20), .S(intadd_22_SUM_0_) );
  fad1_hd intadd_22_U20 ( .A(n2038), .B(intadd_35_SUM_0_), .CI(intadd_22_n20), 
        .CO(intadd_22_n19), .S(intadd_22_SUM_1_) );
  fad1_hd intadd_22_U19 ( .A(intadd_35_SUM_1_), .B(intadd_22_B_2_), .CI(
        intadd_22_n19), .CO(intadd_22_n18), .S(intadd_22_SUM_2_) );
  fad1_hd intadd_22_U18 ( .A(intadd_35_SUM_2_), .B(intadd_22_B_3_), .CI(
        intadd_22_n18), .CO(intadd_22_n17), .S(intadd_22_SUM_3_) );
  fad1_hd intadd_22_U17 ( .A(intadd_35_n1), .B(n1209), .CI(intadd_22_n17), 
        .CO(intadd_22_n16), .S(intadd_22_SUM_4_) );
  fad1_hd intadd_22_U16 ( .A(n1207), .B(intadd_22_B_5_), .CI(intadd_22_n16), 
        .CO(intadd_22_n15), .S(intadd_22_SUM_5_) );
  fad1_hd intadd_22_U15 ( .A(n1200), .B(intadd_22_B_6_), .CI(intadd_22_n15), 
        .CO(intadd_22_n14), .S(intadd_22_SUM_6_) );
  fad1_hd intadd_22_U14 ( .A(n1199), .B(n1196), .CI(intadd_22_n14), .CO(
        intadd_22_n13), .S(intadd_22_SUM_7_) );
  fad1_hd intadd_23_U20 ( .A(intadd_23_A_0_), .B(intadd_23_B_0_), .CI(
        intadd_23_CI), .CO(intadd_23_n19), .S(intadd_21_A_3_) );
  fad1_hd intadd_23_U19 ( .A(intadd_23_A_1_), .B(intadd_23_B_1_), .CI(
        intadd_23_n19), .CO(intadd_23_n18), .S(intadd_21_A_4_) );
  fad1_hd intadd_23_U16 ( .A(intadd_23_A_4_), .B(intadd_23_B_4_), .CI(
        intadd_23_n16), .CO(intadd_23_n15), .S(intadd_21_A_7_) );
  fad1_hd intadd_23_U15 ( .A(intadd_23_A_5_), .B(intadd_23_B_5_), .CI(
        intadd_23_n15), .CO(intadd_23_n14), .S(intadd_21_A_8_) );
  fad1_hd intadd_23_U14 ( .A(intadd_23_A_6_), .B(intadd_23_B_6_), .CI(
        intadd_23_n14), .CO(intadd_23_n13), .S(intadd_21_A_9_) );
  fad1_hd intadd_23_U13 ( .A(intadd_23_A_7_), .B(intadd_23_B_7_), .CI(
        intadd_23_n13), .CO(intadd_23_n12), .S(intadd_21_A_10_) );
  fad1_hd intadd_23_U12 ( .A(intadd_23_A_8_), .B(intadd_23_B_8_), .CI(
        intadd_23_n12), .CO(intadd_23_n11), .S(intadd_21_A_11_) );
  fad1_hd intadd_23_U11 ( .A(intadd_23_A_9_), .B(intadd_23_B_9_), .CI(
        intadd_23_n11), .CO(intadd_23_n10), .S(intadd_21_A_12_) );
  fad1_hd intadd_23_U10 ( .A(intadd_23_A_10_), .B(intadd_23_B_10_), .CI(
        intadd_23_n10), .CO(intadd_23_n9), .S(intadd_21_A_13_) );
  fad1_hd intadd_23_U9 ( .A(intadd_23_A_11_), .B(intadd_23_B_11_), .CI(
        intadd_23_n9), .CO(intadd_23_n8), .S(intadd_21_A_14_) );
  fad1_hd intadd_23_U8 ( .A(intadd_23_A_12_), .B(intadd_23_B_12_), .CI(
        intadd_23_n8), .CO(intadd_23_n7), .S(intadd_21_A_15_) );
  fad1_hd intadd_23_U7 ( .A(intadd_23_A_13_), .B(intadd_23_B_13_), .CI(
        intadd_23_n7), .CO(intadd_23_n6), .S(intadd_21_A_16_) );
  fad1_hd intadd_23_U6 ( .A(intadd_23_A_14_), .B(intadd_23_B_14_), .CI(
        intadd_23_n6), .CO(intadd_23_n5), .S(intadd_21_A_17_) );
  fad1_hd intadd_23_U5 ( .A(intadd_23_A_15_), .B(intadd_23_B_15_), .CI(
        intadd_23_n5), .CO(intadd_23_n4), .S(intadd_21_A_18_) );
  fad1_hd intadd_23_U4 ( .A(intadd_23_A_16_), .B(intadd_23_B_16_), .CI(
        intadd_23_n4), .CO(intadd_23_n3), .S(intadd_21_A_19_) );
  fad1_hd intadd_25_U18 ( .A(intadd_25_A_0_), .B(intadd_25_B_0_), .CI(
        intadd_25_CI), .CO(intadd_25_n17), .S(intadd_23_A_3_) );
  fad1_hd intadd_25_U17 ( .A(intadd_25_A_1_), .B(intadd_25_B_1_), .CI(
        intadd_25_n17), .CO(intadd_25_n16), .S(intadd_23_A_4_) );
  fad1_hd intadd_25_U16 ( .A(intadd_25_A_2_), .B(intadd_25_B_2_), .CI(
        intadd_25_n16), .CO(intadd_25_n15), .S(intadd_23_A_5_) );
  fad1_hd intadd_25_U15 ( .A(intadd_26_SUM_0_), .B(intadd_25_B_3_), .CI(
        intadd_25_n15), .CO(intadd_25_n14), .S(intadd_23_A_6_) );
  fad1_hd intadd_25_U14 ( .A(intadd_26_SUM_1_), .B(intadd_25_B_4_), .CI(
        intadd_25_n14), .CO(intadd_25_n13), .S(intadd_23_A_7_) );
  fad1_hd intadd_25_U13 ( .A(intadd_26_SUM_2_), .B(intadd_25_B_5_), .CI(
        intadd_25_n13), .CO(intadd_25_n12), .S(intadd_23_A_8_) );
  fad1_hd intadd_25_U12 ( .A(intadd_26_SUM_3_), .B(intadd_25_B_6_), .CI(
        intadd_25_n12), .CO(intadd_25_n11), .S(intadd_23_A_9_) );
  fad1_hd intadd_25_U11 ( .A(intadd_26_SUM_4_), .B(intadd_25_B_7_), .CI(
        intadd_25_n11), .CO(intadd_25_n10), .S(intadd_23_B_10_) );
  fad1_hd intadd_25_U10 ( .A(intadd_26_SUM_5_), .B(intadd_25_B_8_), .CI(
        intadd_25_n10), .CO(intadd_25_n9), .S(intadd_23_A_11_) );
  fad1_hd intadd_25_U9 ( .A(intadd_26_SUM_6_), .B(intadd_25_B_9_), .CI(
        intadd_25_n9), .CO(intadd_25_n8), .S(intadd_23_A_12_) );
  fad1_hd intadd_25_U8 ( .A(intadd_25_A_10_), .B(intadd_26_SUM_7_), .CI(
        intadd_25_n8), .CO(intadd_25_n7), .S(intadd_23_B_13_) );
  fad1_hd intadd_25_U7 ( .A(intadd_26_SUM_8_), .B(intadd_25_B_11_), .CI(
        intadd_25_n7), .CO(intadd_25_n6), .S(intadd_23_A_14_) );
  fad1_hd intadd_25_U6 ( .A(intadd_26_SUM_9_), .B(intadd_25_B_12_), .CI(
        intadd_25_n6), .CO(intadd_25_n5), .S(intadd_23_A_15_) );
  fad1_hd intadd_25_U5 ( .A(intadd_25_A_13_), .B(intadd_26_SUM_10_), .CI(
        intadd_25_n5), .CO(intadd_25_n4), .S(intadd_23_A_16_) );
  fad1_hd intadd_25_U4 ( .A(intadd_26_SUM_11_), .B(intadd_25_B_14_), .CI(
        intadd_25_n4), .CO(intadd_25_n3), .S(intadd_23_A_17_) );
  fad1_hd intadd_25_U3 ( .A(intadd_25_A_15_), .B(intadd_26_SUM_12_), .CI(
        intadd_25_n3), .CO(intadd_25_n2), .S(intadd_23_B_18_) );
  fad1_hd intadd_25_U2 ( .A(intadd_26_SUM_13_), .B(intadd_25_B_16_), .CI(
        intadd_25_n2), .CO(intadd_25_n1), .S(intadd_21_A_22_) );
  fad1_hd intadd_21_U5 ( .A(intadd_21_A_21_), .B(intadd_21_B_21_), .CI(
        intadd_21_n5), .CO(intadd_21_n4), .S(intadd_21_SUM_21_) );
  fad1_hd intadd_21_U6 ( .A(intadd_21_A_20_), .B(intadd_21_B_20_), .CI(
        intadd_21_n6), .CO(intadd_21_n5), .S(intadd_21_SUM_20_) );
  fad1_hd intadd_41_U2 ( .A(intadd_27_SUM_11_), .B(intadd_41_B_2_), .CI(
        intadd_41_n2), .CO(intadd_41_n1), .S(intadd_41_SUM_2_) );
  fad1_hd intadd_26_U3 ( .A(intadd_26_A_15_), .B(intadd_26_B_15_), .CI(
        intadd_26_n3), .CO(intadd_26_n2), .S(intadd_26_SUM_15_) );
  fad1_hd intadd_26_U2 ( .A(intadd_26_A_16_), .B(intadd_26_B_16_), .CI(
        intadd_26_n2), .CO(intadd_26_n1), .S(intadd_26_SUM_16_) );
  fad1_hd intadd_30_U9 ( .A(n1134), .B(intadd_30_B_0_), .CI(intadd_30_CI), 
        .CO(intadd_30_n8), .S(intadd_30_SUM_0_) );
  fad1_hd intadd_39_U2 ( .A(n1192), .B(intadd_39_B_2_), .CI(intadd_39_n2), 
        .CO(intadd_39_n1), .S(intadd_39_SUM_2_) );
  fad1_hd intadd_21_U4 ( .A(intadd_21_A_22_), .B(intadd_23_n1), .CI(
        intadd_21_n4), .CO(intadd_21_n3), .S(intadd_21_SUM_22_) );
  fd1qd1_hd o_Z_STB_reg ( .D(n358), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd a_m_reg_18_ ( .D(n331), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n334), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n337), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n340), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n252), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_7_ ( .D(n253), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n254), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_5_ ( .D(n255), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_4_ ( .D(n256), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd round_bit_reg ( .D(n284), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd b_m_reg_20_ ( .D(n288), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n290), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n291), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n294), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n296), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n300), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n302), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n303), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n287), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n309), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n289), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n292), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n293), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n295), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n297), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n298), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n299), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n301), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n304), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n305), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n306), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n307), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n349), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n354), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n328), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n330), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n333), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n336), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n339), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n342), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n345), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n348), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n343), .CK(i_CLK), .Q(a_m[6]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n346), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd state_reg_1_ ( .D(n352), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n285), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_reg_22_ ( .D(n238), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd z_reg_30_ ( .D(n230), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n232), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n234), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n236), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n237), .CK(i_CLK), .Q(z[23]) );
  fad1_hd intadd_23_U2 ( .A(intadd_23_A_18_), .B(intadd_23_B_18_), .CI(
        intadd_23_n2), .CO(intadd_23_n1), .S(intadd_21_A_21_) );
  fad1_hd intadd_23_U3 ( .A(intadd_23_A_17_), .B(intadd_23_B_17_), .CI(
        intadd_23_n3), .CO(intadd_23_n2), .S(intadd_21_A_20_) );
  fad1_hd intadd_23_U18 ( .A(intadd_23_A_2_), .B(intadd_23_B_2_), .CI(
        intadd_23_n18), .CO(intadd_23_n17), .S(intadd_21_A_5_) );
  fad1_hd intadd_23_U17 ( .A(intadd_23_A_3_), .B(intadd_23_B_3_), .CI(
        intadd_23_n17), .CO(intadd_23_n16), .S(intadd_21_A_6_) );
  fad1_hd intadd_21_U3 ( .A(intadd_21_A_23_), .B(intadd_25_n1), .CI(
        intadd_21_n3), .CO(intadd_21_n2), .S(intadd_21_SUM_23_) );
  fd1qd2_hd a_m_reg_20_ ( .D(n329), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n332), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n338), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n341), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n344), .CK(i_CLK), .Q(a_m[5]) );
  fad1_hd intadd_32_U2 ( .A(n1195), .B(intadd_32_B_5_), .CI(intadd_32_n2), 
        .CO(intadd_32_n1), .S(intadd_32_SUM_5_) );
  fad1_hd intadd_37_U2 ( .A(intadd_32_SUM_3_), .B(intadd_37_B_2_), .CI(
        intadd_37_n2), .CO(intadd_37_n1), .S(intadd_37_SUM_2_) );
  fad1_hd intadd_38_U2 ( .A(intadd_31_SUM_7_), .B(intadd_38_B_2_), .CI(
        intadd_38_n2), .CO(intadd_38_n1), .S(intadd_38_SUM_2_) );
  fad1_hd intadd_22_U13 ( .A(n1193), .B(intadd_22_B_8_), .CI(intadd_22_n13), 
        .CO(intadd_22_n12), .S(intadd_22_SUM_8_) );
  fad1_hd DP_OP_125J3_130_6300_U9 ( .A(DP_OP_125J3_130_6300_n26), .B(n1112), 
        .CI(DP_OP_125J3_130_6300_n9), .CO(DP_OP_125J3_130_6300_n8), .S(N468)
         );
  fad1_hd DP_OP_125J3_130_6300_U8 ( .A(DP_OP_125J3_130_6300_n27), .B(n1112), 
        .CI(DP_OP_125J3_130_6300_n8), .CO(DP_OP_125J3_130_6300_n7), .S(N469)
         );
  fad1_hd DP_OP_125J3_130_6300_U7 ( .A(DP_OP_125J3_130_6300_n28), .B(n1112), 
        .CI(DP_OP_125J3_130_6300_n7), .CO(DP_OP_125J3_130_6300_n6), .S(N470)
         );
  fad1_hd DP_OP_125J3_130_6300_U6 ( .A(DP_OP_125J3_130_6300_n29), .B(n1112), 
        .CI(DP_OP_125J3_130_6300_n6), .CO(DP_OP_125J3_130_6300_n5), .S(N471)
         );
  fad1_hd DP_OP_125J3_130_6300_U5 ( .A(DP_OP_125J3_130_6300_n30), .B(n1112), 
        .CI(DP_OP_125J3_130_6300_n5), .CO(DP_OP_125J3_130_6300_n4), .S(N472)
         );
  fad1_hd DP_OP_125J3_130_6300_U4 ( .A(DP_OP_125J3_130_6300_n31), .B(n1112), 
        .CI(DP_OP_125J3_130_6300_n4), .CO(DP_OP_125J3_130_6300_n3), .S(N473)
         );
  fad1_hd DP_OP_125J3_130_6300_U3 ( .A(DP_OP_125J3_130_6300_n32), .B(n1112), 
        .CI(DP_OP_125J3_130_6300_n3), .CO(DP_OP_125J3_130_6300_n2), .S(N474)
         );
  fad1_hd intadd_34_U2 ( .A(n1190), .B(intadd_34_B_2_), .CI(intadd_34_n2), 
        .CO(intadd_34_n1), .S(intadd_34_SUM_2_) );
  fad1_hd intadd_33_U2 ( .A(n1194), .B(intadd_33_B_4_), .CI(intadd_33_n2), 
        .CO(intadd_33_n1), .S(intadd_33_SUM_4_) );
  fad1_hd intadd_36_U4 ( .A(n1221), .B(intadd_36_B_0_), .CI(intadd_36_CI), 
        .CO(intadd_36_n3), .S(intadd_36_SUM_0_) );
  fad1_hd intadd_24_U11 ( .A(n1040), .B(n1039), .CI(intadd_24_n11), .CO(
        intadd_24_n10), .S(intadd_24_SUM_8_) );
  fad1_hd intadd_24_U12 ( .A(n1039), .B(n1037), .CI(intadd_24_n12), .CO(
        intadd_24_n11), .S(intadd_24_SUM_7_) );
  fad1_hd intadd_24_U14 ( .A(n1036), .B(n1034), .CI(intadd_24_n14), .CO(
        intadd_24_n13), .S(intadd_24_SUM_5_) );
  fad1_hd intadd_24_U13 ( .A(n1037), .B(n1036), .CI(intadd_24_n13), .CO(
        intadd_24_n12), .S(intadd_24_SUM_6_) );
  fad1_hd intadd_24_U15 ( .A(n1034), .B(n1032), .CI(intadd_24_n15), .CO(
        intadd_24_n14), .S(intadd_24_SUM_4_) );
  fad1_hd intadd_24_U16 ( .A(n1032), .B(n1031), .CI(intadd_24_n16), .CO(
        intadd_24_n15), .S(intadd_24_SUM_3_) );
  fad1_hd intadd_24_U17 ( .A(n1031), .B(n1030), .CI(intadd_24_n17), .CO(
        intadd_24_n16), .S(intadd_24_SUM_2_) );
  fad1_hd intadd_24_U18 ( .A(n1030), .B(n1011), .CI(intadd_24_n18), .CO(
        intadd_24_n17), .S(intadd_24_SUM_1_) );
  fad1_hd intadd_24_U19 ( .A(n1011), .B(n1027), .CI(intadd_24_CI), .CO(
        intadd_24_n18), .S(intadd_24_SUM_0_) );
  fad1_hd intadd_21_U2 ( .A(intadd_21_A_24_), .B(n1133), .CI(intadd_21_n2), 
        .CO(intadd_21_n1), .S(intadd_21_SUM_24_) );
  fad1_hd intadd_30_U7 ( .A(n1128), .B(n1129), .CI(intadd_30_n7), .CO(
        intadd_30_n6), .S(N206) );
  fad1_hd intadd_30_U6 ( .A(n2024), .B(n1127), .CI(intadd_30_n6), .CO(
        intadd_30_n5), .S(N207) );
  fad1_hd intadd_30_U5 ( .A(n1126), .B(n2023), .CI(intadd_30_n5), .CO(
        intadd_30_n4), .S(N208) );
  fad1_hd intadd_30_U4 ( .A(n1185), .B(n1125), .CI(intadd_30_n4), .CO(
        intadd_30_n3), .S(N209) );
  fad1_hd intadd_22_U5 ( .A(n2029), .B(intadd_34_n1), .CI(intadd_22_n5), .CO(
        intadd_22_n4), .S(N219) );
  fad1_hd intadd_22_U4 ( .A(n1189), .B(n2028), .CI(intadd_22_n4), .CO(
        intadd_22_n3), .S(N220) );
  fad1_hd intadd_22_U3 ( .A(n2037), .B(n1188), .CI(intadd_22_n3), .CO(
        intadd_22_n2), .S(N221) );
  fad1_hd intadd_22_U2 ( .A(n2036), .B(intadd_22_B_19_), .CI(intadd_22_n2), 
        .CO(intadd_22_n1), .S(N222) );
  fad1_hd intadd_22_U6 ( .A(intadd_34_SUM_2_), .B(n1186), .CI(intadd_22_n6), 
        .CO(intadd_22_n5), .S(N218) );
  fad1_hd intadd_30_U8 ( .A(n1131), .B(n1130), .CI(intadd_30_n8), .CO(
        intadd_30_n7), .S(N205) );
  fad1_hd intadd_30_U3 ( .A(n2035), .B(n1184), .CI(intadd_30_n3), .CO(
        intadd_30_n2), .S(N210) );
  fad1_hd intadd_30_U2 ( .A(intadd_22_SUM_8_), .B(n2034), .CI(intadd_30_n2), 
        .CO(intadd_30_n1), .S(N211) );
  fad1_hd intadd_22_U12 ( .A(n1183), .B(intadd_30_n1), .CI(intadd_22_n12), 
        .CO(intadd_22_n11), .S(N212) );
  fad1_hd intadd_22_U11 ( .A(n2033), .B(n1182), .CI(intadd_22_n11), .CO(
        intadd_22_n10), .S(N213) );
  fad1_hd intadd_22_U10 ( .A(intadd_33_SUM_4_), .B(n2032), .CI(intadd_22_n10), 
        .CO(intadd_22_n9), .S(N214) );
  fad1_hd intadd_22_U9 ( .A(n1181), .B(intadd_33_n1), .CI(intadd_22_n9), .CO(
        intadd_22_n8), .S(N215) );
  fad1_hd intadd_22_U8 ( .A(n2031), .B(n1180), .CI(intadd_22_n8), .CO(
        intadd_22_n7), .S(N216) );
  fad1_hd intadd_22_U7 ( .A(n1187), .B(n2030), .CI(intadd_22_n7), .CO(
        intadd_22_n6), .S(N217) );
  fd1qd1_hd sticky_reg ( .D(n283), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n350), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd a_m_reg_23_ ( .D(n355), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd z_reg_31_ ( .D(n229), .CK(i_CLK), .Q(z[31]) );
  fd1qd2_hd b_m_reg_23_ ( .D(n310), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n335), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n347), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd2_hd b_m_reg_0_ ( .D(n308), .CK(i_CLK), .Q(n1022) );
  fad1_hd intadd_24_U5 ( .A(n1050), .B(n1048), .CI(intadd_24_n5), .CO(
        intadd_24_n4), .S(intadd_24_SUM_14_) );
  fad1_hd intadd_24_U7 ( .A(n1046), .B(n1044), .CI(intadd_24_n7), .CO(
        intadd_24_n6), .S(intadd_24_SUM_12_) );
  fad1_hd intadd_24_U6 ( .A(n1048), .B(n1046), .CI(intadd_24_n6), .CO(
        intadd_24_n5), .S(intadd_24_SUM_13_) );
  fad1_hd intadd_24_U2 ( .A(n1055), .B(n1053), .CI(intadd_24_n2), .CO(
        intadd_24_n1), .S(intadd_24_SUM_17_) );
  fad1_hd intadd_24_U4 ( .A(n1051), .B(n1050), .CI(intadd_24_n4), .CO(
        intadd_24_n3), .S(intadd_24_SUM_15_) );
  fad1_hd intadd_24_U3 ( .A(n1053), .B(n1051), .CI(intadd_24_n3), .CO(
        intadd_24_n2), .S(intadd_24_SUM_16_) );
  fad1_hd intadd_24_U10 ( .A(n1041), .B(n1040), .CI(intadd_24_n10), .CO(
        intadd_24_n9), .S(intadd_24_SUM_9_) );
  fad1_hd intadd_24_U9 ( .A(n1043), .B(n1041), .CI(intadd_24_n9), .CO(
        intadd_24_n8), .S(intadd_24_SUM_10_) );
  fad1_hd intadd_24_U8 ( .A(n1044), .B(n1043), .CI(intadd_24_n8), .CO(
        intadd_24_n7), .S(intadd_24_SUM_11_) );
  clknd2d1_hd U367 ( .A(n1176), .B(n1857), .Y(n1140) );
  ivd1_hd U368 ( .A(n1022), .Y(n1014) );
  clknd2d1_hd U369 ( .A(n1060), .B(n1022), .Y(n1910) );
  clknd2d1_hd U370 ( .A(n1354), .B(a_m[20]), .Y(n1343) );
  clknd2d1_hd U371 ( .A(n1022), .B(n1356), .Y(n1404) );
  clknd2d1_hd U372 ( .A(a_m[23]), .B(n1012), .Y(n1912) );
  clknd2d1_hd U373 ( .A(a_m[23]), .B(n1031), .Y(intadd_31_B_2_) );
  clknd2d1_hd U374 ( .A(a_m[23]), .B(n1030), .Y(intadd_31_CI) );
  clknd2d1_hd U375 ( .A(n1374), .B(a_m[17]), .Y(n1375) );
  clknd2d1_hd U376 ( .A(n1022), .B(n1338), .Y(n1378) );
  clknd2d1_hd U377 ( .A(n1034), .B(intadd_31_A_2_), .Y(n1415) );
  clknd2d1_hd U378 ( .A(n1022), .B(n1332), .Y(n1381) );
  clknd2d1_hd U379 ( .A(n1330), .B(a_m[14]), .Y(n1329) );
  clknd2d1_hd U380 ( .A(n1060), .B(n1040), .Y(intadd_32_B_1_) );
  clknd2d1_hd U381 ( .A(a_m[23]), .B(n1036), .Y(n2039) );
  clknd2d1_hd U382 ( .A(a_m[23]), .B(n1039), .Y(n1443) );
  clknd2d1_hd U383 ( .A(a_m[23]), .B(n1523), .Y(n1414) );
  clknd2d1_hd U384 ( .A(n1035), .B(n1033), .Y(n1523) );
  clknd2d1_hd U385 ( .A(n1022), .B(n1284), .Y(n1335) );
  clknd2d1_hd U386 ( .A(n1294), .B(a_m[11]), .Y(n1295) );
  clknd2d1_hd U387 ( .A(n1060), .B(n1044), .Y(intadd_34_A_0_) );
  clknd2d1_hd U388 ( .A(n1043), .B(intadd_32_A_1_), .Y(n1437) );
  clknd2d1_hd U389 ( .A(n1022), .B(n1280), .Y(n1305) );
  clknd2d1_hd U390 ( .A(n1257), .B(a_m[8]), .Y(n1258) );
  clknd2d1_hd U391 ( .A(n1026), .B(n1025), .Y(n1524) );
  clknd2d1_hd U392 ( .A(n1086), .B(n1088), .Y(n1408) );
  clknd2d1_hd U393 ( .A(n1060), .B(n1050), .Y(intadd_36_B_1_) );
  clknd2d1_hd U394 ( .A(n1049), .B(n1045), .Y(n1531) );
  clknd2d1_hd U395 ( .A(n1437), .B(n1436), .Y(n1438) );
  clknd2d1_hd U396 ( .A(b_m[23]), .B(n1058), .Y(n1119) );
  clknd2d1_hd U397 ( .A(n1055), .B(intadd_24_n1), .Y(n1117) );
  clknd2d1_hd U398 ( .A(n1507), .B(n1506), .Y(n1521) );
  clknd2d1_hd U399 ( .A(n1743), .B(n1538), .Y(n1535) );
  clknd2d1_hd U400 ( .A(n1836), .B(n1536), .Y(n1537) );
  clknd2d1_hd U401 ( .A(n1760), .B(n1842), .Y(n1508) );
  clknd2d1_hd U402 ( .A(n1546), .B(n1495), .Y(n1610) );
  clknd2d1_hd U403 ( .A(n1022), .B(n1169), .Y(n1268) );
  clknd2d1_hd U404 ( .A(n1159), .B(a_m[5]), .Y(n1090) );
  clknd2d1_hd U405 ( .A(n1022), .B(n1086), .Y(n1211) );
  clknd2d1_hd U406 ( .A(n1493), .B(n1492), .Y(n1555) );
  clknd2d1_hd U407 ( .A(z_e[7]), .B(z_e[8]), .Y(n1554) );
  clknd2d1_hd U408 ( .A(n1546), .B(n1545), .Y(n1586) );
  clknd2d1_hd U409 ( .A(n1057), .B(n1056), .Y(n1111) );
  clknd2d1_hd U410 ( .A(n1356), .B(n1238), .Y(n1240) );
  clknd2d1_hd U411 ( .A(b_m[23]), .B(n1177), .Y(n1136) );
  clknd2d1_hd U412 ( .A(n1052), .B(n1054), .Y(n1855) );
  clknd2d1_hd U413 ( .A(n1279), .B(n1278), .Y(n1477) );
  xo2d1_hd U414 ( .A(intadd_24_n1), .B(n1217), .Y(n1937) );
  xo2d1_hd U415 ( .A(n1122), .B(n1121), .Y(n1460) );
  clknd2d1_hd U416 ( .A(n1119), .B(n1118), .Y(n1121) );
  clknd2d1_hd U417 ( .A(n1117), .B(n1116), .Y(n1122) );
  clknd2d1_hd U418 ( .A(n1057), .B(n1059), .Y(n1118) );
  ivd1_hd U419 ( .A(b_m[22]), .Y(n1058) );
  clknd2d1_hd U420 ( .A(a_m[0]), .B(n1062), .Y(n1150) );
  ao21d1_hd U421 ( .A(n1058), .B(n1117), .C(n1059), .Y(n1929) );
  clknd2d1_hd U422 ( .A(n1545), .B(n1803), .Y(n1543) );
  clknd2d1_hd U423 ( .A(n1538), .B(n1537), .Y(n1539) );
  clknd2d1_hd U424 ( .A(n1536), .B(n1535), .Y(n1541) );
  ivd2_hd U425 ( .A(n1025), .Y(n1024) );
  ivd2_hd U426 ( .A(n1026), .Y(n1012) );
  ivd1_hd U427 ( .A(b_m[1]), .Y(n1025) );
  ivd1_hd U428 ( .A(b_m[2]), .Y(n1026) );
  ivd2_hd U429 ( .A(n1029), .Y(n1011) );
  ivd2_hd U430 ( .A(n1033), .Y(n1032) );
  nid2_hd U431 ( .A(b_m[9]), .Y(n1036) );
  ivd2_hd U432 ( .A(n1038), .Y(n1037) );
  ivd2_hd U433 ( .A(n1042), .Y(n1041) );
  ivd2_hd U434 ( .A(n1045), .Y(n1044) );
  ivd2_hd U435 ( .A(n1047), .Y(n1046) );
  ivd2_hd U436 ( .A(n1052), .Y(n1051) );
  ivd2_hd U437 ( .A(n1056), .Y(n1055) );
  ivd1_hd U438 ( .A(b_m[21]), .Y(n1056) );
  ivd2_hd U439 ( .A(n1058), .Y(n1057) );
  ivd1_hd U440 ( .A(b_m[7]), .Y(n1033) );
  ivd2_hd U441 ( .A(n1035), .Y(n1034) );
  nid2_hd U442 ( .A(b_m[11]), .Y(n1039) );
  nid2_hd U443 ( .A(b_m[12]), .Y(n1040) );
  nid2_hd U444 ( .A(b_m[14]), .Y(n1043) );
  ivd2_hd U445 ( .A(n1049), .Y(n1048) );
  nid2_hd U446 ( .A(b_m[18]), .Y(n1050) );
  ivd2_hd U447 ( .A(n1054), .Y(n1053) );
  ivd2_hd U448 ( .A(a_m[8]), .Y(n1787) );
  ivd2_hd U449 ( .A(a_m[11]), .Y(n1939) );
  ivd2_hd U450 ( .A(a_m[14]), .Y(n1870) );
  clknd2d1_hd U451 ( .A(n1007), .B(n1832), .Y(n1786) );
  clknd2d1_hd U452 ( .A(N34), .B(n1845), .Y(n1847) );
  clknd2d1_hd U453 ( .A(n1709), .B(n1664), .Y(n1672) );
  clknd2d1_hd U454 ( .A(n1709), .B(n1673), .Y(n1679) );
  clknd2d1_hd U455 ( .A(n1709), .B(n1646), .Y(n1654) );
  clknd2d1_hd U456 ( .A(n1709), .B(n1637), .Y(n1642) );
  clknd2d1_hd U457 ( .A(n1709), .B(n1655), .Y(n1660) );
  clknd2d1_hd U458 ( .A(n1821), .B(n1809), .Y(n1813) );
  clknd2d1_hd U459 ( .A(n1495), .B(n1821), .Y(n1498) );
  clknd2d1_hd U460 ( .A(n1809), .B(n1803), .Y(n1808) );
  clknd2d1_hd U461 ( .A(n1821), .B(n1810), .Y(n1762) );
  clknd2d1_hd U462 ( .A(n1709), .B(n1609), .Y(n1618) );
  clknd2d1_hd U463 ( .A(n1709), .B(n1628), .Y(n1636) );
  clknd2d1_hd U464 ( .A(n1709), .B(n1619), .Y(n1624) );
  clknd2d1_hd U465 ( .A(n1821), .B(n1545), .Y(n1699) );
  clknd2d1_hd U466 ( .A(n1546), .B(n1810), .Y(n1818) );
  clknd2d1_hd U467 ( .A(n1709), .B(n1600), .Y(n1605) );
  clknd2d1_hd U468 ( .A(n1597), .B(n1595), .Y(n1712) );
  clknd2d1_hd U469 ( .A(n1709), .B(n1596), .Y(n1595) );
  clknd2d1_hd U470 ( .A(n1069), .B(n1068), .Y(n1070) );
  clknd2d1_hd U471 ( .A(n1211), .B(n1070), .Y(n1075) );
  clknd2d1_hd U472 ( .A(n1074), .B(n1075), .Y(intadd_21_A_0_) );
  clknd2d1_hd U473 ( .A(n1580), .B(n1576), .Y(n1575) );
  clknd2d1_hd U474 ( .A(n1572), .B(n1569), .Y(n1568) );
  clknd2d1_hd U475 ( .A(n1565), .B(n1562), .Y(n1561) );
  clknd2d1_hd U476 ( .A(n1056), .B(n1059), .Y(n1525) );
  clknd2d1_hd U477 ( .A(n1219), .B(n1111), .Y(n1076) );
  ivd2_hd U478 ( .A(n1060), .Y(n1061) );
  clknd2d1_hd U479 ( .A(n1053), .B(intadd_36_A_1_), .Y(n1856) );
  clknd2d1_hd U480 ( .A(n1140), .B(n1136), .Y(n1144) );
  clknd2d1_hd U481 ( .A(state[1]), .B(state[0]), .Y(n1820) );
  clknd2d1_hd U482 ( .A(n1833), .B(a_e[7]), .Y(n1744) );
  clknd2d1_hd U483 ( .A(n1013), .B(n1548), .Y(n1549) );
  clknd2d1_hd U484 ( .A(n1810), .B(n1803), .Y(n1805) );
  clknd2d1_hd U485 ( .A(n1016), .B(z[23]), .Y(n1583) );
  clknd2d1_hd U486 ( .A(n1016), .B(z[24]), .Y(n1581) );
  clknd2d1_hd U487 ( .A(n1016), .B(z[26]), .Y(n1573) );
  clknd2d1_hd U488 ( .A(n1016), .B(z[28]), .Y(n1566) );
  clknd2d1_hd U489 ( .A(z_e[7]), .B(n1561), .Y(n1559) );
  clknd2d1_hd U490 ( .A(n1016), .B(z[22]), .Y(n1588) );
  clknd2d1_hd U491 ( .A(state[2]), .B(state[3]), .Y(n1827) );
  clknd2d1_hd U492 ( .A(n1750), .B(n138), .Y(n317) );
  clknd2d1_hd U493 ( .A(n1766), .B(n148), .Y(n326) );
  clknd2d1_hd U494 ( .A(n1708), .B(n1687), .Y(n1690) );
  clknd2d1_hd U495 ( .A(n1688), .B(n1687), .Y(n1685) );
  clknd2d1_hd U496 ( .A(z_m[0]), .B(n1709), .Y(n1683) );
  clknd2d1_hd U497 ( .A(n1709), .B(n1814), .Y(n1716) );
  clknd2d1_hd U498 ( .A(z_m[23]), .B(n1591), .Y(n1500) );
  clknd2d1_hd U499 ( .A(n1840), .B(n1839), .Y(n1837) );
  clknd2d1_hd U500 ( .A(b_e[9]), .B(n1850), .Y(n1839) );
  clknd2d1_hd U501 ( .A(n1756), .B(n1755), .Y(n1753) );
  clknd2d1_hd U502 ( .A(n1748), .B(n138), .Y(n311) );
  clknd2d1_hd U503 ( .A(b_e[8]), .B(n1763), .Y(n1764) );
  clknd2d1_hd U504 ( .A(n1499), .B(n1699), .Y(n105) );
  clknd2d1_hd U505 ( .A(a_m[2]), .B(N176), .Y(n1064) );
  clknd2d1_hd U506 ( .A(n1584), .B(n1579), .Y(n235) );
  clknd2d1_hd U507 ( .A(n1552), .B(n1843), .Y(n148) );
  clknd2d1_hd U508 ( .A(n1552), .B(n1759), .Y(n138) );
  ivd1_hd U509 ( .A(b_m[23]), .Y(n1059) );
  ivd1_hd U510 ( .A(intadd_21_n1), .Y(n1131) );
  scg16d2_hd U512 ( .A(n1117), .B(n1119), .C(n1091), .Y(n1857) );
  xo2d1_hd U513 ( .A(n1028), .B(n1072), .Y(n1396) );
  ivd1_hd U514 ( .A(b_m[8]), .Y(n1035) );
  ivd1_hd U515 ( .A(b_m[17]), .Y(n1049) );
  nr2d2_hd U516 ( .A(n1284), .B(n1232), .Y(n1868) );
  nr2d2_hd U517 ( .A(n1279), .B(n1281), .Y(n1936) );
  nr2d2_hd U518 ( .A(n1332), .B(n1229), .Y(n1880) );
  scg12d2_hd U519 ( .A(n1228), .B(n1229), .C(n1332), .Y(n1889) );
  ivd1_hd U520 ( .A(b_m[15]), .Y(n1045) );
  ivd1_hd U521 ( .A(b_m[19]), .Y(n1052) );
  xo2d1_hd U522 ( .A(n1019), .B(n1293), .Y(intadd_25_B_16_) );
  xo2d1_hd U523 ( .A(n1019), .B(n1246), .Y(intadd_23_A_18_) );
  xo2d1_hd U524 ( .A(n1337), .B(n1336), .Y(intadd_26_CI) );
  xo2d1_hd U525 ( .A(n1270), .B(n1269), .Y(intadd_23_CI) );
  xo2d1_hd U526 ( .A(n1216), .B(n1214), .Y(intadd_21_CI) );
  xo2d1_hd U527 ( .A(n1361), .B(n1360), .Y(intadd_27_CI) );
  nid2_hd U528 ( .A(n1933), .Y(n1009) );
  xo2d1_hd U529 ( .A(n1787), .B(n1422), .Y(intadd_31_B_3_) );
  ivd2_hd U530 ( .A(n1150), .Y(n1176) );
  ivd2_hd U531 ( .A(n1408), .Y(n1290) );
  ad2d2_hd U532 ( .A(n1226), .B(n1338), .Y(n1919) );
  nr2d2_hd U533 ( .A(n1086), .B(n1085), .Y(n1292) );
  nr2d2_hd U534 ( .A(n1169), .B(n1094), .Y(n1486) );
  ivd1_hd U535 ( .A(b_m[20]), .Y(n1054) );
  ivd1_hd U536 ( .A(b_m[3]), .Y(n1028) );
  ivd1_hd U537 ( .A(b_m[16]), .Y(n1047) );
  nid2_hd U538 ( .A(a_m[23]), .Y(n1060) );
  ivd1_hd U539 ( .A(b_m[13]), .Y(n1042) );
  ivd1_hd U540 ( .A(b_m[10]), .Y(n1038) );
  xo2d1_hd U541 ( .A(n1939), .B(n1478), .Y(intadd_39_B_2_) );
  xo2d1_hd U542 ( .A(n1787), .B(n1489), .Y(intadd_41_B_2_) );
  xo2d1_hd U543 ( .A(n1939), .B(n1352), .Y(intadd_27_B_13_) );
  xo2d1_hd U544 ( .A(a_m[14]), .B(n1236), .Y(intadd_22_B_8_) );
  xo2d1_hd U545 ( .A(a_m[5]), .B(n1410), .Y(intadd_30_B_0_) );
  xo2d1_hd U546 ( .A(n1021), .B(n1123), .Y(intadd_21_B_19_) );
  xo2d1_hd U547 ( .A(n1061), .B(n1461), .Y(intadd_36_B_2_) );
  xo2d1_hd U548 ( .A(a_m[17]), .B(n1446), .Y(intadd_33_B_4_) );
  xo2d1_hd U549 ( .A(n1870), .B(n1472), .Y(intadd_38_B_2_) );
  xo2d1_hd U550 ( .A(a_m[20]), .B(n1452), .Y(intadd_34_B_2_) );
  xo2d1_hd U551 ( .A(n1061), .B(n1860), .Y(n1862) );
  xo2d1_hd U552 ( .A(n1787), .B(n1327), .Y(intadd_26_B_16_) );
  xo2d1_hd U553 ( .A(n1019), .B(n1093), .Y(n1099) );
  xo2d1_hd U554 ( .A(n1020), .B(n1467), .Y(intadd_37_B_2_) );
  xo2d1_hd U555 ( .A(n1892), .B(n1440), .Y(intadd_32_B_5_) );
  xo2d1_hd U556 ( .A(a_m[11]), .B(n1866), .Y(n1873) );
  xo2d1_hd U557 ( .A(a_m[8]), .B(n1932), .Y(n1942) );
  xo2d1_hd U558 ( .A(a_m[20]), .B(n1897), .Y(n1901) );
  xo2d1_hd U559 ( .A(a_m[14]), .B(n1878), .Y(n1885) );
  xo2d1_hd U560 ( .A(a_m[17]), .B(n1890), .Y(n1895) );
  xo2d1_hd U561 ( .A(n1870), .B(n1869), .Y(n1872) );
  xo2d1_hd U562 ( .A(n1061), .B(n1898), .Y(n1900) );
  xo2d1_hd U563 ( .A(n1939), .B(n1938), .Y(n1941) );
  xo2d1_hd U564 ( .A(n1021), .B(n1115), .Y(intadd_21_B_18_) );
  xo2d1_hd U565 ( .A(n1892), .B(n1891), .Y(n1894) );
  xo2d1_hd U566 ( .A(n1020), .B(n1881), .Y(n1884) );
  xo2d1_hd U567 ( .A(a_m[8]), .B(n1412), .Y(intadd_30_CI) );
  xo2d1_hd U568 ( .A(n1021), .B(n1110), .Y(intadd_21_B_17_) );
  xo2d1_hd U569 ( .A(a_m[14]), .B(n1235), .Y(intadd_22_B_6_) );
  xo2d1_hd U570 ( .A(n1019), .B(n1256), .Y(intadd_23_B_17_) );
  xo2d1_hd U571 ( .A(n1939), .B(n1351), .Y(intadd_27_B_11_) );
  xo2d1_hd U572 ( .A(n1787), .B(n1097), .Y(n1098) );
  xo2d1_hd U573 ( .A(n1020), .B(n1425), .Y(intadd_31_B_7_) );
  xo2d1_hd U574 ( .A(n1892), .B(n1439), .Y(intadd_32_B_3_) );
  xo2d1_hd U575 ( .A(n1061), .B(n1462), .Y(intadd_36_CI) );
  xo2d1_hd U576 ( .A(n1892), .B(n1465), .Y(intadd_37_B_1_) );
  xo2d1_hd U577 ( .A(n1020), .B(n1469), .Y(intadd_38_B_1_) );
  xo2d1_hd U578 ( .A(n1870), .B(n1475), .Y(intadd_39_B_1_) );
  xo2d1_hd U579 ( .A(n1787), .B(n1311), .Y(intadd_26_A_13_) );
  xo2d1_hd U580 ( .A(n1019), .B(n1255), .Y(intadd_23_B_16_) );
  xo2d1_hd U581 ( .A(n1939), .B(n1485), .Y(intadd_41_A_1_) );
  xo2d1_hd U582 ( .A(n1021), .B(n1109), .Y(intadd_21_B_16_) );
  xo2d1_hd U583 ( .A(n1060), .B(n1448), .Y(intadd_34_A_1_) );
  xo2d1_hd U584 ( .A(n1939), .B(n1490), .Y(intadd_41_CI) );
  xo2d1_hd U585 ( .A(n1787), .B(n1276), .Y(intadd_25_A_15_) );
  xo2d1_hd U586 ( .A(n1060), .B(n1453), .Y(intadd_34_CI) );
  xo2d1_hd U587 ( .A(n1892), .B(n1464), .Y(intadd_37_B_0_) );
  xo2d1_hd U588 ( .A(n1021), .B(n1108), .Y(intadd_21_B_15_) );
  xo2d1_hd U589 ( .A(n1019), .B(n1254), .Y(intadd_23_B_15_) );
  xo2d1_hd U590 ( .A(n1870), .B(n1479), .Y(intadd_39_CI) );
  xo2d1_hd U591 ( .A(n1020), .B(n1473), .Y(intadd_38_CI) );
  xo2d1_hd U592 ( .A(n1787), .B(n1288), .Y(intadd_25_B_14_) );
  xo2d1_hd U593 ( .A(n1021), .B(n1107), .Y(intadd_21_B_14_) );
  xo2d1_hd U594 ( .A(a_m[20]), .B(n1445), .Y(intadd_33_B_2_) );
  xo2d1_hd U595 ( .A(n1019), .B(n1253), .Y(intadd_23_B_14_) );
  xo2d1_hd U596 ( .A(n1939), .B(n1323), .Y(n1326) );
  xo2d1_hd U597 ( .A(n1870), .B(n1403), .Y(intadd_29_B_8_) );
  xo2d1_hd U598 ( .A(n1060), .B(n1429), .Y(n1431) );
  xo2d1_hd U599 ( .A(n1020), .B(n1482), .Y(intadd_40_B_2_) );
  xo2d1_hd U600 ( .A(n1021), .B(n1105), .Y(intadd_21_B_13_) );
  xo2d1_hd U601 ( .A(n1892), .B(n1424), .Y(intadd_31_B_6_) );
  xo2d1_hd U602 ( .A(n1939), .B(n1364), .Y(intadd_28_A_10_) );
  xo2d1_hd U603 ( .A(n1061), .B(n1426), .Y(intadd_32_A_2_) );
  xo2d1_hd U604 ( .A(n1019), .B(n1245), .Y(intadd_23_A_13_) );
  xo2d1_hd U605 ( .A(a_m[17]), .B(n1231), .Y(intadd_22_B_5_) );
  xo2d1_hd U606 ( .A(n1787), .B(n1275), .Y(intadd_25_A_13_) );
  xo2d1_hd U607 ( .A(n1870), .B(n1341), .Y(intadd_27_A_10_) );
  xo2d1_hd U608 ( .A(n1787), .B(n1287), .Y(intadd_25_B_12_) );
  xo2d1_hd U609 ( .A(n1061), .B(n1463), .Y(intadd_37_A_0_) );
  xo2d1_hd U610 ( .A(n1019), .B(n1252), .Y(intadd_23_B_12_) );
  xo2d1_hd U611 ( .A(n1021), .B(n1104), .Y(intadd_21_B_12_) );
  xo2d1_hd U612 ( .A(n1870), .B(n1484), .Y(intadd_41_A_0_) );
  xo2d1_hd U613 ( .A(n1020), .B(n1474), .Y(intadd_39_B_0_) );
  xo2d1_hd U614 ( .A(n1892), .B(n1468), .Y(intadd_38_B_0_) );
  xo2d1_hd U615 ( .A(n1939), .B(n1322), .Y(intadd_26_B_12_) );
  xo2d1_hd U616 ( .A(n1939), .B(n1310), .Y(intadd_26_A_11_) );
  xo2d1_hd U617 ( .A(n1019), .B(n1251), .Y(intadd_23_B_11_) );
  xo2d1_hd U618 ( .A(n1061), .B(n1441), .Y(intadd_32_CI) );
  xo2d1_hd U619 ( .A(n1870), .B(n1324), .Y(n1325) );
  xo2d1_hd U620 ( .A(n1892), .B(n1423), .Y(intadd_31_B_4_) );
  xo2d1_hd U621 ( .A(n1787), .B(n1286), .Y(intadd_25_B_11_) );
  xo2d1_hd U622 ( .A(n1021), .B(n1103), .Y(intadd_21_B_11_) );
  xo2d1_hd U623 ( .A(a_m[17]), .B(n1230), .Y(intadd_22_B_3_) );
  xo2d1_hd U624 ( .A(n1787), .B(n1274), .Y(intadd_25_A_10_) );
  xo2d1_hd U625 ( .A(n1020), .B(n1402), .Y(intadd_29_B_7_) );
  xo2d1_hd U626 ( .A(n1870), .B(n1348), .Y(intadd_27_A_7_) );
  xo2d1_hd U627 ( .A(n1939), .B(n1321), .Y(intadd_26_B_10_) );
  xo2d1_hd U628 ( .A(n1021), .B(n1102), .Y(intadd_21_B_10_) );
  xo2d1_hd U629 ( .A(n1892), .B(n1481), .Y(intadd_40_B_1_) );
  xo2d1_hd U630 ( .A(n1060), .B(n1442), .Y(intadd_33_A_1_) );
  xo2d1_hd U631 ( .A(n1019), .B(n1244), .Y(intadd_23_A_10_) );
  xo2d1_hd U632 ( .A(n1870), .B(n1380), .Y(intadd_28_B_9_) );
  xo2d1_hd U633 ( .A(n1939), .B(n1319), .Y(intadd_26_A_9_) );
  xo2d1_hd U634 ( .A(n1892), .B(n1483), .Y(intadd_40_CI) );
  xo2d1_hd U635 ( .A(a_m[23]), .B(n1447), .Y(intadd_33_CI) );
  xo2d1_hd U636 ( .A(n1021), .B(n1202), .Y(intadd_21_B_9_) );
  xo2d1_hd U637 ( .A(n1019), .B(n1267), .Y(intadd_23_B_9_) );
  xo2d1_hd U638 ( .A(n1020), .B(n1359), .Y(intadd_27_B_9_) );
  xo2d1_hd U639 ( .A(a_m[20]), .B(n1455), .Y(intadd_35_B_2_) );
  xo2d1_hd U640 ( .A(n1020), .B(n1349), .Y(intadd_27_A_8_) );
  xo2d1_hd U641 ( .A(a_m[23]), .B(n1416), .Y(n1418) );
  xo2d1_hd U642 ( .A(n1021), .B(n1175), .Y(intadd_21_B_8_) );
  xo2d1_hd U643 ( .A(n1939), .B(n1334), .Y(intadd_26_B_8_) );
  xo2d1_hd U644 ( .A(n1019), .B(n1266), .Y(intadd_23_B_8_) );
  xo2d1_hd U645 ( .A(n1870), .B(n1372), .Y(intadd_28_A_8_) );
  xo2d1_hd U646 ( .A(DP_OP_125J3_130_6300_n2), .B(n1083), .Y(n1084) );
  xo2d1_hd U647 ( .A(a_m[20]), .B(n1227), .Y(intadd_22_B_2_) );
  xo2d1_hd U648 ( .A(n1021), .B(n1174), .Y(intadd_21_B_7_) );
  xo2d1_hd U649 ( .A(n1061), .B(n1413), .Y(intadd_31_A_3_) );
  xo2d1_hd U650 ( .A(n1020), .B(n1393), .Y(intadd_29_A_4_) );
  xo2d1_hd U651 ( .A(n1870), .B(n1371), .Y(intadd_28_A_7_) );
  xo2d1_hd U652 ( .A(n1019), .B(n1265), .Y(intadd_23_B_7_) );
  xo2d1_hd U653 ( .A(n1061), .B(n1480), .Y(intadd_40_B_0_) );
  xo2d1_hd U654 ( .A(n1020), .B(n1358), .Y(intadd_27_B_6_) );
  xo2d1_hd U655 ( .A(n1019), .B(n1264), .Y(intadd_23_B_6_) );
  xo2d1_hd U656 ( .A(n1021), .B(n1173), .Y(intadd_21_B_6_) );
  xo2d1_hd U657 ( .A(n1870), .B(n1370), .Y(intadd_28_A_6_) );
  xo2d1_hd U658 ( .A(n1892), .B(n1401), .Y(intadd_29_B_6_) );
  xo2d1_hd U659 ( .A(n1061), .B(n1421), .Y(intadd_31_B_1_) );
  xo2d1_hd U660 ( .A(n1021), .B(n1172), .Y(intadd_21_B_5_) );
  xo2d1_hd U661 ( .A(n1019), .B(n1263), .Y(intadd_23_B_5_) );
  xo2d1_hd U662 ( .A(n1892), .B(n1400), .Y(n1851) );
  xo2d1_hd U663 ( .A(n1020), .B(n1347), .Y(intadd_27_A_5_) );
  xo2d1_hd U664 ( .A(n1870), .B(n1369), .Y(intadd_28_A_5_) );
  xo2d1_hd U665 ( .A(n1021), .B(n1171), .Y(intadd_21_B_4_) );
  xo2d1_hd U666 ( .A(n1019), .B(n1262), .Y(intadd_23_B_4_) );
  xo2d1_hd U667 ( .A(n1020), .B(n1346), .Y(intadd_27_A_4_) );
  xo2d1_hd U668 ( .A(n1870), .B(n1368), .Y(intadd_28_A_4_) );
  xo2d1_hd U669 ( .A(a_m[20]), .B(n1923), .Y(n1925) );
  scg2d1_hd U670 ( .A(z_e[8]), .B(n1844), .C(n1010), .D(
        DP_OP_125J3_130_6300_n42), .Y(DP_OP_125J3_130_6300_n32) );
  xo2d1_hd U671 ( .A(n1892), .B(n1398), .Y(intadd_29_B_3_) );
  xo2d1_hd U672 ( .A(n1163), .B(n1090), .Y(intadd_21_A_1_) );
  xo2d1_hd U673 ( .A(n1296), .B(n1295), .Y(intadd_25_B_1_) );
  xo2d1_hd U674 ( .A(n1019), .B(n1261), .Y(intadd_23_B_3_) );
  xo2d1_hd U675 ( .A(n1259), .B(n1258), .Y(intadd_23_B_1_) );
  xo2d1_hd U676 ( .A(n1021), .B(n1170), .Y(intadd_21_B_3_) );
  xo2d1_hd U677 ( .A(n1870), .B(n1367), .Y(intadd_28_A_3_) );
  xo2d1_hd U678 ( .A(n1020), .B(n1345), .Y(intadd_27_A_3_) );
  xo2d1_hd U679 ( .A(n1020), .B(n1344), .Y(intadd_27_A_2_) );
  xo2d1_hd U680 ( .A(n1892), .B(n1392), .Y(intadd_29_A_2_) );
  xo2d1_hd U681 ( .A(n1355), .B(n1343), .Y(intadd_27_A_1_) );
  xo2d1_hd U682 ( .A(n1870), .B(n1366), .Y(intadd_28_A_2_) );
  xo2d1_hd U683 ( .A(n1376), .B(n1375), .Y(intadd_28_B_1_) );
  xo2d1_hd U684 ( .A(n1019), .B(n1260), .Y(intadd_23_B_2_) );
  scg2d1_hd U685 ( .A(z_e[7]), .B(n1844), .C(n1010), .D(
        DP_OP_125J3_130_6300_n41), .Y(DP_OP_125J3_130_6300_n31) );
  xo2d1_hd U686 ( .A(n1331), .B(n1329), .Y(intadd_26_B_1_) );
  xo2d1_hd U687 ( .A(n1021), .B(n1100), .Y(intadd_21_A_2_) );
  xo2d1_hd U688 ( .A(n1892), .B(n1395), .Y(intadd_29_B_1_) );
  xo2d1_hd U689 ( .A(n1019), .B(n1247), .Y(intadd_23_A_1_) );
  xo2d1_hd U690 ( .A(n1406), .B(n1405), .Y(intadd_29_CI) );
  xo2d1_hd U691 ( .A(n1870), .B(n1365), .Y(intadd_28_A_1_) );
  xo2d1_hd U692 ( .A(n1020), .B(n1353), .Y(intadd_27_B_1_) );
  xo2d1_hd U693 ( .A(n1307), .B(n1306), .Y(intadd_25_CI) );
  xo2d1_hd U694 ( .A(n1061), .B(n1399), .Y(n1913) );
  scg6d1_hd U695 ( .A(n1552), .B(n1547), .C(n1551), .Y(n1013) );
  scg2d1_hd U696 ( .A(z_e[6]), .B(n1844), .C(n1010), .D(
        DP_OP_125J3_130_6300_n40), .Y(DP_OP_125J3_130_6300_n30) );
  xo2d1_hd U697 ( .A(n1019), .B(n1250), .Y(intadd_23_B_0_) );
  xo2d1_hd U698 ( .A(n1060), .B(n1907), .Y(n1918) );
  xo2d1_hd U699 ( .A(n1892), .B(n1394), .Y(intadd_29_B_0_) );
  xo2d1_hd U700 ( .A(n1383), .B(n1382), .Y(intadd_28_CI) );
  xo2d1_hd U701 ( .A(n1061), .B(n1387), .Y(n1391) );
  xo2d1_hd U702 ( .A(n1020), .B(n1350), .Y(intadd_27_B_0_) );
  scg2d1_hd U703 ( .A(n1388), .B(n1290), .C(n1024), .D(n1291), .Y(n1089) );
  scg2d1_hd U704 ( .A(n1388), .B(n1930), .C(n1024), .D(n1411), .Y(n1249) );
  scg2d1_hd U705 ( .A(n1388), .B(n1936), .C(n1022), .D(n1935), .Y(n1282) );
  scg2d1_hd U706 ( .A(n1388), .B(n1903), .C(n1024), .D(n1906), .Y(n1389) );
  xo2d1_hd U707 ( .A(n1870), .B(n1438), .Y(intadd_32_B_2_) );
  scg2d1_hd U708 ( .A(n1388), .B(n1919), .C(n1024), .D(n1922), .Y(n1342) );
  ivd2_hd U709 ( .A(n1240), .Y(n1903) );
  ad2bd2_hd U710 ( .B(n1096), .AN(n1095), .Y(n1930) );
  nr2bd2_hd U711 ( .AN(n1332), .B(n1228), .Y(n1879) );
  ivd6_hd U712 ( .A(n1817), .Y(n2022) );
  ao21d1_hd U713 ( .A(n1022), .B(n1024), .C(n1012), .Y(n1271) );
  nr2d4_hd U714 ( .A(a_m[0]), .B(n1800), .Y(n1177) );
  nr2bd1_hd U715 ( .AN(state[0]), .B(state[1]), .Y(n1495) );
  xo2d1_hd U716 ( .A(a_s), .B(b_s), .Y(N35) );
  oa22ad1_hd U717 ( .A(a_m[21]), .B(a_m[22]), .C(a_m[22]), .D(a_m[21]), .Y(
        n1239) );
  xo3d1_hd U718 ( .A(n1079), .B(intadd_22_n1), .C(n1078), .Y(N223) );
  xn2d1_hd U719 ( .A(n1219), .B(n1218), .Y(intadd_22_B_19_) );
  xo2d1_hd U720 ( .A(n1084), .B(n1813), .Y(N475) );
  xo2d1_hd U721 ( .A(n1787), .B(n1304), .Y(intadd_25_B_9_) );
  xo2d1_hd U722 ( .A(n1787), .B(n1303), .Y(intadd_25_B_8_) );
  xo2d1_hd U723 ( .A(n1939), .B(n1318), .Y(intadd_26_A_7_) );
  xo2d1_hd U724 ( .A(n1787), .B(n1302), .Y(intadd_25_B_7_) );
  scg2d1_hd U725 ( .A(b_e[2]), .B(n1765), .C(n1838), .D(C82_DATA2_2), .Y(n325)
         );
  xo2d1_hd U726 ( .A(n1787), .B(n1301), .Y(intadd_25_B_6_) );
  scg2d1_hd U727 ( .A(b_e[6]), .B(n1765), .C(n1838), .D(C82_DATA2_6), .Y(n321)
         );
  scg2d1_hd U728 ( .A(b_e[5]), .B(n1765), .C(n1838), .D(C82_DATA2_5), .Y(n322)
         );
  scg2d1_hd U729 ( .A(b_e[4]), .B(n1765), .C(n1838), .D(C82_DATA2_4), .Y(n323)
         );
  xo2d1_hd U730 ( .A(n1939), .B(n1317), .Y(intadd_26_A_6_) );
  scg2d1_hd U731 ( .A(b_e[3]), .B(n1765), .C(n1838), .D(C82_DATA2_3), .Y(n324)
         );
  scg2d1_hd U732 ( .A(a_e[6]), .B(n1749), .C(C81_DATA2_6), .D(n1754), .Y(n312)
         );
  xo2d1_hd U733 ( .A(n1939), .B(n1316), .Y(intadd_26_A_5_) );
  xo2d1_hd U734 ( .A(n1787), .B(n1300), .Y(intadd_25_B_5_) );
  scg2d1_hd U735 ( .A(z_m[15]), .B(n1590), .C(n1016), .D(z[15]), .Y(n245) );
  scg2d1_hd U736 ( .A(z_m[18]), .B(n1590), .C(n1016), .D(z[18]), .Y(n242) );
  scg2d1_hd U737 ( .A(z_m[9]), .B(n1590), .C(n1016), .D(z[9]), .Y(n251) );
  scg2d1_hd U738 ( .A(z_m[14]), .B(n1590), .C(n1016), .D(z[14]), .Y(n246) );
  scg2d1_hd U739 ( .A(a_e[5]), .B(n1749), .C(C81_DATA2_5), .D(n1754), .Y(n313)
         );
  scg2d1_hd U740 ( .A(z_m[10]), .B(n1590), .C(n1016), .D(z[10]), .Y(n250) );
  scg2d1_hd U741 ( .A(z_m[17]), .B(n1590), .C(n1016), .D(z[17]), .Y(n243) );
  scg2d1_hd U742 ( .A(z_m[11]), .B(n1590), .C(n1016), .D(z[11]), .Y(n249) );
  scg2d1_hd U743 ( .A(z_m[13]), .B(n1590), .C(n1016), .D(z[13]), .Y(n247) );
  scg2d1_hd U744 ( .A(z_m[12]), .B(n1590), .C(n1016), .D(z[12]), .Y(n248) );
  scg2d1_hd U745 ( .A(z_m[16]), .B(n1590), .C(n1016), .D(z[16]), .Y(n244) );
  scg2d1_hd U746 ( .A(a_e[2]), .B(n1749), .C(C81_DATA2_2), .D(n1754), .Y(n316)
         );
  scg2d1_hd U747 ( .A(z_m[20]), .B(n1590), .C(n1016), .D(z[20]), .Y(n240) );
  scg2d1_hd U748 ( .A(a_e[3]), .B(n1749), .C(C81_DATA2_3), .D(n1754), .Y(n315)
         );
  scg2d1_hd U749 ( .A(z_m[21]), .B(n1590), .C(n1016), .D(z[21]), .Y(n239) );
  scg9d1_hd U750 ( .A(n1075), .B(n1074), .C(intadd_21_A_0_), .Y(N179) );
  scg2d1_hd U751 ( .A(a_e[4]), .B(n1749), .C(C81_DATA2_4), .D(n1754), .Y(n314)
         );
  scg10d1_hd U752 ( .A(n1589), .B(n1549), .C(z[31]), .D(n1013), .Y(n229) );
  scg2d1_hd U753 ( .A(z_m[19]), .B(n1590), .C(n1016), .D(z[19]), .Y(n241) );
  xo2d1_hd U754 ( .A(n1787), .B(n1299), .Y(intadd_25_B_4_) );
  xo2d1_hd U755 ( .A(a_m[23]), .B(n1454), .Y(intadd_35_A_1_) );
  xo2d1_hd U756 ( .A(n1939), .B(n1315), .Y(intadd_26_A_4_) );
  scg2d1_hd U757 ( .A(z_m[5]), .B(n1590), .C(n1016), .D(z[5]), .Y(n255) );
  scg2d1_hd U758 ( .A(z_m[6]), .B(n1590), .C(n1016), .D(z[6]), .Y(n254) );
  scg2d1_hd U759 ( .A(z_m[7]), .B(n1590), .C(n1016), .D(z[7]), .Y(n253) );
  scg2d1_hd U760 ( .A(z_m[8]), .B(n1590), .C(n1016), .D(z[8]), .Y(n252) );
  xo2d1_hd U761 ( .A(a_m[23]), .B(n1456), .Y(intadd_35_CI) );
  xo2d1_hd U762 ( .A(n1939), .B(n1314), .Y(intadd_26_A_3_) );
  xo2d1_hd U763 ( .A(n1787), .B(n1298), .Y(intadd_25_B_3_) );
  xo2d1_hd U764 ( .A(n1787), .B(n1297), .Y(intadd_25_B_2_) );
  scg9d1_hd U765 ( .A(n1069), .B(n1068), .C(n1070), .Y(N178) );
  xo2d1_hd U766 ( .A(n1939), .B(n1313), .Y(intadd_26_A_2_) );
  or2d1_hd U767 ( .A(n1391), .B(n1390), .Y(n1909) );
  xo2d1_hd U768 ( .A(a_m[23]), .B(n1241), .Y(intadd_22_CI) );
  xo2d1_hd U769 ( .A(n1021), .B(n1124), .Y(intadd_21_B_1_) );
  xo2d1_hd U770 ( .A(n1939), .B(n1320), .Y(intadd_26_B_0_) );
  xo2d1_hd U771 ( .A(n1939), .B(n1312), .Y(intadd_26_A_1_) );
  xo2d1_hd U772 ( .A(a_m[11]), .B(n1283), .Y(n1308) );
  xo2d1_hd U773 ( .A(n1870), .B(n1373), .Y(intadd_28_B_0_) );
  xo2d1_hd U774 ( .A(n1787), .B(n1277), .Y(intadd_25_A_1_) );
  xo2d1_hd U775 ( .A(a_m[14]), .B(n1333), .Y(n1362) );
  scg2d1_hd U776 ( .A(n1120), .B(a[0]), .C(n1830), .D(a_m[0]), .Y(n349) );
  xo2d1_hd U777 ( .A(a_m[2]), .B(n1073), .Y(n1074) );
  xo2d1_hd U778 ( .A(a_m[5]), .B(n1167), .Y(n1242) );
  xo2d1_hd U779 ( .A(a_m[20]), .B(n1357), .Y(n1384) );
  xo2d1_hd U780 ( .A(a_m[17]), .B(n1340), .Y(n1377) );
  xo2d1_hd U781 ( .A(n1021), .B(n1101), .Y(intadd_21_B_0_) );
  xo2d1_hd U782 ( .A(a_m[2]), .B(n1067), .Y(n1068) );
  xn2d1_hd U783 ( .A(n1065), .B(n1064), .Y(N177) );
  xo2d1_hd U784 ( .A(a_m[8]), .B(n1248), .Y(n1272) );
  xo2d1_hd U785 ( .A(n1061), .B(n1397), .Y(n1908) );
  scg2d1_hd U786 ( .A(n1388), .B(n1876), .C(n1024), .D(n1867), .Y(n1328) );
  xo2d1_hd U787 ( .A(n1787), .B(n1285), .Y(intadd_25_B_0_) );
  scg2d1_hd U788 ( .A(n1120), .B(b[0]), .C(n1022), .D(n1018), .Y(n308) );
  scg2d1_hd U789 ( .A(n1120), .B(b[28]), .C(b_e[5]), .D(n1850), .Y(n774) );
  scg2d1_hd U790 ( .A(n1120), .B(b[27]), .C(b_e[4]), .D(n1850), .Y(n773) );
  scg2d1_hd U791 ( .A(n1120), .B(b[26]), .C(b_e[3]), .D(n1850), .Y(n772) );
  scg2d1_hd U792 ( .A(n1120), .B(b[25]), .C(b_e[2]), .D(n1850), .Y(n771) );
  scg2d1_hd U793 ( .A(n1120), .B(b[24]), .C(b_e[1]), .D(n1850), .Y(n770) );
  scg2d1_hd U794 ( .A(n1120), .B(b[23]), .C(b_e[0]), .D(n1850), .Y(n769) );
  scg2d1_hd U795 ( .A(n1120), .B(b[29]), .C(b_e[6]), .D(n1850), .Y(n775) );
  scg2d1_hd U796 ( .A(n1120), .B(a[28]), .C(n1833), .D(a_e[5]), .Y(C1_Z_5) );
  scg2d1_hd U797 ( .A(n1120), .B(a[27]), .C(n1833), .D(a_e[4]), .Y(C1_Z_4) );
  scg2d1_hd U798 ( .A(n1120), .B(a[26]), .C(n1833), .D(a_e[3]), .Y(C1_Z_3) );
  scg2d1_hd U799 ( .A(n1120), .B(a[25]), .C(n1833), .D(a_e[2]), .Y(C1_Z_2) );
  scg2d1_hd U800 ( .A(n1120), .B(a[24]), .C(n1833), .D(a_e[1]), .Y(C1_Z_1) );
  scg2d1_hd U801 ( .A(n1120), .B(a[29]), .C(n1833), .D(a_e[6]), .Y(C1_Z_6) );
  nr2d2_hd U802 ( .A(n1234), .B(n1233), .Y(n1867) );
  scg2d1_hd U803 ( .A(n1388), .B(n1888), .C(n1024), .D(n1879), .Y(n1339) );
  nr2d2_hd U804 ( .A(n1226), .B(n1223), .Y(n1922) );
  nr2d2_hd U805 ( .A(n1238), .B(n1237), .Y(n1906) );
  nid4_hd U806 ( .A(n1113), .Y(n1010) );
  xo2d1_hd U807 ( .A(n1939), .B(n1444), .Y(intadd_33_B_1_) );
  nr2d2_hd U808 ( .A(n1096), .B(n1095), .Y(n1411) );
  xo2d1_hd U809 ( .A(n1892), .B(n1457), .Y(intadd_36_A_2_) );
  xo2d1_hd U810 ( .A(a_m[17]), .B(n1449), .Y(intadd_34_B_1_) );
  nr2d2_hd U811 ( .A(n1088), .B(n1087), .Y(n1291) );
  ivd2_hd U812 ( .A(n1699), .Y(n1710) );
  ivd4_hd U813 ( .A(n1007), .Y(n1120) );
  nr2d2_hd U814 ( .A(n1356), .B(n1239), .Y(n1904) );
  nr2d2_hd U815 ( .A(n1338), .B(n1220), .Y(n1920) );
  or4d1_hd U816 ( .A(n1768), .B(n1760), .C(n1842), .D(b_e[4]), .Y(n1522) );
  or4d1_hd U817 ( .A(product[3]), .B(product[10]), .C(product[11]), .D(
        product[6]), .Y(n1696) );
  clknd2d1_hd U818 ( .A(n1584), .B(n1564), .Y(n231) );
  clknd2d1_hd U819 ( .A(n1584), .B(n1571), .Y(n233) );
  oa21d2_hd U820 ( .A(n1749), .B(n1808), .C(n1007), .Y(n1754) );
  ao21d2_hd U821 ( .A(n1836), .B(n1741), .C(n1786), .Y(n1749) );
  scg2d1_hd U822 ( .A(z_e[1]), .B(n1844), .C(n1113), .D(
        DP_OP_125J3_130_6300_n35), .Y(DP_OP_125J3_130_6300_n25) );
  scg2d1_hd U823 ( .A(z_e[2]), .B(n1844), .C(n1113), .D(
        DP_OP_125J3_130_6300_n36), .Y(DP_OP_125J3_130_6300_n26) );
  scg2d1_hd U824 ( .A(z_e[3]), .B(n1844), .C(n1010), .D(
        DP_OP_125J3_130_6300_n37), .Y(DP_OP_125J3_130_6300_n27) );
  scg2d1_hd U825 ( .A(z_e[4]), .B(n1844), .C(n1010), .D(
        DP_OP_125J3_130_6300_n38), .Y(DP_OP_125J3_130_6300_n28) );
  scg2d1_hd U826 ( .A(z_e[5]), .B(n1844), .C(n1010), .D(
        DP_OP_125J3_130_6300_n39), .Y(DP_OP_125J3_130_6300_n29) );
  oa21d2_hd U827 ( .A(state[1]), .B(n1806), .C(n1813), .Y(n1844) );
  nr2d2_hd U828 ( .A(n1062), .B(n1802), .Y(n1179) );
  scg2d1_hd U829 ( .A(z_m[0]), .B(n1590), .C(n1016), .D(z[0]), .Y(n260) );
  scg2d1_hd U830 ( .A(z_m[1]), .B(n1590), .C(n1016), .D(z[1]), .Y(n259) );
  scg2d1_hd U831 ( .A(z_m[2]), .B(n1590), .C(n1016), .D(z[2]), .Y(n258) );
  scg2d1_hd U832 ( .A(z_m[3]), .B(n1590), .C(n1016), .D(z[3]), .Y(n257) );
  scg2d1_hd U833 ( .A(z_m[4]), .B(n1590), .C(n1016), .D(z[4]), .Y(n256) );
  nr2d4_hd U834 ( .A(n1587), .B(n1586), .Y(n1590) );
  nr2ad1_hd U835 ( .A(n1705), .B(n1813), .Y(n1711) );
  clknd2d2_hd U836 ( .A(n1495), .B(n1803), .Y(n1007) );
  oa211d2_hd U837 ( .A(n1717), .B(n1500), .C(n1499), .D(n1498), .Y(n110) );
  nr2ad1_hd U838 ( .A(n1591), .B(n105), .Y(n1705) );
  ivd2_hd U839 ( .A(n1028), .Y(n1027) );
  ivd1_hd U840 ( .A(b_m[4]), .Y(n1029) );
  nid2_hd U841 ( .A(b_m[5]), .Y(n1030) );
  scg4d1_hd U842 ( .A(n1055), .B(n1906), .C(n1053), .D(n1904), .E(n1051), .F(
        n1905), .G(n1903), .H(intadd_24_SUM_17_), .Y(n1462) );
  ivd1_hd U843 ( .A(n1929), .Y(n1407) );
  nid2_hd U844 ( .A(b_m[6]), .Y(n1031) );
  ivd1_hd U845 ( .A(n1808), .Y(n1833) );
  ivd1_hd U846 ( .A(n1762), .Y(n1850) );
  ivd1_hd U847 ( .A(n1813), .Y(n1112) );
  nid2_hd U848 ( .A(n359), .Y(n1023) );
  ivd1_hd U849 ( .A(n1711), .Y(n1708) );
  ivd1_hd U850 ( .A(n1767), .Y(n1838) );
  ivd1_hd U851 ( .A(n1765), .Y(n1843) );
  scg6d1_hd U852 ( .A(n1850), .B(n1059), .C(n1120), .Y(n1015) );
  nid2_hd U853 ( .A(n1703), .Y(n1017) );
  ivd1_hd U854 ( .A(n105), .Y(n1701) );
  ivd1_hd U855 ( .A(n1709), .Y(n1684) );
  ivd1_hd U856 ( .A(n1498), .Y(n1113) );
  ivd1_hd U857 ( .A(n1820), .Y(n1809) );
  ivd1_hd U858 ( .A(n1875), .Y(n2034) );
  ivd1_hd U859 ( .A(n1887), .Y(n2032) );
  ivd1_hd U860 ( .A(intadd_32_n1), .Y(n1186) );
  ivd1_hd U861 ( .A(intadd_36_n1), .Y(n1188) );
  nid2_hd U862 ( .A(n1882), .Y(n1020) );
  ivd1_hd U863 ( .A(n1865), .Y(n2036) );
  ivd2_hd U864 ( .A(n1015), .Y(n1018) );
  clknd2d2_hd U865 ( .A(n1850), .B(n1015), .Y(n1740) );
  ivd2_hd U866 ( .A(n1013), .Y(n1016) );
  ivd1_hd U867 ( .A(n1586), .Y(n1551) );
  ivd1_hd U868 ( .A(n1749), .Y(n1759) );
  clknd2d2_hd U869 ( .A(n1833), .B(n1061), .Y(n1832) );
  ivd1_hd U870 ( .A(n1543), .Y(n1552) );
  ao21d1_hd U871 ( .A(n1743), .B(n1741), .C(n1015), .Y(n1765) );
  nr2d1_hd U872 ( .A(n1547), .B(n1543), .Y(n1741) );
  nr2d1_hd U873 ( .A(n1504), .B(n1503), .Y(n1836) );
  nr2d1_hd U874 ( .A(n1701), .B(n1818), .Y(n1703) );
  nr2ad1_hd U875 ( .A(n1705), .B(n1610), .Y(n1709) );
  ivd1_hd U876 ( .A(n1601), .Y(n1600) );
  ivd1_hd U877 ( .A(n1611), .Y(n1609) );
  ivd1_hd U878 ( .A(n1620), .Y(n1619) );
  ivd1_hd U879 ( .A(n1629), .Y(n1628) );
  ivd1_hd U880 ( .A(n1638), .Y(n1637) );
  scg14d1_hd U881 ( .A(n1388), .B(n1176), .C(n1063), .Y(n1065) );
  nid2_hd U882 ( .A(n1793), .Y(n1019) );
  ivd1_hd U883 ( .A(n1169), .Y(n1095) );
  ad2d2_hd U884 ( .A(n1281), .B(n1280), .Y(n1934) );
  nid2_hd U885 ( .A(n1914), .Y(n1021) );
  ivd1_hd U886 ( .A(intadd_38_SUM_2_), .Y(n1183) );
  ivd1_hd U887 ( .A(n1883), .Y(n2033) );
  ivd1_hd U888 ( .A(a_m[12]), .Y(n1781) );
  ivd1_hd U889 ( .A(intadd_37_SUM_2_), .Y(n1181) );
  ivd1_hd U890 ( .A(n1896), .Y(n2030) );
  ivd1_hd U891 ( .A(intadd_32_SUM_5_), .Y(n1187) );
  ivd1_hd U892 ( .A(n1899), .Y(n2029) );
  ivd1_hd U893 ( .A(a_m[19]), .Y(n1771) );
  ivd1_hd U894 ( .A(a_m[18]), .Y(n1773) );
  ivd1_hd U895 ( .A(a_m[17]), .Y(n1882) );
  ivd1_hd U896 ( .A(n1861), .Y(n2037) );
  ivd1_hd U897 ( .A(n1356), .Y(n1237) );
  ivd1_hd U898 ( .A(n1741), .Y(n1835) );
  scg17d1_hd U899 ( .A(z_m[6]), .B(n1711), .C(n1663), .D(n1662), .Y(n276) );
  ivd1_hd U900 ( .A(n1578), .Y(n1585) );
  ao21d1_hd U901 ( .A(n1558), .B(n1557), .C(n1586), .Y(n1578) );
  ao22d1_hd U902 ( .A(n1553), .B(n1552), .C(n1587), .D(n1551), .Y(n1584) );
  scg20d1_hd U903 ( .A(z_e[7]), .B(z_e[8]), .C(z_e[9]), .Y(n1587) );
  scg17d1_hd U904 ( .A(z_m[14]), .B(n1711), .C(n1627), .D(n1626), .Y(n268) );
  ivd2_hd U905 ( .A(n1786), .Y(n1830) );
  scg17d1_hd U906 ( .A(z_m[10]), .B(n1711), .C(n1645), .D(n1644), .Y(n272) );
  scg17d1_hd U907 ( .A(z_m[2]), .B(n1711), .C(n1682), .D(n1681), .Y(n280) );
  scg2d1_hd U908 ( .A(state[0]), .B(n1829), .C(n1828), .D(n1827), .Y(n353) );
  nr2d1_hd U909 ( .A(n1806), .B(n1820), .Y(n359) );
  scg17d1_hd U910 ( .A(z_m[18]), .B(n1711), .C(n1608), .D(n1607), .Y(n264) );
  oa21d1_hd U911 ( .A(n1120), .B(n1850), .C(n1843), .Y(n1767) );
  nr2d1_hd U912 ( .A(state[2]), .B(state[3]), .Y(n1803) );
  nd3d1_hd U913 ( .A(n1550), .B(n1537), .C(n1535), .Y(n1547) );
  nr2d1_hd U914 ( .A(n1522), .B(n1521), .Y(n1743) );
  ivd1_hd U915 ( .A(b_e[8]), .Y(n1760) );
  ivd1_hd U916 ( .A(b_e[0]), .Y(n1768) );
  scg17d1_hd U917 ( .A(z_m[20]), .B(n1711), .C(n1599), .D(n1598), .Y(n262) );
  nr2d1_hd U918 ( .A(state[0]), .B(n1825), .Y(n1545) );
  ivd1_hd U919 ( .A(state[1]), .Y(n1825) );
  ivd1_hd U920 ( .A(a_e[9]), .Y(n1758) );
  ivd1_hd U921 ( .A(b_e[9]), .Y(n1842) );
  ivd1_hd U922 ( .A(n1546), .Y(n1806) );
  ivd1_hd U923 ( .A(z_m[23]), .Y(n1814) );
  nr2d1_hd U924 ( .A(n1822), .B(state[3]), .Y(n1821) );
  ivd1_hd U925 ( .A(state[2]), .Y(n1822) );
  nr2d1_hd U926 ( .A(state[2]), .B(n1846), .Y(n1546) );
  ivd1_hd U927 ( .A(state[3]), .Y(n1846) );
  ivd1_hd U928 ( .A(z_m[0]), .Y(n1496) );
  ivd1_hd U929 ( .A(a_m[0]), .Y(n1802) );
  ivd1_hd U930 ( .A(a_m[1]), .Y(n1800) );
  ad2d2_hd U931 ( .A(n1515), .B(a_m[2]), .Y(n1178) );
  ivd1_hd U932 ( .A(a_m[7]), .Y(n1789) );
  ivd1_hd U933 ( .A(a_m[5]), .Y(n1793) );
  ivd1_hd U934 ( .A(a_m[6]), .Y(n1791) );
  ivd1_hd U935 ( .A(n1066), .Y(n1071) );
  fad1_hd U936 ( .A(n1874), .B(n1873), .CI(n1872), .CO(n1875), .S(n1871) );
  ivd1_hd U937 ( .A(a_m[10]), .Y(n1783) );
  ivd1_hd U938 ( .A(a_m[9]), .Y(n1785) );
  ivd1_hd U939 ( .A(a_m[2]), .Y(n1914) );
  fad1_hd U940 ( .A(n1886), .B(n1885), .CI(n1884), .CO(n1887), .S(n1883) );
  ivd1_hd U941 ( .A(a_m[13]), .Y(n1779) );
  ivd1_hd U942 ( .A(a_m[15]), .Y(n1777) );
  ivd1_hd U943 ( .A(a_m[16]), .Y(n1775) );
  fad1_hd U944 ( .A(intadd_36_SUM_1_), .B(n1901), .CI(n1900), .CO(n1902), .S(
        n1899) );
  ivd2_hd U945 ( .A(a_m[20]), .Y(n1892) );
  fad1_hd U946 ( .A(n1864), .B(n1863), .CI(n1862), .CO(n1865), .S(n1861) );
  nr2d1_hd U947 ( .A(state[1]), .B(state[0]), .Y(n1810) );
  nr2d1_hd U948 ( .A(n1802), .B(n1014), .Y(N176) );
  ivd2_hd U949 ( .A(n1409), .Y(n1289) );
  ivd2_hd U950 ( .A(n1488), .Y(n1931) );
  ivd2_hd U951 ( .A(n1477), .Y(n1935) );
  ivd2_hd U952 ( .A(n1471), .Y(n1877) );
  ivd2_hd U953 ( .A(n1451), .Y(n1921) );
  ivd2_hd U954 ( .A(n1859), .Y(n1905) );
  nr2d1_hd U955 ( .A(n1061), .B(n1056), .Y(n1863) );
  ad2d2_hd U956 ( .A(n1234), .B(n1284), .Y(n1876) );
  ad2d2_hd U957 ( .A(n1332), .B(n1228), .Y(n1888) );
  nr2d1_hd U958 ( .A(n1022), .B(n1025), .Y(n1066) );
  oa21d1_hd U959 ( .A(n1014), .B(n1024), .C(n1071), .Y(n1388) );
  ao22d1_hd U960 ( .A(a_m[2]), .B(a_m[1]), .C(n1800), .D(n1914), .Y(n1062) );
  ao22d1_hd U961 ( .A(n1022), .B(n1177), .C(n1024), .D(n1179), .Y(n1063) );
  nr3d1_hd U962 ( .A(N176), .B(n1065), .C(n1021), .Y(n1069) );
  nr2d1_hd U963 ( .A(a_m[0]), .B(a_m[1]), .Y(n1515) );
  ao22d1_hd U964 ( .A(n1012), .B(n1066), .C(n1071), .D(n1026), .Y(n1386) );
  scg4d1_hd U965 ( .A(n1022), .B(n1178), .C(n1024), .D(n1177), .E(n1386), .F(
        n1176), .G(n1179), .H(n1012), .Y(n1067) );
  nr2d1_hd U966 ( .A(a_m[3]), .B(a_m[2]), .Y(n1510) );
  ao21d1_hd U967 ( .A(a_m[2]), .B(a_m[3]), .C(n1510), .Y(n1086) );
  oa211d1_hd U968 ( .A(n1025), .B(n1026), .C(n1524), .D(n1071), .Y(n1072) );
  scg4d1_hd U969 ( .A(n1027), .B(n1179), .C(n1024), .D(n1178), .E(n1177), .F(
        n1012), .G(n1396), .H(n1176), .Y(n1073) );
  nr2d1_hd U970 ( .A(n1057), .B(n1056), .Y(n1114) );
  nr2d1_hd U971 ( .A(n1061), .B(n1114), .Y(n1077) );
  nr2d1_hd U972 ( .A(a_m[21]), .B(a_m[20]), .Y(n1509) );
  ao21d1_hd U973 ( .A(a_m[20]), .B(a_m[21]), .C(n1509), .Y(n1356) );
  nr2d1_hd U974 ( .A(a_m[23]), .B(a_m[22]), .Y(n1512) );
  ao21d1_hd U975 ( .A(a_m[22]), .B(n1060), .C(n1512), .Y(n1238) );
  nd3d1_hd U976 ( .A(n1239), .B(n1237), .C(n1238), .Y(n1859) );
  oa22d1_hd U977 ( .A(n1059), .B(n1859), .C(n1240), .D(n1407), .Y(n1219) );
  oa22d1_hd U978 ( .A(n1077), .B(n1219), .C(n1061), .D(n1076), .Y(n1079) );
  oa22ad1_hd U979 ( .A(n1061), .B(n1525), .C(b_m[23]), .D(n1863), .Y(n1078) );
  ao22d1_hd U980 ( .A(a_e[9]), .B(b_e[9]), .C(n1842), .D(n1758), .Y(n1081) );
  nr2d1_hd U981 ( .A(DP_OP_125J3_130_6300_n12), .B(n1081), .Y(n1080) );
  ao211d1_hd U982 ( .A(DP_OP_125J3_130_6300_n12), .B(n1081), .C(n1498), .D(
        n1080), .Y(n1082) );
  ao21d1_hd U983 ( .A(z_e[9]), .B(n1844), .C(n1082), .Y(n1083) );
  ivd1_hd U984 ( .A(n1086), .Y(n1087) );
  ivd1_hd U985 ( .A(a_m[4]), .Y(n1795) );
  ivd1_hd U986 ( .A(a_m[3]), .Y(n1797) );
  oa22d1_hd U987 ( .A(n1795), .B(n1797), .C(a_m[3]), .D(a_m[4]), .Y(n1085) );
  nr2d1_hd U988 ( .A(a_m[5]), .B(a_m[4]), .Y(n1511) );
  ao21d1_hd U989 ( .A(a_m[4]), .B(a_m[5]), .C(n1511), .Y(n1088) );
  nd3d1_hd U990 ( .A(n1087), .B(n1085), .C(n1088), .Y(n1409) );
  scg4d1_hd U991 ( .A(n1022), .B(n1289), .C(n1024), .D(n1292), .E(n1386), .F(
        n1290), .G(n1012), .H(n1291), .Y(n1163) );
  ao21d1_hd U992 ( .A(n1022), .B(n1292), .C(n1089), .Y(n1216) );
  nd3d1_hd U993 ( .A(n1216), .B(a_m[5]), .C(n1211), .Y(n1159) );
  oa211d1_hd U994 ( .A(n1055), .B(intadd_24_n1), .C(n1057), .D(n1059), .Y(
        n1091) );
  ao22d1_hd U995 ( .A(b_m[23]), .B(n1292), .C(n1290), .D(n1857), .Y(n1092) );
  oa21d1_hd U996 ( .A(n1409), .B(n1058), .C(n1092), .Y(n1093) );
  ao22d1_hd U997 ( .A(a_m[8]), .B(a_m[7]), .C(n1789), .D(n1787), .Y(n1096) );
  ao22d1_hd U998 ( .A(a_m[5]), .B(a_m[6]), .C(n1791), .D(n1793), .Y(n1169) );
  nr2d1_hd U999 ( .A(a_m[7]), .B(a_m[6]), .Y(n1513) );
  scg6d1_hd U1000 ( .A(a_m[6]), .B(a_m[7]), .C(n1513), .Y(n1094) );
  nd3d1_hd U1001 ( .A(n1095), .B(n1094), .C(n1096), .Y(n1488) );
  scg4d1_hd U1002 ( .A(n1055), .B(n1411), .C(n1053), .D(n1486), .E(n1051), .F(
        n1931), .G(n1930), .H(intadd_24_SUM_17_), .Y(n1097) );
  fad1_hd U1003 ( .A(intadd_26_SUM_14_), .B(n1099), .CI(n1098), .CO(
        intadd_21_A_24_), .S(intadd_21_A_23_) );
  scg4d1_hd U1004 ( .A(n1011), .B(n1178), .C(n1031), .D(n1179), .E(n1030), .F(
        n1177), .G(n1176), .H(intadd_24_SUM_2_), .Y(n1100) );
  scg4d1_hd U1005 ( .A(n1011), .B(n1179), .C(n1012), .D(n1178), .E(n1177), .F(
        n1027), .G(n1176), .H(intadd_24_SUM_0_), .Y(n1101) );
  scg4d1_hd U1006 ( .A(n1043), .B(n1179), .C(n1040), .D(n1178), .E(n1177), .F(
        n1041), .G(n1176), .H(intadd_24_SUM_10_), .Y(n1102) );
  scg4d1_hd U1007 ( .A(n1044), .B(n1179), .C(n1041), .D(n1178), .E(n1177), .F(
        n1043), .G(n1176), .H(intadd_24_SUM_11_), .Y(n1103) );
  scg4d1_hd U1008 ( .A(n1046), .B(n1179), .C(n1043), .D(n1178), .E(n1177), .F(
        n1044), .G(n1176), .H(intadd_24_SUM_12_), .Y(n1104) );
  scg4d1_hd U1009 ( .A(n1048), .B(n1179), .C(n1044), .D(n1178), .E(n1177), .F(
        n1046), .G(n1176), .H(intadd_24_SUM_13_), .Y(n1105) );
  scg4d1_hd U1010 ( .A(n1048), .B(n1177), .C(n1050), .D(n1179), .E(n1178), .F(
        n1046), .G(n1176), .H(intadd_24_SUM_14_), .Y(n1107) );
  scg4d1_hd U1011 ( .A(n1048), .B(n1178), .C(n1050), .D(n1177), .E(n1051), .F(
        n1179), .G(n1176), .H(intadd_24_SUM_15_), .Y(n1108) );
  scg4d1_hd U1012 ( .A(n1051), .B(n1177), .C(n1050), .D(n1178), .E(n1053), .F(
        n1179), .G(n1176), .H(intadd_24_SUM_16_), .Y(n1109) );
  scg4d1_hd U1013 ( .A(n1055), .B(n1179), .C(n1053), .D(n1177), .E(n1178), .F(
        n1051), .G(n1176), .H(intadd_24_SUM_17_), .Y(n1110) );
  nd2bd1_hd U1014 ( .AN(n1114), .B(n1111), .Y(n1217) );
  scg4d1_hd U1015 ( .A(n1937), .B(n1176), .C(n1055), .D(n1177), .E(n1179), .F(
        n1057), .G(n1178), .H(n1053), .Y(n1115) );
  oa21d1_hd U1016 ( .A(intadd_24_n1), .B(n1055), .C(n1057), .Y(n1116) );
  scg4d1_hd U1017 ( .A(n1057), .B(n1177), .C(b_m[23]), .D(n1179), .E(n1178), 
        .F(n1055), .G(n1176), .H(n1460), .Y(n1123) );
  scg4d1_hd U1018 ( .A(n1011), .B(n1177), .C(n1027), .D(n1178), .E(n1030), .F(
        n1179), .G(n1176), .H(intadd_24_SUM_1_), .Y(n1124) );
  ao21d1_hd U1019 ( .A(n1515), .B(n1057), .C(n1021), .Y(n1146) );
  mx2id1_hd U1020 ( .D0(n1146), .D1(n1021), .S(n1144), .YN(intadd_21_B_20_) );
  ao22d1_hd U1021 ( .A(b_m[23]), .B(n1178), .C(n1176), .D(n1929), .Y(n1155) );
  nr2d1_hd U1022 ( .A(n1150), .B(n1407), .Y(n1153) );
  ao22d1_hd U1023 ( .A(a_m[2]), .B(n1155), .C(n1153), .D(n1021), .Y(
        intadd_21_B_21_) );
  nr2d1_hd U1024 ( .A(n1163), .B(n1159), .Y(n1243) );
  scg4d1_hd U1025 ( .A(n1027), .B(n1291), .C(n1024), .D(n1289), .E(n1292), .F(
        n1012), .G(n1396), .H(n1290), .Y(n1167) );
  xo3d1_hd U1026 ( .A(n1243), .B(n1242), .C(n1268), .Y(intadd_21_B_2_) );
  scg4d1_hd U1027 ( .A(n1030), .B(n1178), .C(n1031), .D(n1177), .E(n1032), .F(
        n1179), .G(n1176), .H(intadd_24_SUM_3_), .Y(n1170) );
  scg4d1_hd U1028 ( .A(n1034), .B(n1179), .C(n1031), .D(n1178), .E(n1177), .F(
        n1032), .G(n1176), .H(intadd_24_SUM_4_), .Y(n1171) );
  scg4d1_hd U1029 ( .A(n1034), .B(n1177), .C(n1036), .D(n1179), .E(n1178), .F(
        n1032), .G(n1176), .H(intadd_24_SUM_5_), .Y(n1172) );
  scg4d1_hd U1030 ( .A(n1034), .B(n1178), .C(n1037), .D(n1179), .E(n1036), .F(
        n1177), .G(n1176), .H(intadd_24_SUM_6_), .Y(n1173) );
  scg4d1_hd U1031 ( .A(n1039), .B(n1179), .C(n1037), .D(n1177), .E(n1178), .F(
        n1036), .G(n1176), .H(intadd_24_SUM_7_), .Y(n1174) );
  scg4d1_hd U1032 ( .A(n1040), .B(n1179), .C(n1037), .D(n1178), .E(n1177), .F(
        n1039), .G(n1176), .H(intadd_24_SUM_8_), .Y(n1175) );
  scg4d1_hd U1033 ( .A(n1041), .B(n1179), .C(n1039), .D(n1178), .E(n1177), .F(
        n1040), .G(n1176), .H(intadd_24_SUM_9_), .Y(n1202) );
  nr2d1_hd U1034 ( .A(n1019), .B(n1211), .Y(n1214) );
  nr2d1_hd U1035 ( .A(n1061), .B(n1028), .Y(intadd_22_B_0_) );
  nr2d1_hd U1036 ( .A(n1061), .B(n1217), .Y(n1218) );
  oa22d1_hd U1037 ( .A(n1771), .B(a_m[20]), .C(n1892), .D(a_m[19]), .Y(n1226)
         );
  ao22d1_hd U1038 ( .A(a_m[17]), .B(a_m[18]), .C(n1773), .D(n1882), .Y(n1338)
         );
  ivd1_hd U1039 ( .A(n1338), .Y(n1223) );
  oa22d1_hd U1040 ( .A(n1771), .B(n1773), .C(a_m[18]), .D(a_m[19]), .Y(n1220)
         );
  nd3d1_hd U1041 ( .A(n1223), .B(n1220), .C(n1226), .Y(n1451) );
  scg4d1_hd U1042 ( .A(n1039), .B(n1922), .C(n1037), .D(n1920), .E(n1036), .F(
        n1921), .G(n1919), .H(intadd_24_SUM_7_), .Y(n1227) );
  nr2d1_hd U1043 ( .A(a_m[15]), .B(a_m[14]), .Y(n1514) );
  ao21d1_hd U1044 ( .A(a_m[14]), .B(a_m[15]), .C(n1514), .Y(n1332) );
  oa22d1_hd U1045 ( .A(n1775), .B(a_m[17]), .C(n1882), .D(a_m[16]), .Y(n1228)
         );
  oa22d1_hd U1046 ( .A(n1775), .B(n1777), .C(a_m[15]), .D(a_m[16]), .Y(n1229)
         );
  scg4d1_hd U1047 ( .A(n1044), .B(n1879), .C(n1041), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_11_), .G(n1043), .H(n1880), .Y(n1230) );
  scg4d1_hd U1048 ( .A(n1048), .B(n1879), .C(n1044), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_13_), .G(n1046), .H(n1880), .Y(n1231) );
  oa22d1_hd U1049 ( .A(n1779), .B(a_m[14]), .C(n1870), .D(a_m[13]), .Y(n1234)
         );
  ao22d1_hd U1050 ( .A(a_m[11]), .B(a_m[12]), .C(n1781), .D(n1939), .Y(n1284)
         );
  ivd1_hd U1051 ( .A(n1284), .Y(n1233) );
  oa22d1_hd U1052 ( .A(n1779), .B(n1781), .C(a_m[12]), .D(a_m[13]), .Y(n1232)
         );
  nd3d1_hd U1053 ( .A(n1233), .B(n1232), .C(n1234), .Y(n1471) );
  scg4d1_hd U1054 ( .A(n1055), .B(n1867), .C(n1053), .D(n1868), .E(n1051), .F(
        n1877), .G(n1876), .H(intadd_24_SUM_17_), .Y(n1235) );
  scg4d1_hd U1055 ( .A(n1057), .B(n1868), .C(b_m[23]), .D(n1867), .E(n1055), 
        .F(n1877), .G(n1876), .H(n1460), .Y(n1236) );
  scg4d1_hd U1056 ( .A(n1011), .B(n1905), .C(n1031), .D(n1906), .E(n1904), .F(
        n1030), .G(n1903), .H(intadd_24_SUM_2_), .Y(n1241) );
  scg16d1_hd U1057 ( .A(n1268), .B(n1243), .C(n1242), .Y(intadd_23_A_0_) );
  scg4d1_hd U1058 ( .A(n1043), .B(n1291), .C(n1040), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_10_), .G(n1041), .H(n1292), .Y(n1244) );
  scg4d1_hd U1059 ( .A(n1048), .B(n1291), .C(n1044), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_13_), .G(n1046), .H(n1292), .Y(n1245) );
  scg4d1_hd U1060 ( .A(n1937), .B(n1290), .C(n1055), .D(n1292), .E(n1291), .F(
        n1057), .G(n1289), .H(n1053), .Y(n1246) );
  scg4d1_hd U1061 ( .A(n1011), .B(n1292), .C(n1027), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_1_), .G(n1291), .H(n1030), .Y(n1247) );
  scg4d1_hd U1062 ( .A(n1027), .B(n1411), .C(n1024), .D(n1931), .E(n1396), .F(
        n1930), .G(n1486), .H(n1012), .Y(n1248) );
  ao22d1_hd U1063 ( .A(a_m[8]), .B(n1785), .C(a_m[9]), .D(n1787), .Y(n1279) );
  ivd1_hd U1064 ( .A(n1279), .Y(n1280) );
  scg4d1_hd U1065 ( .A(n1022), .B(n1931), .C(n1024), .D(n1486), .E(n1012), .F(
        n1411), .G(n1386), .H(n1930), .Y(n1259) );
  ao21d1_hd U1066 ( .A(n1022), .B(n1486), .C(n1249), .Y(n1270) );
  nd3d1_hd U1067 ( .A(a_m[8]), .B(n1270), .C(n1268), .Y(n1257) );
  nr2d1_hd U1068 ( .A(n1259), .B(n1257), .Y(n1273) );
  xo3d1_hd U1069 ( .A(n1272), .B(n1305), .C(n1273), .Y(intadd_23_A_2_) );
  scg4d1_hd U1070 ( .A(n1011), .B(n1291), .C(n1012), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_0_), .G(n1027), .H(n1292), .Y(n1250) );
  scg4d1_hd U1071 ( .A(n1044), .B(n1291), .C(n1041), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_11_), .G(n1043), .H(n1292), .Y(n1251) );
  scg4d1_hd U1072 ( .A(n1046), .B(n1291), .C(n1043), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_12_), .G(n1044), .H(n1292), .Y(n1252) );
  scg4d1_hd U1073 ( .A(n1048), .B(n1292), .C(n1050), .D(n1291), .E(n1290), .F(
        intadd_24_SUM_14_), .G(n1046), .H(n1289), .Y(n1253) );
  scg4d1_hd U1074 ( .A(n1048), .B(n1289), .C(n1050), .D(n1292), .E(n1290), .F(
        intadd_24_SUM_15_), .G(n1291), .H(n1051), .Y(n1254) );
  scg4d1_hd U1075 ( .A(n1051), .B(n1292), .C(n1050), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_16_), .G(n1291), .H(n1053), .Y(n1255) );
  scg4d1_hd U1076 ( .A(n1055), .B(n1291), .C(n1053), .D(n1292), .E(n1290), .F(
        intadd_24_SUM_17_), .G(n1051), .H(n1289), .Y(n1256) );
  scg4d1_hd U1077 ( .A(n1011), .B(n1289), .C(n1031), .D(n1291), .E(n1290), .F(
        intadd_24_SUM_2_), .G(n1292), .H(n1030), .Y(n1260) );
  scg4d1_hd U1078 ( .A(n1030), .B(n1289), .C(n1031), .D(n1292), .E(n1290), .F(
        intadd_24_SUM_3_), .G(n1291), .H(n1032), .Y(n1261) );
  scg4d1_hd U1079 ( .A(n1034), .B(n1291), .C(n1031), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_4_), .G(n1032), .H(n1292), .Y(n1262) );
  scg4d1_hd U1080 ( .A(n1034), .B(n1292), .C(n1036), .D(n1291), .E(n1290), .F(
        intadd_24_SUM_5_), .G(n1032), .H(n1289), .Y(n1263) );
  scg4d1_hd U1081 ( .A(n1034), .B(n1289), .C(n1037), .D(n1291), .E(n1290), .F(
        intadd_24_SUM_6_), .G(n1292), .H(n1036), .Y(n1264) );
  scg4d1_hd U1082 ( .A(n1039), .B(n1291), .C(n1037), .D(n1292), .E(n1290), .F(
        intadd_24_SUM_7_), .G(n1036), .H(n1289), .Y(n1265) );
  scg4d1_hd U1083 ( .A(n1040), .B(n1291), .C(n1037), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_8_), .G(n1039), .H(n1292), .Y(n1266) );
  scg4d1_hd U1084 ( .A(n1041), .B(n1291), .C(n1039), .D(n1289), .E(n1290), .F(
        intadd_24_SUM_9_), .G(n1040), .H(n1292), .Y(n1267) );
  nr2d1_hd U1085 ( .A(n1787), .B(n1268), .Y(n1269) );
  oa22d1_hd U1086 ( .A(n1271), .B(n1028), .C(n1026), .D(n1025), .Y(
        intadd_24_CI) );
  scg16d1_hd U1087 ( .A(n1305), .B(n1273), .C(n1272), .Y(intadd_25_A_0_) );
  scg4d1_hd U1088 ( .A(n1043), .B(n1411), .C(n1040), .D(n1931), .E(n1041), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_10_), .Y(n1274) );
  scg4d1_hd U1089 ( .A(n1048), .B(n1411), .C(n1044), .D(n1931), .E(n1046), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_13_), .Y(n1275) );
  scg4d1_hd U1090 ( .A(n1048), .B(n1931), .C(n1050), .D(n1486), .E(n1411), .F(
        n1051), .G(n1930), .H(intadd_24_SUM_15_), .Y(n1276) );
  scg4d1_hd U1091 ( .A(n1011), .B(n1486), .C(n1027), .D(n1931), .E(n1411), .F(
        n1030), .G(n1930), .H(intadd_24_SUM_1_), .Y(n1277) );
  nr2d1_hd U1092 ( .A(a_m[10]), .B(a_m[9]), .Y(n1516) );
  ao21d1_hd U1093 ( .A(a_m[9]), .B(a_m[10]), .C(n1516), .Y(n1278) );
  ao22d1_hd U1094 ( .A(a_m[11]), .B(n1783), .C(a_m[10]), .D(n1939), .Y(n1281)
         );
  nr3d1_hd U1095 ( .A(n1280), .B(n1278), .C(n1281), .Y(n1933) );
  scg4d1_hd U1096 ( .A(n1022), .B(n1009), .C(n1024), .D(n1935), .E(n1386), .F(
        n1936), .G(n1012), .H(n1934), .Y(n1296) );
  ao21d1_hd U1097 ( .A(n1024), .B(n1934), .C(n1282), .Y(n1307) );
  nd3d1_hd U1098 ( .A(a_m[11]), .B(n1307), .C(n1305), .Y(n1294) );
  nr2d1_hd U1099 ( .A(n1296), .B(n1294), .Y(n1309) );
  scg4d1_hd U1100 ( .A(n1027), .B(n1934), .C(n1024), .D(n1009), .E(n1935), .F(
        n1012), .G(n1396), .H(n1936), .Y(n1283) );
  xo3d1_hd U1101 ( .A(n1309), .B(n1308), .C(n1335), .Y(intadd_25_A_2_) );
  scg4d1_hd U1102 ( .A(n1011), .B(n1411), .C(n1012), .D(n1931), .E(n1027), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_0_), .Y(n1285) );
  scg4d1_hd U1103 ( .A(n1044), .B(n1411), .C(n1041), .D(n1931), .E(n1043), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_11_), .Y(n1286) );
  scg4d1_hd U1104 ( .A(n1046), .B(n1411), .C(n1043), .D(n1931), .E(n1044), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_12_), .Y(n1287) );
  scg4d1_hd U1105 ( .A(n1048), .B(n1486), .C(n1050), .D(n1411), .E(n1931), .F(
        n1046), .G(n1930), .H(intadd_24_SUM_14_), .Y(n1288) );
  scg4d1_hd U1106 ( .A(n1057), .B(n1292), .C(b_m[23]), .D(n1291), .E(n1290), 
        .F(n1460), .G(n1055), .H(n1289), .Y(n1293) );
  scg4d1_hd U1107 ( .A(n1011), .B(n1931), .C(n1031), .D(n1411), .E(n1030), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_2_), .Y(n1297) );
  scg4d1_hd U1108 ( .A(n1030), .B(n1931), .C(n1031), .D(n1486), .E(n1411), .F(
        n1032), .G(n1930), .H(intadd_24_SUM_3_), .Y(n1298) );
  scg4d1_hd U1109 ( .A(n1034), .B(n1411), .C(n1031), .D(n1931), .E(n1032), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_4_), .Y(n1299) );
  scg4d1_hd U1110 ( .A(n1034), .B(n1486), .C(n1036), .D(n1411), .E(n1931), .F(
        n1032), .G(n1930), .H(intadd_24_SUM_5_), .Y(n1300) );
  scg4d1_hd U1111 ( .A(n1034), .B(n1931), .C(n1037), .D(n1411), .E(n1036), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_6_), .Y(n1301) );
  scg4d1_hd U1112 ( .A(n1039), .B(n1411), .C(n1037), .D(n1486), .E(n1036), .F(
        n1931), .G(n1930), .H(intadd_24_SUM_7_), .Y(n1302) );
  scg4d1_hd U1113 ( .A(n1040), .B(n1411), .C(n1037), .D(n1931), .E(n1039), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_8_), .Y(n1303) );
  scg4d1_hd U1114 ( .A(n1041), .B(n1411), .C(n1039), .D(n1931), .E(n1040), .F(
        n1486), .G(n1930), .H(intadd_24_SUM_9_), .Y(n1304) );
  nr2d1_hd U1115 ( .A(n1939), .B(n1305), .Y(n1306) );
  scg16d1_hd U1116 ( .A(n1335), .B(n1309), .C(n1308), .Y(intadd_26_A_0_) );
  scg4d1_hd U1117 ( .A(n1044), .B(n1934), .C(n1041), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_11_), .G(n1043), .H(n1935), .Y(n1310) );
  scg4d1_hd U1118 ( .A(n1051), .B(n1486), .C(n1050), .D(n1931), .E(n1411), .F(
        n1053), .G(n1930), .H(intadd_24_SUM_16_), .Y(n1311) );
  scg4d1_hd U1119 ( .A(n1011), .B(n1935), .C(n1027), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_1_), .G(n1934), .H(n1030), .Y(n1312) );
  scg4d1_hd U1120 ( .A(n1011), .B(n1009), .C(n1031), .D(n1934), .E(n1936), .F(
        intadd_24_SUM_2_), .G(n1935), .H(n1030), .Y(n1313) );
  scg4d1_hd U1121 ( .A(n1030), .B(n1009), .C(n1031), .D(n1935), .E(n1936), .F(
        intadd_24_SUM_3_), .G(n1934), .H(n1032), .Y(n1314) );
  scg4d1_hd U1122 ( .A(n1034), .B(n1934), .C(n1031), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_4_), .G(n1032), .H(n1935), .Y(n1315) );
  scg4d1_hd U1123 ( .A(n1034), .B(n1935), .C(n1036), .D(n1934), .E(n1936), .F(
        intadd_24_SUM_5_), .G(n1032), .H(n1009), .Y(n1316) );
  scg4d1_hd U1124 ( .A(n1034), .B(n1009), .C(n1037), .D(n1934), .E(n1936), .F(
        intadd_24_SUM_6_), .G(n1935), .H(n1036), .Y(n1317) );
  scg4d1_hd U1125 ( .A(n1039), .B(n1934), .C(n1037), .D(n1935), .E(n1936), .F(
        intadd_24_SUM_7_), .G(n1036), .H(n1009), .Y(n1318) );
  scg4d1_hd U1126 ( .A(n1041), .B(n1934), .C(n1039), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_9_), .G(n1040), .H(n1935), .Y(n1319) );
  scg4d1_hd U1127 ( .A(n1011), .B(n1934), .C(n1012), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_0_), .G(n1027), .H(n1935), .Y(n1320) );
  scg4d1_hd U1128 ( .A(n1043), .B(n1934), .C(n1040), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_10_), .G(n1041), .H(n1935), .Y(n1321) );
  scg4d1_hd U1129 ( .A(n1046), .B(n1934), .C(n1043), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_12_), .G(n1044), .H(n1935), .Y(n1322) );
  scg4d1_hd U1130 ( .A(n1048), .B(n1935), .C(n1050), .D(n1934), .E(n1936), .F(
        intadd_24_SUM_14_), .G(n1046), .H(n1009), .Y(n1323) );
  scg4d1_hd U1131 ( .A(n1044), .B(n1867), .C(n1041), .D(n1877), .E(n1868), .F(
        n1043), .G(n1876), .H(intadd_24_SUM_11_), .Y(n1324) );
  fad1_hd U1132 ( .A(intadd_27_SUM_8_), .B(n1326), .CI(n1325), .CO(
        intadd_26_B_15_), .S(intadd_26_B_14_) );
  scg4d1_hd U1133 ( .A(n1057), .B(n1486), .C(b_m[23]), .D(n1411), .E(n1931), 
        .F(n1055), .G(n1930), .H(n1460), .Y(n1327) );
  scg4d1_hd U1134 ( .A(n1022), .B(n1877), .C(n1024), .D(n1868), .E(n1867), .F(
        n1012), .G(n1386), .H(n1876), .Y(n1331) );
  ao21d1_hd U1135 ( .A(n1022), .B(n1868), .C(n1328), .Y(n1337) );
  nd3d1_hd U1136 ( .A(a_m[14]), .B(n1337), .C(n1335), .Y(n1330) );
  nr2d1_hd U1137 ( .A(n1331), .B(n1330), .Y(n1363) );
  scg4d1_hd U1138 ( .A(n1027), .B(n1867), .C(n1024), .D(n1877), .E(n1012), .F(
        n1868), .G(n1396), .H(n1876), .Y(n1333) );
  xo3d1_hd U1139 ( .A(n1363), .B(n1381), .C(n1362), .Y(intadd_26_B_2_) );
  scg4d1_hd U1140 ( .A(n1040), .B(n1934), .C(n1037), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_8_), .G(n1039), .H(n1935), .Y(n1334) );
  nr2d1_hd U1141 ( .A(n1870), .B(n1335), .Y(n1336) );
  scg4d1_hd U1142 ( .A(n1022), .B(n1889), .C(n1024), .D(n1880), .E(n1879), .F(
        n1012), .G(n1386), .H(n1888), .Y(n1376) );
  ao21d1_hd U1143 ( .A(n1022), .B(n1880), .C(n1339), .Y(n1383) );
  nd3d1_hd U1144 ( .A(a_m[17]), .B(n1383), .C(n1381), .Y(n1374) );
  nr2d1_hd U1145 ( .A(n1376), .B(n1374), .Y(n1379) );
  scg4d1_hd U1146 ( .A(n1027), .B(n1879), .C(n1024), .D(n1889), .E(n1012), .F(
        n1880), .G(n1888), .H(n1396), .Y(n1340) );
  scg16d1_hd U1147 ( .A(n1378), .B(n1379), .C(n1377), .Y(intadd_27_A_0_) );
  scg4d1_hd U1148 ( .A(n1048), .B(n1867), .C(n1044), .D(n1877), .E(n1868), .F(
        n1046), .G(n1876), .H(intadd_24_SUM_13_), .Y(n1341) );
  scg4d1_hd U1149 ( .A(n1022), .B(n1921), .C(n1024), .D(n1920), .E(n1919), .F(
        n1386), .G(n1922), .H(n1012), .Y(n1355) );
  ao21d1_hd U1150 ( .A(n1022), .B(n1920), .C(n1342), .Y(n1361) );
  nd3d1_hd U1151 ( .A(a_m[20]), .B(n1361), .C(n1378), .Y(n1354) );
  scg4d1_hd U1152 ( .A(n1011), .B(n1889), .C(n1031), .D(n1879), .E(n1888), .F(
        intadd_24_SUM_2_), .G(n1030), .H(n1880), .Y(n1344) );
  scg4d1_hd U1153 ( .A(n1030), .B(n1889), .C(n1031), .D(n1880), .E(n1888), .F(
        intadd_24_SUM_3_), .G(n1032), .H(n1879), .Y(n1345) );
  scg4d1_hd U1154 ( .A(n1034), .B(n1879), .C(n1031), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_4_), .G(n1032), .H(n1880), .Y(n1346) );
  scg4d1_hd U1155 ( .A(n1034), .B(n1880), .C(n1036), .D(n1879), .E(n1888), .F(
        intadd_24_SUM_5_), .G(n1889), .H(n1032), .Y(n1347) );
  scg4d1_hd U1156 ( .A(n1043), .B(n1867), .C(n1040), .D(n1877), .E(n1868), .F(
        n1041), .G(n1876), .H(intadd_24_SUM_10_), .Y(n1348) );
  scg4d1_hd U1157 ( .A(n1040), .B(n1879), .C(n1037), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_8_), .G(n1039), .H(n1880), .Y(n1349) );
  scg4d1_hd U1158 ( .A(n1011), .B(n1879), .C(n1012), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_0_), .G(n1027), .H(n1880), .Y(n1350) );
  scg4d1_hd U1159 ( .A(n1055), .B(n1934), .C(n1053), .D(n1935), .E(n1936), .F(
        intadd_24_SUM_17_), .G(n1051), .H(n1009), .Y(n1351) );
  scg4d1_hd U1160 ( .A(n1057), .B(n1935), .C(b_m[23]), .D(n1934), .E(n1936), 
        .F(n1460), .G(n1055), .H(n1009), .Y(n1352) );
  scg4d1_hd U1161 ( .A(n1011), .B(n1880), .C(n1027), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_1_), .G(n1879), .H(n1030), .Y(n1353) );
  nr2d1_hd U1162 ( .A(n1355), .B(n1354), .Y(n1385) );
  scg4d1_hd U1163 ( .A(n1027), .B(n1922), .C(n1024), .D(n1921), .E(n1919), .F(
        n1396), .G(n1920), .H(n1012), .Y(n1357) );
  xo3d1_hd U1164 ( .A(n1385), .B(n1404), .C(n1384), .Y(intadd_27_B_2_) );
  scg4d1_hd U1165 ( .A(n1034), .B(n1889), .C(n1037), .D(n1879), .E(n1888), .F(
        intadd_24_SUM_6_), .G(n1036), .H(n1880), .Y(n1358) );
  scg4d1_hd U1166 ( .A(n1041), .B(n1879), .C(n1039), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_9_), .G(n1040), .H(n1880), .Y(n1359) );
  nr2d1_hd U1167 ( .A(n1892), .B(n1378), .Y(n1360) );
  scg16d1_hd U1168 ( .A(n1381), .B(n1363), .C(n1362), .Y(intadd_28_A_0_) );
  scg4d1_hd U1169 ( .A(n1048), .B(n1934), .C(n1044), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_13_), .G(n1046), .H(n1935), .Y(n1364) );
  scg4d1_hd U1170 ( .A(n1011), .B(n1868), .C(n1027), .D(n1877), .E(n1030), .F(
        n1867), .G(n1876), .H(intadd_24_SUM_1_), .Y(n1365) );
  scg4d1_hd U1171 ( .A(n1011), .B(n1877), .C(n1031), .D(n1867), .E(n1868), .F(
        n1030), .G(n1876), .H(intadd_24_SUM_2_), .Y(n1366) );
  scg4d1_hd U1172 ( .A(n1030), .B(n1877), .C(n1031), .D(n1868), .E(n1867), .F(
        n1032), .G(n1876), .H(intadd_24_SUM_3_), .Y(n1367) );
  scg4d1_hd U1173 ( .A(n1034), .B(n1867), .C(n1031), .D(n1877), .E(n1868), .F(
        n1032), .G(n1876), .H(intadd_24_SUM_4_), .Y(n1368) );
  scg4d1_hd U1174 ( .A(n1034), .B(n1868), .C(n1036), .D(n1867), .E(n1032), .F(
        n1877), .G(n1876), .H(intadd_24_SUM_5_), .Y(n1369) );
  scg4d1_hd U1175 ( .A(n1034), .B(n1877), .C(n1037), .D(n1867), .E(n1868), .F(
        n1036), .G(n1876), .H(intadd_24_SUM_6_), .Y(n1370) );
  scg4d1_hd U1176 ( .A(n1039), .B(n1867), .C(n1037), .D(n1868), .E(n1036), .F(
        n1877), .G(n1876), .H(intadd_24_SUM_7_), .Y(n1371) );
  scg4d1_hd U1177 ( .A(n1040), .B(n1867), .C(n1037), .D(n1877), .E(n1868), .F(
        n1039), .G(n1876), .H(intadd_24_SUM_8_), .Y(n1372) );
  scg4d1_hd U1178 ( .A(n1011), .B(n1867), .C(n1012), .D(n1877), .E(n1868), .F(
        n1027), .G(n1876), .H(intadd_24_SUM_0_), .Y(n1373) );
  xo3d1_hd U1179 ( .A(n1379), .B(n1378), .C(n1377), .Y(intadd_28_B_2_) );
  scg4d1_hd U1180 ( .A(n1041), .B(n1867), .C(n1039), .D(n1877), .E(n1868), .F(
        n1040), .G(n1876), .H(intadd_24_SUM_9_), .Y(n1380) );
  nr2d1_hd U1181 ( .A(n1020), .B(n1381), .Y(n1382) );
  scg16d1_hd U1182 ( .A(n1404), .B(n1385), .C(n1384), .Y(intadd_29_A_0_) );
  scg4d1_hd U1183 ( .A(n1022), .B(n1905), .C(n1024), .D(n1904), .E(n1906), .F(
        n1012), .G(n1386), .H(n1903), .Y(n1387) );
  ao21d1_hd U1184 ( .A(n1022), .B(n1904), .C(n1389), .Y(n1406) );
  nd3d1_hd U1185 ( .A(n1060), .B(n1406), .C(n1404), .Y(n1390) );
  scg14d1_hd U1186 ( .A(n1391), .B(n1390), .C(n1909), .Y(intadd_29_A_1_) );
  scg4d1_hd U1187 ( .A(n1011), .B(n1921), .C(n1031), .D(n1922), .E(n1919), .F(
        intadd_24_SUM_2_), .G(n1030), .H(n1920), .Y(n1392) );
  scg4d1_hd U1188 ( .A(n1039), .B(n1879), .C(n1037), .D(n1880), .E(n1888), .F(
        intadd_24_SUM_7_), .G(n1889), .H(n1036), .Y(n1393) );
  scg4d1_hd U1189 ( .A(n1011), .B(n1922), .C(n1012), .D(n1921), .E(n1027), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_0_), .Y(n1394) );
  scg4d1_hd U1190 ( .A(n1011), .B(n1920), .C(n1027), .D(n1921), .E(n1922), .F(
        n1030), .G(n1919), .H(intadd_24_SUM_1_), .Y(n1395) );
  scg4d1_hd U1191 ( .A(n1027), .B(n1906), .C(n1024), .D(n1905), .E(n1012), .F(
        n1904), .G(n1903), .H(n1396), .Y(n1397) );
  xo3d1_hd U1192 ( .A(n1909), .B(n1910), .C(n1908), .Y(intadd_29_B_2_) );
  scg4d1_hd U1193 ( .A(n1030), .B(n1921), .C(n1031), .D(n1920), .E(n1922), .F(
        n1032), .G(n1919), .H(intadd_24_SUM_3_), .Y(n1398) );
  ivd1_hd U1194 ( .A(intadd_22_SUM_0_), .Y(n1853) );
  scg4d1_hd U1195 ( .A(n1011), .B(n1904), .C(n1027), .D(n1905), .E(n1906), .F(
        n1030), .G(n1903), .H(intadd_24_SUM_1_), .Y(n1399) );
  scg4d1_hd U1196 ( .A(n1034), .B(n1920), .C(n1036), .D(n1922), .E(n1919), .F(
        intadd_24_SUM_5_), .G(n1921), .H(n1032), .Y(n1400) );
  scg4d1_hd U1197 ( .A(n1034), .B(n1921), .C(n1037), .D(n1922), .E(n1919), .F(
        intadd_24_SUM_6_), .G(n1036), .H(n1920), .Y(n1401) );
  scg4d1_hd U1198 ( .A(n1043), .B(n1879), .C(n1040), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_10_), .G(n1041), .H(n1880), .Y(n1402) );
  scg4d1_hd U1199 ( .A(n1048), .B(n1868), .C(n1050), .D(n1867), .E(n1046), .F(
        n1877), .G(n1876), .H(intadd_24_SUM_14_), .Y(n1403) );
  nr2d1_hd U1200 ( .A(n1061), .B(n1404), .Y(n1405) );
  oa22d1_hd U1201 ( .A(n1059), .B(n1409), .C(n1408), .D(n1407), .Y(n1410) );
  scg4d1_hd U1202 ( .A(n1937), .B(n1930), .C(n1055), .D(n1486), .E(n1411), .F(
        n1057), .G(n1931), .H(n1053), .Y(n1412) );
  nr2d1_hd U1203 ( .A(n1061), .B(n1033), .Y(intadd_31_A_2_) );
  scg4d1_hd U1204 ( .A(n1039), .B(n1906), .C(n1037), .D(n1904), .E(n1036), .F(
        n1905), .G(n1903), .H(intadd_24_SUM_7_), .Y(n1413) );
  ao21d1_hd U1205 ( .A(a_m[8]), .B(n1415), .C(n1414), .Y(n1419) );
  scg4d1_hd U1206 ( .A(n1040), .B(n1906), .C(n1037), .D(n1905), .E(n1039), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_8_), .Y(n1416) );
  ivd1_hd U1207 ( .A(n1417), .Y(intadd_31_A_4_) );
  fad1_hd U1208 ( .A(n2039), .B(n1419), .CI(n1418), .CO(n1420), .S(n1417) );
  ivd1_hd U1209 ( .A(n1420), .Y(intadd_31_A_5_) );
  scg4d1_hd U1210 ( .A(n1034), .B(n1904), .C(n1036), .D(n1906), .E(n1032), .F(
        n1905), .G(n1903), .H(intadd_24_SUM_5_), .Y(n1421) );
  oa211d1_hd U1211 ( .A(n1035), .B(n1033), .C(a_m[23]), .D(n1523), .Y(n1422)
         );
  scg4d1_hd U1212 ( .A(n1044), .B(n1922), .C(n1041), .D(n1921), .E(n1043), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_11_), .Y(n1423) );
  scg4d1_hd U1213 ( .A(n1048), .B(n1922), .C(n1044), .D(n1921), .E(n1046), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_13_), .Y(n1424) );
  scg4d1_hd U1214 ( .A(n1055), .B(n1879), .C(n1053), .D(n1880), .E(n1888), .F(
        intadd_24_SUM_17_), .G(n1889), .H(n1051), .Y(n1425) );
  nr2d1_hd U1215 ( .A(n1061), .B(n1042), .Y(intadd_32_A_1_) );
  scg4d1_hd U1216 ( .A(n1048), .B(n1906), .C(n1044), .D(n1905), .E(n1046), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_13_), .Y(n1426) );
  nr2d1_hd U1217 ( .A(n1043), .B(n1041), .Y(n1427) );
  nr2d1_hd U1218 ( .A(n1427), .B(n1061), .Y(n1436) );
  ivd1_hd U1219 ( .A(n1436), .Y(n1428) );
  ao21d1_hd U1220 ( .A(a_m[14]), .B(n1437), .C(n1428), .Y(n1432) );
  scg4d1_hd U1221 ( .A(n1048), .B(n1904), .C(n1050), .D(n1906), .E(n1046), .F(
        n1905), .G(n1903), .H(intadd_24_SUM_14_), .Y(n1429) );
  ivd1_hd U1222 ( .A(n1430), .Y(intadd_32_A_3_) );
  fad1_hd U1223 ( .A(intadd_34_A_0_), .B(n1432), .CI(n1431), .CO(n1433), .S(
        n1430) );
  ivd1_hd U1224 ( .A(n1433), .Y(intadd_32_A_4_) );
  ivd1_hd U1225 ( .A(n2039), .Y(n1435) );
  nr2d1_hd U1226 ( .A(a_m[11]), .B(n1443), .Y(n1434) );
  oa22d1_hd U1227 ( .A(n1039), .B(n1939), .C(n1435), .D(n1434), .Y(
        intadd_32_B_0_) );
  scg4d1_hd U1228 ( .A(n1055), .B(n1922), .C(n1053), .D(n1920), .E(n1051), .F(
        n1921), .G(n1919), .H(intadd_24_SUM_17_), .Y(n1439) );
  scg4d1_hd U1229 ( .A(n1057), .B(n1920), .C(b_m[23]), .D(n1922), .E(n1919), 
        .F(n1460), .G(n1921), .H(n1055), .Y(n1440) );
  scg4d1_hd U1230 ( .A(n1044), .B(n1906), .C(n1041), .D(n1905), .E(n1043), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_11_), .Y(n1441) );
  scg4d1_hd U1231 ( .A(n1043), .B(n1906), .C(n1040), .D(n1905), .E(n1041), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_10_), .Y(n1442) );
  nr2d1_hd U1232 ( .A(n1061), .B(n1038), .Y(intadd_33_B_0_) );
  oa22d1_hd U1233 ( .A(n1036), .B(n1443), .C(n1039), .D(n2039), .Y(n1444) );
  scg4d1_hd U1234 ( .A(n1048), .B(n1920), .C(n1050), .D(n1922), .E(n1919), .F(
        intadd_24_SUM_14_), .G(n1921), .H(n1046), .Y(n1445) );
  scg4d1_hd U1235 ( .A(n1057), .B(n1880), .C(b_m[23]), .D(n1879), .E(n1888), 
        .F(n1460), .G(n1889), .H(n1055), .Y(n1446) );
  scg4d1_hd U1236 ( .A(n1041), .B(n1906), .C(n1039), .D(n1905), .E(n1040), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_9_), .Y(n1447) );
  scg4d1_hd U1237 ( .A(n1051), .B(n1904), .C(n1050), .D(n1905), .E(n1906), .F(
        n1053), .G(n1903), .H(intadd_24_SUM_16_), .Y(n1448) );
  nr2d1_hd U1238 ( .A(n1061), .B(n1047), .Y(intadd_34_B_0_) );
  oa211d1_hd U1239 ( .A(n1049), .B(n1045), .C(n1060), .D(n1531), .Y(n1449) );
  ao22d1_hd U1240 ( .A(b_m[23]), .B(n1920), .C(n1919), .D(n1857), .Y(n1450) );
  oa21d1_hd U1241 ( .A(n1058), .B(n1451), .C(n1450), .Y(n1452) );
  scg4d1_hd U1242 ( .A(n1048), .B(n1905), .C(n1050), .D(n1904), .E(n1906), .F(
        n1051), .G(n1903), .H(intadd_24_SUM_15_), .Y(n1453) );
  scg4d1_hd U1243 ( .A(n1034), .B(n1906), .C(n1031), .D(n1905), .E(n1032), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_4_), .Y(n1454) );
  nr2d1_hd U1244 ( .A(n1061), .B(n1029), .Y(intadd_35_B_0_) );
  scg4d1_hd U1245 ( .A(n1040), .B(n1922), .C(n1037), .D(n1921), .E(n1039), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_8_), .Y(n1455) );
  scg4d1_hd U1246 ( .A(n1030), .B(n1905), .C(n1031), .D(n1904), .E(n1906), .F(
        n1032), .G(n1903), .H(intadd_24_SUM_3_), .Y(n1456) );
  nr2d1_hd U1247 ( .A(n1061), .B(n1052), .Y(intadd_36_A_1_) );
  oa211d1_hd U1248 ( .A(n1052), .B(n1054), .C(n1060), .D(n1855), .Y(n1457) );
  ivd1_hd U1249 ( .A(intadd_34_A_0_), .Y(n1459) );
  nr3d1_hd U1250 ( .A(a_m[17]), .B(n1061), .C(n1049), .Y(n1458) );
  oa22d1_hd U1251 ( .A(n1048), .B(n1020), .C(n1459), .D(n1458), .Y(
        intadd_36_B_0_) );
  scg4d1_hd U1252 ( .A(n1057), .B(n1904), .C(b_m[23]), .D(n1906), .E(n1055), 
        .F(n1905), .G(n1903), .H(n1460), .Y(n1461) );
  scg4d1_hd U1253 ( .A(n1046), .B(n1906), .C(n1043), .D(n1905), .E(n1044), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_12_), .Y(n1463) );
  scg4d1_hd U1254 ( .A(n1048), .B(n1921), .C(n1050), .D(n1920), .E(n1922), .F(
        n1051), .G(n1919), .H(intadd_24_SUM_15_), .Y(n1464) );
  scg4d1_hd U1255 ( .A(n1051), .B(n1920), .C(n1050), .D(n1921), .E(n1922), .F(
        n1053), .G(n1919), .H(intadd_24_SUM_16_), .Y(n1465) );
  ao22d1_hd U1256 ( .A(b_m[23]), .B(n1880), .C(n1888), .D(n1857), .Y(n1466) );
  scg14d1_hd U1257 ( .A(n1889), .B(n1057), .C(n1466), .Y(n1467) );
  scg4d1_hd U1258 ( .A(n1046), .B(n1922), .C(n1043), .D(n1921), .E(n1044), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_12_), .Y(n1468) );
  scg4d1_hd U1259 ( .A(n1051), .B(n1880), .C(n1050), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_16_), .G(n1879), .H(n1053), .Y(n1469) );
  ao22d1_hd U1260 ( .A(b_m[23]), .B(n1868), .C(n1876), .D(n1857), .Y(n1470) );
  oa21d1_hd U1261 ( .A(n1471), .B(n1058), .C(n1470), .Y(n1472) );
  scg4d1_hd U1262 ( .A(n1048), .B(n1889), .C(n1050), .D(n1880), .E(n1888), .F(
        intadd_24_SUM_15_), .G(n1051), .H(n1879), .Y(n1473) );
  scg4d1_hd U1263 ( .A(n1046), .B(n1879), .C(n1043), .D(n1889), .E(n1888), .F(
        intadd_24_SUM_12_), .G(n1044), .H(n1880), .Y(n1474) );
  scg4d1_hd U1264 ( .A(n1051), .B(n1868), .C(n1050), .D(n1877), .E(n1053), .F(
        n1867), .G(n1876), .H(intadd_24_SUM_16_), .Y(n1475) );
  ao22d1_hd U1265 ( .A(n1057), .B(n1009), .C(n1936), .D(n1857), .Y(n1476) );
  oa21d1_hd U1266 ( .A(n1059), .B(n1477), .C(n1476), .Y(n1478) );
  scg4d1_hd U1267 ( .A(n1048), .B(n1877), .C(n1050), .D(n1868), .E(n1867), .F(
        n1051), .G(n1876), .H(intadd_24_SUM_15_), .Y(n1479) );
  scg4d1_hd U1268 ( .A(n1034), .B(n1905), .C(n1037), .D(n1906), .E(n1904), .F(
        n1036), .G(n1903), .H(intadd_24_SUM_6_), .Y(n1480) );
  scg4d1_hd U1269 ( .A(n1043), .B(n1922), .C(n1040), .D(n1921), .E(n1041), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_10_), .Y(n1481) );
  scg4d1_hd U1270 ( .A(n1048), .B(n1880), .C(n1050), .D(n1879), .E(n1888), .F(
        intadd_24_SUM_14_), .G(n1889), .H(n1046), .Y(n1482) );
  scg4d1_hd U1271 ( .A(n1041), .B(n1922), .C(n1039), .D(n1921), .E(n1040), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_9_), .Y(n1483) );
  scg4d1_hd U1272 ( .A(n1046), .B(n1867), .C(n1043), .D(n1877), .E(n1868), .F(
        n1044), .G(n1876), .H(intadd_24_SUM_12_), .Y(n1484) );
  scg4d1_hd U1273 ( .A(n1051), .B(n1935), .C(n1050), .D(n1009), .E(n1936), .F(
        intadd_24_SUM_16_), .G(n1934), .H(n1053), .Y(n1485) );
  ao22d1_hd U1274 ( .A(b_m[23]), .B(n1486), .C(n1930), .D(n1857), .Y(n1487) );
  oa21d1_hd U1275 ( .A(n1488), .B(n1058), .C(n1487), .Y(n1489) );
  scg4d1_hd U1276 ( .A(n1048), .B(n1009), .C(n1050), .D(n1935), .E(n1936), .F(
        intadd_24_SUM_15_), .G(n1934), .H(n1051), .Y(n1490) );
  ao22d1_hd U1277 ( .A(n1113), .B(DP_OP_125J3_130_6300_n34), .C(z_e[0]), .D(
        n1844), .Y(n1004) );
  oa22ad1_hd U1278 ( .A(n1818), .B(n1496), .C(n1112), .D(round_bit), .Y(n1491)
         );
  ao21d1_hd U1279 ( .A(n1710), .B(product[25]), .C(n1491), .Y(n104) );
  nr2d1_hd U1280 ( .A(z_e[4]), .B(z_e[3]), .Y(n1493) );
  nr2d1_hd U1281 ( .A(z_e[6]), .B(z_e[5]), .Y(n1492) );
  nr3d1_hd U1282 ( .A(z_e[2]), .B(z_e[1]), .C(n1555), .Y(n1494) );
  oa21d1_hd U1283 ( .A(n1494), .B(n1554), .C(z_e[9]), .Y(n1807) );
  nr2d1_hd U1284 ( .A(n1807), .B(n1818), .Y(n1697) );
  ao21d1_hd U1285 ( .A(n1112), .B(n1814), .C(n1697), .Y(n1499) );
  nd3d1_hd U1286 ( .A(z_m[0]), .B(z_m[1]), .C(z_m[2]), .Y(n1674) );
  ivd1_hd U1287 ( .A(n1674), .Y(n1673) );
  nd3d1_hd U1288 ( .A(n1673), .B(z_m[3]), .C(z_m[4]), .Y(n1665) );
  ivd1_hd U1289 ( .A(n1665), .Y(n1664) );
  nd3d1_hd U1290 ( .A(n1664), .B(z_m[5]), .C(z_m[6]), .Y(n1656) );
  ivd1_hd U1291 ( .A(n1656), .Y(n1655) );
  nd3d1_hd U1292 ( .A(n1655), .B(z_m[7]), .C(z_m[8]), .Y(n1647) );
  ivd1_hd U1293 ( .A(n1647), .Y(n1646) );
  nd3d1_hd U1294 ( .A(n1646), .B(z_m[9]), .C(z_m[10]), .Y(n1638) );
  nd3d1_hd U1295 ( .A(n1637), .B(z_m[11]), .C(z_m[12]), .Y(n1629) );
  nd3d1_hd U1296 ( .A(n1628), .B(z_m[13]), .C(z_m[14]), .Y(n1620) );
  nd3d1_hd U1297 ( .A(n1619), .B(z_m[15]), .C(z_m[16]), .Y(n1611) );
  nd3d1_hd U1298 ( .A(n1609), .B(z_m[17]), .C(z_m[18]), .Y(n1601) );
  nd3d1_hd U1299 ( .A(n1600), .B(z_m[19]), .C(z_m[20]), .Y(n1594) );
  ivd1_hd U1300 ( .A(n1594), .Y(n1592) );
  nd3d1_hd U1301 ( .A(z_m[22]), .B(z_m[21]), .C(n1592), .Y(n1717) );
  nr2d1_hd U1302 ( .A(round_bit), .B(sticky), .Y(n1497) );
  ao211d1_hd U1303 ( .A(n1497), .B(n1496), .C(net922), .D(n1610), .Y(n1591) );
  nr4d1_hd U1304 ( .A(a_e[4]), .B(n10), .C(a_e[6]), .D(a_e[1]), .Y(n1501) );
  scg13d1_hd U1305 ( .A(a_e[3]), .B(a_e[2]), .C(n1501), .Y(n1504) );
  ivd1_hd U1306 ( .A(a_e[5]), .Y(n1502) );
  nd4d1_hd U1307 ( .A(a_e[9]), .B(a_e[8]), .C(a_e[0]), .D(n1502), .Y(n1503) );
  nd2bd1_hd U1308 ( .AN(n1504), .B(n1758), .Y(n1505) );
  nr4d1_hd U1309 ( .A(a_e[8]), .B(a_e[5]), .C(a_e[0]), .D(n1505), .Y(n1542) );
  nr4d1_hd U1310 ( .A(b_e[5]), .B(b_e[2]), .C(b_e[1]), .D(n14), .Y(n1507) );
  nr2d1_hd U1311 ( .A(b_e[6]), .B(b_e[3]), .Y(n1506) );
  nr4d1_hd U1312 ( .A(b_e[4]), .B(b_e[0]), .C(n1521), .D(n1508), .Y(n1540) );
  nr2d1_hd U1313 ( .A(n1542), .B(n1540), .Y(n1550) );
  nd4d1_hd U1314 ( .A(n1779), .B(n1939), .C(n1781), .D(n1775), .Y(n1520) );
  nd4d1_hd U1315 ( .A(n1020), .B(n1771), .C(n1773), .D(n1787), .Y(n1519) );
  nd4d1_hd U1316 ( .A(n1512), .B(n1511), .C(n1510), .D(n1509), .Y(n1518) );
  nd4d1_hd U1317 ( .A(n1516), .B(n1515), .C(n1514), .D(n1513), .Y(n1517) );
  nr4d1_hd U1318 ( .A(n1520), .B(n1519), .C(n1518), .D(n1517), .Y(n1536) );
  nr4d1_hd U1319 ( .A(n1057), .B(n1030), .C(n1027), .D(n1022), .Y(n1529) );
  nr4d1_hd U1320 ( .A(n1525), .B(n1855), .C(n1524), .D(n1523), .Y(n1528) );
  nr4d1_hd U1321 ( .A(n1031), .B(n1039), .C(n1036), .D(n1037), .Y(n1527) );
  nr4d1_hd U1322 ( .A(n1043), .B(n1041), .C(n1050), .D(n1040), .Y(n1526) );
  nd4d1_hd U1323 ( .A(n1529), .B(n1528), .C(n1527), .D(n1526), .Y(n1530) );
  nr4d1_hd U1324 ( .A(n1046), .B(n1011), .C(n1531), .D(n1530), .Y(n1538) );
  ivd1_hd U1325 ( .A(n1744), .Y(n1746) );
  ivd1_hd U1326 ( .A(DP_OP_113J3_124_6892_n3), .Y(n1745) );
  ao22d1_hd U1327 ( .A(DP_OP_113J3_124_6892_n3), .B(n1744), .C(n1746), .D(
        n1745), .Y(n1532) );
  ao22d1_hd U1328 ( .A(n1749), .B(a_e[7]), .C(n1754), .D(n1532), .Y(n141) );
  oa22ad1_hd U1329 ( .A(n1762), .B(n14), .C(n1120), .D(b[30]), .Y(n1534) );
  nr2d1_hd U1330 ( .A(DP_OP_116J3_127_7148_n3), .B(n1534), .Y(n1761) );
  oa22ad1_hd U1331 ( .A(n14), .B(n1843), .C(n1838), .D(n1761), .Y(n1533) );
  ao21d1_hd U1332 ( .A(DP_OP_116J3_127_7148_n3), .B(n1534), .C(n1533), .Y(n151) );
  ao22d1_hd U1333 ( .A(n1542), .B(n1541), .C(n1540), .D(n1539), .Y(n1544) );
  nr2d1_hd U1334 ( .A(n1544), .B(n1543), .Y(n1589) );
  ao22d1_hd U1335 ( .A(n1552), .B(N35), .C(n1551), .D(z_s), .Y(n1548) );
  ivd1_hd U1336 ( .A(n1550), .Y(n1553) );
  nr2d1_hd U1337 ( .A(z_e[1]), .B(z_e[0]), .Y(n1580) );
  ivd1_hd U1338 ( .A(z_e[2]), .Y(n1576) );
  nr2d1_hd U1339 ( .A(z_e[3]), .B(n1575), .Y(n1572) );
  ivd1_hd U1340 ( .A(z_e[4]), .Y(n1569) );
  nr2d1_hd U1341 ( .A(z_e[5]), .B(n1568), .Y(n1565) );
  ivd1_hd U1342 ( .A(z_e[6]), .Y(n1562) );
  nr2d1_hd U1343 ( .A(z_m[23]), .B(z_e[0]), .Y(n1558) );
  ivd1_hd U1344 ( .A(z_e[1]), .Y(n1556) );
  nr4d1_hd U1345 ( .A(z_e[2]), .B(n1556), .C(n1555), .D(n1554), .Y(n1557) );
  oa211d1_hd U1346 ( .A(z_e[7]), .B(n1561), .C(n1578), .D(n1559), .Y(n1560) );
  scg15d1_hd U1347 ( .A(n1016), .B(z[30]), .C(n1584), .D(n1560), .Y(n230) );
  oa21d1_hd U1348 ( .A(n1565), .B(n1562), .C(n1561), .Y(n1563) );
  ao22d1_hd U1349 ( .A(n1016), .B(z[29]), .C(n1578), .D(n1563), .Y(n1564) );
  ao21d1_hd U1350 ( .A(z_e[5]), .B(n1568), .C(n1565), .Y(n1567) );
  oa211d1_hd U1351 ( .A(n1567), .B(n1585), .C(n1584), .D(n1566), .Y(n232) );
  oa21d1_hd U1352 ( .A(n1572), .B(n1569), .C(n1568), .Y(n1570) );
  ao22d1_hd U1353 ( .A(n1016), .B(z[27]), .C(n1578), .D(n1570), .Y(n1571) );
  ao21d1_hd U1354 ( .A(z_e[3]), .B(n1575), .C(n1572), .Y(n1574) );
  oa211d1_hd U1355 ( .A(n1574), .B(n1585), .C(n1584), .D(n1573), .Y(n234) );
  oa21d1_hd U1356 ( .A(n1580), .B(n1576), .C(n1575), .Y(n1577) );
  ao22d1_hd U1357 ( .A(n1016), .B(z[25]), .C(n1578), .D(n1577), .Y(n1579) );
  ao21d1_hd U1358 ( .A(z_e[0]), .B(z_e[1]), .C(n1580), .Y(n1582) );
  oa211d1_hd U1359 ( .A(n1582), .B(n1585), .C(n1584), .D(n1581), .Y(n236) );
  oa211d1_hd U1360 ( .A(z_e[0]), .B(n1585), .C(n1584), .D(n1583), .Y(n237) );
  scg17d1_hd U1361 ( .A(z_m[22]), .B(n1590), .C(n1589), .D(n1588), .Y(n238) );
  ao21d1_hd U1362 ( .A(n1709), .B(n1594), .C(n1705), .Y(n1597) );
  ivd1_hd U1363 ( .A(z_m[21]), .Y(n1596) );
  nr2d1_hd U1364 ( .A(z_m[22]), .B(n1684), .Y(n1713) );
  scg6d1_hd U1365 ( .A(n1592), .B(n1713), .C(n1711), .Y(n1593) );
  scg4d1_hd U1366 ( .A(n1712), .B(z_m[22]), .C(n1593), .D(z_m[21]), .E(n1710), 
        .F(product[48]), .G(z_m[23]), .H(n1703), .Y(n261) );
  oa22d1_hd U1367 ( .A(n1597), .B(n1596), .C(n1595), .D(n1594), .Y(n1599) );
  ao22d1_hd U1368 ( .A(z_m[22]), .B(n1017), .C(n1710), .D(product[47]), .Y(
        n1598) );
  oa21d1_hd U1369 ( .A(z_m[20]), .B(n1605), .C(n1708), .Y(n1603) );
  ao21d1_hd U1370 ( .A(n1701), .B(n1601), .C(n1705), .Y(n1606) );
  oa21d1_hd U1371 ( .A(z_m[19]), .B(n1684), .C(n1606), .Y(n1602) );
  scg4d1_hd U1372 ( .A(n1603), .B(z_m[19]), .C(n1602), .D(z_m[20]), .E(z_m[21]), .F(n1017), .G(n1710), .H(product[46]), .Y(n263) );
  ivd1_hd U1373 ( .A(z_m[19]), .Y(n1604) );
  ao22d1_hd U1374 ( .A(z_m[19]), .B(n1606), .C(n1605), .D(n1604), .Y(n1608) );
  ao22d1_hd U1375 ( .A(n1710), .B(product[45]), .C(z_m[20]), .D(n1017), .Y(
        n1607) );
  oa21d1_hd U1376 ( .A(z_m[18]), .B(n1618), .C(n1708), .Y(n1613) );
  ivd1_hd U1377 ( .A(n1610), .Y(n1675) );
  ao21d1_hd U1378 ( .A(n1675), .B(n1611), .C(n1705), .Y(n1614) );
  oa21d1_hd U1379 ( .A(z_m[17]), .B(n1684), .C(n1614), .Y(n1612) );
  scg4d1_hd U1380 ( .A(n1613), .B(z_m[17]), .C(n1612), .D(z_m[18]), .E(z_m[19]), .F(n1017), .G(n1710), .H(product[44]), .Y(n265) );
  ao22d1_hd U1381 ( .A(n1710), .B(product[43]), .C(z_m[18]), .D(n1703), .Y(
        n1617) );
  ivd1_hd U1382 ( .A(n1614), .Y(n1615) );
  ao22d1_hd U1383 ( .A(z_m[16]), .B(n1711), .C(z_m[17]), .D(n1615), .Y(n1616)
         );
  oa211d1_hd U1384 ( .A(z_m[17]), .B(n1618), .C(n1617), .D(n1616), .Y(n266) );
  oa21d1_hd U1385 ( .A(z_m[16]), .B(n1624), .C(n1708), .Y(n1622) );
  ao21d1_hd U1386 ( .A(n1701), .B(n1620), .C(n1705), .Y(n1625) );
  oa21d1_hd U1387 ( .A(z_m[15]), .B(n1684), .C(n1625), .Y(n1621) );
  scg4d1_hd U1388 ( .A(n1622), .B(z_m[15]), .C(n1621), .D(z_m[16]), .E(z_m[17]), .F(n1017), .G(n1710), .H(product[42]), .Y(n267) );
  ivd1_hd U1389 ( .A(z_m[15]), .Y(n1623) );
  ao22d1_hd U1390 ( .A(z_m[15]), .B(n1625), .C(n1624), .D(n1623), .Y(n1627) );
  ao22d1_hd U1391 ( .A(n1710), .B(product[41]), .C(z_m[16]), .D(n1703), .Y(
        n1626) );
  oa21d1_hd U1392 ( .A(z_m[14]), .B(n1636), .C(n1708), .Y(n1631) );
  ao21d1_hd U1393 ( .A(n1675), .B(n1629), .C(n1705), .Y(n1632) );
  oa21d1_hd U1394 ( .A(z_m[13]), .B(n1684), .C(n1632), .Y(n1630) );
  scg4d1_hd U1395 ( .A(n1631), .B(z_m[13]), .C(n1630), .D(z_m[14]), .E(z_m[15]), .F(n1017), .G(n1710), .H(product[40]), .Y(n269) );
  ao22d1_hd U1396 ( .A(n1710), .B(product[39]), .C(z_m[14]), .D(n1703), .Y(
        n1635) );
  ivd1_hd U1397 ( .A(n1632), .Y(n1633) );
  ao22d1_hd U1398 ( .A(z_m[12]), .B(n1711), .C(z_m[13]), .D(n1633), .Y(n1634)
         );
  oa211d1_hd U1399 ( .A(z_m[13]), .B(n1636), .C(n1635), .D(n1634), .Y(n270) );
  oa21d1_hd U1400 ( .A(z_m[12]), .B(n1642), .C(n1708), .Y(n1640) );
  ao21d1_hd U1401 ( .A(n1675), .B(n1638), .C(n1705), .Y(n1643) );
  oa21d1_hd U1402 ( .A(z_m[11]), .B(n1684), .C(n1643), .Y(n1639) );
  scg4d1_hd U1403 ( .A(n1640), .B(z_m[11]), .C(n1639), .D(z_m[12]), .E(z_m[13]), .F(n1017), .G(n1710), .H(product[38]), .Y(n271) );
  ivd1_hd U1404 ( .A(z_m[11]), .Y(n1641) );
  ao22d1_hd U1405 ( .A(z_m[11]), .B(n1643), .C(n1642), .D(n1641), .Y(n1645) );
  ao22d1_hd U1406 ( .A(n1710), .B(product[37]), .C(z_m[12]), .D(n1017), .Y(
        n1644) );
  oa21d1_hd U1407 ( .A(z_m[10]), .B(n1654), .C(n1708), .Y(n1649) );
  ao21d1_hd U1408 ( .A(n1701), .B(n1647), .C(n1705), .Y(n1650) );
  oa21d1_hd U1409 ( .A(z_m[9]), .B(n1684), .C(n1650), .Y(n1648) );
  scg4d1_hd U1410 ( .A(n1649), .B(z_m[9]), .C(n1648), .D(z_m[10]), .E(z_m[11]), 
        .F(n1017), .G(n1710), .H(product[36]), .Y(n273) );
  ao22d1_hd U1411 ( .A(n1710), .B(product[35]), .C(z_m[10]), .D(n1017), .Y(
        n1653) );
  ivd1_hd U1412 ( .A(n1650), .Y(n1651) );
  ao22d1_hd U1413 ( .A(z_m[8]), .B(n1711), .C(z_m[9]), .D(n1651), .Y(n1652) );
  oa211d1_hd U1414 ( .A(z_m[9]), .B(n1654), .C(n1653), .D(n1652), .Y(n274) );
  oa21d1_hd U1415 ( .A(z_m[8]), .B(n1660), .C(n1708), .Y(n1658) );
  ao21d1_hd U1416 ( .A(n1675), .B(n1656), .C(n1705), .Y(n1661) );
  oa21d1_hd U1417 ( .A(z_m[7]), .B(n1684), .C(n1661), .Y(n1657) );
  scg4d1_hd U1418 ( .A(n1658), .B(z_m[7]), .C(n1657), .D(z_m[8]), .E(z_m[9]), 
        .F(n1017), .G(n1710), .H(product[34]), .Y(n275) );
  ivd1_hd U1419 ( .A(z_m[7]), .Y(n1659) );
  ao22d1_hd U1420 ( .A(z_m[7]), .B(n1661), .C(n1660), .D(n1659), .Y(n1663) );
  ao22d1_hd U1421 ( .A(n1710), .B(product[33]), .C(z_m[8]), .D(n1703), .Y(
        n1662) );
  oa21d1_hd U1422 ( .A(z_m[6]), .B(n1672), .C(n1708), .Y(n1667) );
  ao21d1_hd U1423 ( .A(n1701), .B(n1665), .C(n1705), .Y(n1668) );
  oa21d1_hd U1424 ( .A(z_m[5]), .B(n1684), .C(n1668), .Y(n1666) );
  scg4d1_hd U1425 ( .A(n1667), .B(z_m[5]), .C(n1666), .D(z_m[6]), .E(z_m[7]), 
        .F(n1017), .G(n1710), .H(product[32]), .Y(n277) );
  ao22d1_hd U1426 ( .A(n1710), .B(product[31]), .C(z_m[6]), .D(n1703), .Y(
        n1671) );
  ivd1_hd U1427 ( .A(n1668), .Y(n1669) );
  ao22d1_hd U1428 ( .A(z_m[4]), .B(n1711), .C(z_m[5]), .D(n1669), .Y(n1670) );
  oa211d1_hd U1429 ( .A(z_m[5]), .B(n1672), .C(n1671), .D(n1670), .Y(n278) );
  oa21d1_hd U1430 ( .A(z_m[4]), .B(n1679), .C(n1708), .Y(n1677) );
  ao21d1_hd U1431 ( .A(n1675), .B(n1674), .C(n1705), .Y(n1680) );
  oa21d1_hd U1432 ( .A(z_m[3]), .B(n1684), .C(n1680), .Y(n1676) );
  scg4d1_hd U1433 ( .A(n1677), .B(z_m[3]), .C(n1676), .D(z_m[4]), .E(z_m[5]), 
        .F(n1017), .G(n1710), .H(product[30]), .Y(n279) );
  ivd1_hd U1434 ( .A(z_m[3]), .Y(n1678) );
  ao22d1_hd U1435 ( .A(z_m[3]), .B(n1680), .C(n1679), .D(n1678), .Y(n1682) );
  ao22d1_hd U1436 ( .A(n1710), .B(product[29]), .C(z_m[4]), .D(n1017), .Y(
        n1681) );
  oa21d1_hd U1437 ( .A(z_m[2]), .B(n1683), .C(n1708), .Y(n1686) );
  nr2d1_hd U1438 ( .A(z_m[0]), .B(n1684), .Y(n1704) );
  nr2d1_hd U1439 ( .A(n1705), .B(n1704), .Y(n1688) );
  nd2bd1_hd U1440 ( .AN(z_m[1]), .B(n1709), .Y(n1687) );
  scg4d1_hd U1441 ( .A(n1686), .B(z_m[1]), .C(n1685), .D(z_m[2]), .E(z_m[3]), 
        .F(n1017), .G(n1710), .H(product[28]), .Y(n281) );
  ivd1_hd U1442 ( .A(n1688), .Y(n1689) );
  scg4d1_hd U1443 ( .A(n1690), .B(z_m[0]), .C(n1689), .D(z_m[1]), .E(z_m[2]), 
        .F(n1017), .G(n1710), .H(product[27]), .Y(n282) );
  nr4d1_hd U1444 ( .A(product[14]), .B(product[12]), .C(product[19]), .D(
        product[17]), .Y(n1694) );
  nr4d1_hd U1445 ( .A(product[15]), .B(product[8]), .C(product[20]), .D(
        product[4]), .Y(n1693) );
  nr4d1_hd U1446 ( .A(product[21]), .B(product[2]), .C(product[13]), .D(
        product[16]), .Y(n1692) );
  nr4d1_hd U1447 ( .A(product[23]), .B(product[5]), .C(product[22]), .D(
        product[18]), .Y(n1691) );
  nd4d1_hd U1448 ( .A(n1694), .B(n1693), .C(n1692), .D(n1691), .Y(n1695) );
  nr4d1_hd U1449 ( .A(product[9]), .B(product[7]), .C(n1696), .D(n1695), .Y(
        n1700) );
  ao22d1_hd U1450 ( .A(round_bit), .B(n1697), .C(sticky), .D(n1699), .Y(n1698)
         );
  oa21d1_hd U1451 ( .A(n1700), .B(n1699), .C(n1698), .Y(n283) );
  ao22d1_hd U1452 ( .A(n1710), .B(product[24]), .C(n1701), .D(round_bit), .Y(
        n1702) );
  scg16d1_hd U1453 ( .A(n1017), .B(net922), .C(n1702), .Y(n284) );
  ao22d1_hd U1454 ( .A(n1710), .B(product[26]), .C(z_m[1]), .D(n1703), .Y(
        n1707) );
  ao21d1_hd U1455 ( .A(n1705), .B(z_m[0]), .C(n1704), .Y(n1706) );
  oa211d1_hd U1456 ( .A(net922), .B(n1708), .C(n1707), .D(n1706), .Y(n285) );
  ao22d1_hd U1457 ( .A(z_m[22]), .B(n1711), .C(n1710), .D(product[49]), .Y(
        n1715) );
  oa21d1_hd U1458 ( .A(n1713), .B(n1712), .C(z_m[23]), .Y(n1714) );
  oa211d1_hd U1459 ( .A(n1717), .B(n1716), .C(n1715), .D(n1714), .Y(n286) );
  ao22d1_hd U1460 ( .A(n1120), .B(b[22]), .C(n1057), .D(n1018), .Y(n1718) );
  oa21d1_hd U1461 ( .A(n1056), .B(n1740), .C(n1718), .Y(n287) );
  ao22d1_hd U1462 ( .A(n1120), .B(b[20]), .C(n1053), .D(n1018), .Y(n1719) );
  oa21d1_hd U1463 ( .A(n1052), .B(n1740), .C(n1719), .Y(n288) );
  ao22d1_hd U1464 ( .A(n1120), .B(b[19]), .C(n1051), .D(n1018), .Y(n1720) );
  scg16d1_hd U1465 ( .A(n1050), .B(n1740), .C(n1720), .Y(n289) );
  ao22d1_hd U1466 ( .A(n1120), .B(b[18]), .C(n1050), .D(n1018), .Y(n1721) );
  oa21d1_hd U1467 ( .A(n1049), .B(n1740), .C(n1721), .Y(n290) );
  ao22d1_hd U1468 ( .A(n1120), .B(b[17]), .C(n1048), .D(n1018), .Y(n1722) );
  oa21d1_hd U1469 ( .A(n1047), .B(n1740), .C(n1722), .Y(n291) );
  ao22d1_hd U1470 ( .A(n1120), .B(b[16]), .C(n1046), .D(n1018), .Y(n1723) );
  oa21d1_hd U1471 ( .A(n1045), .B(n1740), .C(n1723), .Y(n292) );
  ao22d1_hd U1472 ( .A(n1120), .B(b[15]), .C(n1044), .D(n1018), .Y(n1724) );
  scg16d1_hd U1473 ( .A(n1043), .B(n1740), .C(n1724), .Y(n293) );
  ao22d1_hd U1474 ( .A(n1120), .B(b[14]), .C(n1043), .D(n1018), .Y(n1725) );
  oa21d1_hd U1475 ( .A(n1042), .B(n1740), .C(n1725), .Y(n294) );
  ao22d1_hd U1476 ( .A(n1120), .B(b[13]), .C(n1041), .D(n1018), .Y(n1726) );
  scg16d1_hd U1477 ( .A(n1040), .B(n1740), .C(n1726), .Y(n295) );
  ao22d1_hd U1478 ( .A(n1120), .B(b[12]), .C(n1040), .D(n1018), .Y(n1727) );
  scg16d1_hd U1479 ( .A(n1039), .B(n1740), .C(n1727), .Y(n296) );
  ao22d1_hd U1480 ( .A(n1120), .B(b[11]), .C(n1039), .D(n1018), .Y(n1728) );
  oa21d1_hd U1481 ( .A(n1038), .B(n1740), .C(n1728), .Y(n297) );
  ao22d1_hd U1482 ( .A(n1120), .B(b[10]), .C(n1037), .D(n1018), .Y(n1729) );
  scg16d1_hd U1483 ( .A(n1036), .B(n1740), .C(n1729), .Y(n298) );
  ao22d1_hd U1484 ( .A(n1120), .B(b[9]), .C(n1036), .D(n1018), .Y(n1730) );
  oa21d1_hd U1485 ( .A(n1035), .B(n1740), .C(n1730), .Y(n299) );
  ao22d1_hd U1486 ( .A(n1120), .B(b[8]), .C(n1034), .D(n1018), .Y(n1731) );
  oa21d1_hd U1487 ( .A(n1033), .B(n1740), .C(n1731), .Y(n300) );
  ao22d1_hd U1488 ( .A(n1120), .B(b[7]), .C(n1032), .D(n1018), .Y(n1732) );
  scg16d1_hd U1489 ( .A(n1031), .B(n1740), .C(n1732), .Y(n301) );
  ao22d1_hd U1490 ( .A(n1120), .B(b[6]), .C(n1031), .D(n1018), .Y(n1733) );
  scg16d1_hd U1491 ( .A(n1030), .B(n1740), .C(n1733), .Y(n302) );
  ao22d1_hd U1492 ( .A(n1120), .B(b[5]), .C(n1030), .D(n1018), .Y(n1734) );
  oa21d1_hd U1493 ( .A(n1029), .B(n1740), .C(n1734), .Y(n303) );
  ao22d1_hd U1494 ( .A(n1120), .B(b[4]), .C(n1011), .D(n1018), .Y(n1735) );
  oa21d1_hd U1495 ( .A(n1028), .B(n1740), .C(n1735), .Y(n304) );
  ao22d1_hd U1496 ( .A(n1120), .B(b[3]), .C(n1027), .D(n1018), .Y(n1736) );
  oa21d1_hd U1497 ( .A(n1026), .B(n1740), .C(n1736), .Y(n305) );
  ao22d1_hd U1498 ( .A(n1120), .B(b[2]), .C(n1012), .D(n1018), .Y(n1737) );
  oa21d1_hd U1499 ( .A(n1025), .B(n1740), .C(n1737), .Y(n306) );
  ao22d1_hd U1500 ( .A(n1120), .B(b[1]), .C(n1024), .D(n1018), .Y(n1738) );
  oa21d1_hd U1501 ( .A(n1014), .B(n1740), .C(n1738), .Y(n307) );
  ao22d1_hd U1502 ( .A(n1120), .B(b[21]), .C(n1055), .D(n1018), .Y(n1739) );
  oa21d1_hd U1503 ( .A(n1054), .B(n1740), .C(n1739), .Y(n309) );
  ao22d1_hd U1504 ( .A(n1850), .B(n1057), .C(b_m[23]), .D(n1007), .Y(n1742) );
  oa21d1_hd U1505 ( .A(n1743), .B(n1835), .C(n1742), .Y(n310) );
  oa211d1_hd U1506 ( .A(n1808), .B(n1745), .C(n1759), .D(n1744), .Y(n1747) );
  ao211d1_hd U1507 ( .A(a_e[8]), .B(n1833), .C(DP_OP_113J3_124_6892_n3), .D(
        n1746), .Y(n1756) );
  ao22d1_hd U1508 ( .A(a_e[8]), .B(n1747), .C(n1756), .D(n1754), .Y(n1748) );
  ao22d1_hd U1509 ( .A(a_e[1]), .B(n1749), .C(C81_DATA2_1), .D(n1754), .Y(
        n1750) );
  ivd1_hd U1510 ( .A(a_e[0]), .Y(n1751) );
  nr2d1_hd U1511 ( .A(n1808), .B(n1751), .Y(n768) );
  ivd1_hd U1512 ( .A(n1754), .Y(n1752) );
  oa22d1_hd U1513 ( .A(n1752), .B(n768), .C(n1751), .D(n1759), .Y(n318) );
  nr2d1_hd U1514 ( .A(n1808), .B(n1758), .Y(n1755) );
  oa211d1_hd U1515 ( .A(n1756), .B(n1755), .C(n1754), .D(n1753), .Y(n1757) );
  oa211d1_hd U1516 ( .A(n1759), .B(n1758), .C(n138), .D(n1757), .Y(n319) );
  oa21d1_hd U1517 ( .A(n1760), .B(n1762), .C(n1761), .Y(n1840) );
  oa21d1_hd U1518 ( .A(n1762), .B(n1761), .C(n1843), .Y(n1763) );
  oa211d1_hd U1519 ( .A(n1840), .B(n1767), .C(n148), .D(n1764), .Y(n320) );
  ao22d1_hd U1520 ( .A(b_e[1]), .B(n1765), .C(n1838), .D(C82_DATA2_1), .Y(
        n1766) );
  oa22d1_hd U1521 ( .A(n1768), .B(n1843), .C(n1767), .D(n769), .Y(n327) );
  ao22d1_hd U1522 ( .A(n1120), .B(a[21]), .C(n1830), .D(a_m[21]), .Y(n1769) );
  oa21d1_hd U1523 ( .A(n1832), .B(n1892), .C(n1769), .Y(n328) );
  ao22d1_hd U1524 ( .A(n1120), .B(a[20]), .C(n1830), .D(a_m[20]), .Y(n1770) );
  oa21d1_hd U1525 ( .A(n1832), .B(n1771), .C(n1770), .Y(n329) );
  ao22d1_hd U1526 ( .A(n1120), .B(a[19]), .C(n1830), .D(a_m[19]), .Y(n1772) );
  oa21d1_hd U1527 ( .A(n1832), .B(n1773), .C(n1772), .Y(n330) );
  oa22d1_hd U1528 ( .A(n1832), .B(n1020), .C(n1786), .D(n1773), .Y(n331) );
  ao22d1_hd U1529 ( .A(n1120), .B(a[17]), .C(n1830), .D(a_m[17]), .Y(n1774) );
  oa21d1_hd U1530 ( .A(n1832), .B(n1775), .C(n1774), .Y(n332) );
  ao22d1_hd U1531 ( .A(n1120), .B(a[16]), .C(n1830), .D(a_m[16]), .Y(n1776) );
  oa21d1_hd U1532 ( .A(n1832), .B(n1777), .C(n1776), .Y(n333) );
  oa22d1_hd U1533 ( .A(n1832), .B(n1870), .C(n1786), .D(n1777), .Y(n334) );
  ao22d1_hd U1534 ( .A(n1120), .B(a[14]), .C(n1830), .D(a_m[14]), .Y(n1778) );
  oa21d1_hd U1535 ( .A(n1832), .B(n1779), .C(n1778), .Y(n335) );
  ao22d1_hd U1536 ( .A(n1120), .B(a[13]), .C(n1830), .D(a_m[13]), .Y(n1780) );
  oa21d1_hd U1537 ( .A(n1832), .B(n1781), .C(n1780), .Y(n336) );
  oa22d1_hd U1538 ( .A(n1832), .B(n1939), .C(n1786), .D(n1781), .Y(n337) );
  ao22d1_hd U1539 ( .A(n1120), .B(a[11]), .C(n1830), .D(a_m[11]), .Y(n1782) );
  oa21d1_hd U1540 ( .A(n1832), .B(n1783), .C(n1782), .Y(n338) );
  ao22d1_hd U1541 ( .A(n1120), .B(a[10]), .C(n1830), .D(a_m[10]), .Y(n1784) );
  oa21d1_hd U1542 ( .A(n1832), .B(n1785), .C(n1784), .Y(n339) );
  oa22d1_hd U1543 ( .A(n1832), .B(n1787), .C(n1786), .D(n1785), .Y(n340) );
  ao22d1_hd U1544 ( .A(n1120), .B(a[8]), .C(n1830), .D(a_m[8]), .Y(n1788) );
  oa21d1_hd U1545 ( .A(n1832), .B(n1789), .C(n1788), .Y(n341) );
  ao22d1_hd U1546 ( .A(n1120), .B(a[7]), .C(n1830), .D(a_m[7]), .Y(n1790) );
  oa21d1_hd U1547 ( .A(n1832), .B(n1791), .C(n1790), .Y(n342) );
  ao22d1_hd U1548 ( .A(n1120), .B(a[6]), .C(n1830), .D(a_m[6]), .Y(n1792) );
  oa21d1_hd U1549 ( .A(n1832), .B(n1019), .C(n1792), .Y(n343) );
  ao22d1_hd U1550 ( .A(n1120), .B(a[5]), .C(n1830), .D(a_m[5]), .Y(n1794) );
  oa21d1_hd U1551 ( .A(n1832), .B(n1795), .C(n1794), .Y(n344) );
  ao22d1_hd U1552 ( .A(n1120), .B(a[4]), .C(n1830), .D(a_m[4]), .Y(n1796) );
  oa21d1_hd U1553 ( .A(n1832), .B(n1797), .C(n1796), .Y(n345) );
  ao22d1_hd U1554 ( .A(n1120), .B(a[3]), .C(n1830), .D(a_m[3]), .Y(n1798) );
  oa21d1_hd U1555 ( .A(n1832), .B(n1021), .C(n1798), .Y(n346) );
  ao22d1_hd U1556 ( .A(n1120), .B(a[2]), .C(n1830), .D(a_m[2]), .Y(n1799) );
  oa21d1_hd U1557 ( .A(n1832), .B(n1800), .C(n1799), .Y(n347) );
  ao22d1_hd U1558 ( .A(n1120), .B(a[1]), .C(n1830), .D(a_m[1]), .Y(n1801) );
  oa21d1_hd U1559 ( .A(n1832), .B(n1802), .C(n1801), .Y(n348) );
  nd4d1_hd U1560 ( .A(n1810), .B(n1803), .C(o_AB_ACK), .D(i_AB_STB), .Y(n1817)
         );
  ivd1_hd U1561 ( .A(o_AB_ACK), .Y(n1804) );
  ao211d1_hd U1562 ( .A(n1805), .B(n1804), .C(i_RST), .D(n2022), .Y(n350) );
  ivd1_hd U1563 ( .A(n1807), .Y(n1819) );
  nr2d1_hd U1564 ( .A(n1808), .B(n1061), .Y(n1816) );
  ao211d1_hd U1565 ( .A(state[3]), .B(state[2]), .C(n1810), .D(n1809), .Y(
        n1824) );
  nd3d1_hd U1566 ( .A(o_Z_STB), .B(i_Z_ACK), .C(n1023), .Y(n1811) );
  nd2bd1_hd U1567 ( .AN(i_RST), .B(n1811), .Y(n1849) );
  ao211d1_hd U1568 ( .A(n1850), .B(b_m[23]), .C(n1824), .D(n1849), .Y(n1812)
         );
  oa21d1_hd U1569 ( .A(n1814), .B(n1813), .C(n1812), .Y(n1815) );
  nr2d1_hd U1570 ( .A(n1816), .B(n1815), .Y(n1829) );
  oa211d1_hd U1571 ( .A(n1819), .B(n1818), .C(n1829), .D(n1817), .Y(n1845) );
  ao22d1_hd U1572 ( .A(n1821), .B(n1820), .C(n1833), .D(n1845), .Y(n1823) );
  oa22d1_hd U1573 ( .A(n1005), .B(n1823), .C(n1822), .D(n1845), .Y(n351) );
  ivd1_hd U1574 ( .A(n1824), .Y(n1826) );
  oa22d1_hd U1575 ( .A(n1005), .B(n1826), .C(n1825), .D(n1845), .Y(n352) );
  nr2d1_hd U1576 ( .A(state[0]), .B(n1847), .Y(n1828) );
  ao22d1_hd U1577 ( .A(n1120), .B(a[22]), .C(n1830), .D(a_m[22]), .Y(n1831) );
  scg16d1_hd U1578 ( .A(a_m[21]), .B(n1832), .C(n1831), .Y(n354) );
  ao22d1_hd U1579 ( .A(a_m[22]), .B(n1833), .C(n1060), .D(n1007), .Y(n1834) );
  oa21d1_hd U1580 ( .A(n1836), .B(n1835), .C(n1834), .Y(n355) );
  oa211d1_hd U1581 ( .A(n1840), .B(n1839), .C(n1838), .D(n1837), .Y(n1841) );
  oa211d1_hd U1582 ( .A(n1843), .B(n1842), .C(n148), .D(n1841), .Y(n356) );
  nr2d1_hd U1583 ( .A(n1013), .B(n1844), .Y(n1848) );
  oa22d1_hd U1584 ( .A(n1848), .B(n1847), .C(n1846), .D(n1845), .Y(n357) );
  scg20d1_hd U1585 ( .A(o_Z_STB), .B(n1023), .C(n1849), .Y(n358) );
  fad1_hd U1586 ( .A(n1853), .B(n1852), .CI(n1851), .CO(n1854), .S(
        intadd_29_B_5_) );
  ivd1_hd U1587 ( .A(n1854), .Y(n2038) );
  scg15d1_hd U1588 ( .A(n1856), .B(a_m[20]), .C(n1060), .D(n1855), .Y(n1864)
         );
  ao22d1_hd U1589 ( .A(b_m[23]), .B(n1904), .C(n1903), .D(n1857), .Y(n1858) );
  oa21d1_hd U1590 ( .A(n1058), .B(n1859), .C(n1858), .Y(n1860) );
  ivd1_hd U1591 ( .A(intadd_22_SUM_7_), .Y(n1874) );
  ao22d1_hd U1592 ( .A(b_m[23]), .B(n1009), .C(n1936), .D(n1929), .Y(n1866) );
  scg4d1_hd U1593 ( .A(n1937), .B(n1876), .C(n1055), .D(n1868), .E(n1867), .F(
        n1057), .G(n1053), .H(n1877), .Y(n1869) );
  ivd1_hd U1594 ( .A(n1871), .Y(n2035) );
  ivd1_hd U1595 ( .A(intadd_33_SUM_3_), .Y(n1886) );
  ao22d1_hd U1596 ( .A(b_m[23]), .B(n1877), .C(n1876), .D(n1929), .Y(n1878) );
  scg4d1_hd U1597 ( .A(n1937), .B(n1888), .C(n1055), .D(n1880), .E(n1879), .F(
        n1057), .G(n1053), .H(n1889), .Y(n1881) );
  ao22d1_hd U1598 ( .A(b_m[23]), .B(n1889), .C(n1888), .D(n1929), .Y(n1890) );
  scg4d1_hd U1599 ( .A(n1937), .B(n1919), .C(n1055), .D(n1920), .E(n1922), .F(
        n1057), .G(n1053), .H(n1921), .Y(n1891) );
  ivd1_hd U1600 ( .A(n1893), .Y(n2031) );
  fad1_hd U1601 ( .A(intadd_32_SUM_4_), .B(n1895), .CI(n1894), .CO(n1896), .S(
        n1893) );
  ao22d1_hd U1602 ( .A(b_m[23]), .B(n1921), .C(n1919), .D(n1929), .Y(n1897) );
  scg4d1_hd U1603 ( .A(n1937), .B(n1903), .C(n1055), .D(n1904), .E(n1906), .F(
        n1057), .G(n1053), .H(n1905), .Y(n1898) );
  ivd1_hd U1604 ( .A(n1902), .Y(n2028) );
  scg4d1_hd U1605 ( .A(n1011), .B(n1906), .C(n1012), .D(n1905), .E(n1027), .F(
        n1904), .G(n1903), .H(intadd_24_SUM_0_), .Y(n1907) );
  ao21d1_hd U1606 ( .A(n1910), .B(n1909), .C(n1908), .Y(n1917) );
  nr2d1_hd U1607 ( .A(n1061), .B(n1025), .Y(n1916) );
  ivd1_hd U1608 ( .A(n1911), .Y(n2027) );
  fad1_hd U1609 ( .A(n1021), .B(n1913), .CI(n1912), .CO(n1852), .S(n1915) );
  ivd1_hd U1610 ( .A(n1915), .Y(n1927) );
  fad1_hd U1611 ( .A(n1918), .B(n1917), .CI(n1916), .CO(n1926), .S(n1911) );
  scg4d1_hd U1612 ( .A(n1034), .B(n1922), .C(n1031), .D(n1921), .E(n1032), .F(
        n1920), .G(n1919), .H(intadd_24_SUM_4_), .Y(n1923) );
  ivd1_hd U1613 ( .A(n1924), .Y(n2026) );
  fad1_hd U1614 ( .A(n1927), .B(n1926), .CI(n1925), .CO(n1928), .S(n1924) );
  ivd1_hd U1615 ( .A(n1928), .Y(n2025) );
  ao22d1_hd U1616 ( .A(b_m[23]), .B(n1931), .C(n1930), .D(n1929), .Y(n1932) );
  scg4d1_hd U1617 ( .A(n1937), .B(n1936), .C(n1055), .D(n1935), .E(n1934), .F(
        n1057), .G(n1009), .H(n1053), .Y(n1938) );
  ivd1_hd U1618 ( .A(n1940), .Y(n2024) );
  fad1_hd U1619 ( .A(intadd_27_SUM_12_), .B(n1942), .CI(n1941), .CO(n1943), 
        .S(n1940) );
  ivd1_hd U1620 ( .A(n1943), .Y(n2023) );
  ivd1_hd U1621 ( .A(intadd_31_B_2_), .Y(n1225) );
  ivd1_hd U1622 ( .A(intadd_31_SUM_0_), .Y(n1224) );
  ivd1_hd U1623 ( .A(intadd_32_B_1_), .Y(n1222) );
  ivd1_hd U1624 ( .A(intadd_36_B_1_), .Y(n1221) );
  ivd1_hd U1625 ( .A(intadd_22_SUM_1_), .Y(n1215) );
  ivd1_hd U1626 ( .A(intadd_31_SUM_1_), .Y(n1213) );
  ivd1_hd U1627 ( .A(intadd_22_SUM_2_), .Y(n1212) );
  ivd1_hd U1628 ( .A(intadd_33_SUM_0_), .Y(n1210) );
  ivd1_hd U1629 ( .A(intadd_40_SUM_0_), .Y(n1209) );
  ivd1_hd U1630 ( .A(intadd_33_SUM_1_), .Y(n1208) );
  ivd1_hd U1631 ( .A(intadd_40_SUM_1_), .Y(n1207) );
  ivd1_hd U1632 ( .A(intadd_22_SUM_3_), .Y(n1206) );
  ivd1_hd U1633 ( .A(intadd_22_SUM_4_), .Y(n1205) );
  ivd1_hd U1634 ( .A(intadd_32_SUM_0_), .Y(n1204) );
  ivd1_hd U1635 ( .A(intadd_22_SUM_5_), .Y(n1203) );
  ivd1_hd U1636 ( .A(intadd_33_SUM_2_), .Y(n1201) );
  ivd1_hd U1637 ( .A(intadd_40_SUM_2_), .Y(n1200) );
  ivd1_hd U1638 ( .A(intadd_40_n1), .Y(n1199) );
  ivd1_hd U1639 ( .A(intadd_34_SUM_0_), .Y(n1198) );
  ivd1_hd U1640 ( .A(intadd_37_SUM_0_), .Y(n1197) );
  ivd1_hd U1641 ( .A(intadd_38_SUM_0_), .Y(n1196) );
  ivd1_hd U1642 ( .A(intadd_34_SUM_1_), .Y(n1195) );
  ivd1_hd U1643 ( .A(intadd_37_SUM_1_), .Y(n1194) );
  ivd1_hd U1644 ( .A(intadd_38_SUM_1_), .Y(n1193) );
  ivd1_hd U1645 ( .A(intadd_22_SUM_6_), .Y(n1192) );
  ivd1_hd U1646 ( .A(intadd_31_n1), .Y(n1191) );
  ivd1_hd U1647 ( .A(intadd_36_SUM_0_), .Y(n1190) );
  ivd1_hd U1648 ( .A(intadd_36_SUM_2_), .Y(n1189) );
  ivd1_hd U1649 ( .A(intadd_39_SUM_2_), .Y(n1185) );
  ivd1_hd U1650 ( .A(intadd_39_n1), .Y(n1184) );
  ivd1_hd U1651 ( .A(intadd_38_n1), .Y(n1182) );
  ivd1_hd U1652 ( .A(intadd_37_n1), .Y(n1180) );
  ivd1_hd U1653 ( .A(intadd_21_SUM_0_), .Y(n1168) );
  ivd1_hd U1654 ( .A(intadd_21_SUM_1_), .Y(n1166) );
  ivd1_hd U1655 ( .A(intadd_21_SUM_2_), .Y(n1165) );
  ivd1_hd U1656 ( .A(intadd_21_SUM_3_), .Y(n1164) );
  ivd1_hd U1657 ( .A(intadd_21_SUM_4_), .Y(n1162) );
  ivd1_hd U1658 ( .A(intadd_21_SUM_5_), .Y(n1161) );
  ivd1_hd U1659 ( .A(intadd_21_SUM_6_), .Y(n1160) );
  ivd1_hd U1660 ( .A(intadd_21_SUM_7_), .Y(n1158) );
  ivd1_hd U1661 ( .A(intadd_21_SUM_8_), .Y(n1157) );
  ivd1_hd U1662 ( .A(intadd_21_SUM_9_), .Y(n1156) );
  ivd1_hd U1663 ( .A(intadd_21_SUM_10_), .Y(n1154) );
  ivd1_hd U1664 ( .A(intadd_21_SUM_11_), .Y(n1152) );
  ivd1_hd U1665 ( .A(intadd_21_SUM_12_), .Y(n1151) );
  ivd1_hd U1666 ( .A(intadd_21_SUM_13_), .Y(n1149) );
  ivd1_hd U1667 ( .A(intadd_21_SUM_14_), .Y(n1148) );
  ivd1_hd U1668 ( .A(intadd_21_SUM_15_), .Y(n1147) );
  ivd1_hd U1669 ( .A(intadd_21_SUM_16_), .Y(n1145) );
  ivd1_hd U1670 ( .A(intadd_21_SUM_17_), .Y(n1143) );
  ivd1_hd U1671 ( .A(intadd_21_SUM_18_), .Y(n1142) );
  ivd1_hd U1672 ( .A(intadd_21_SUM_19_), .Y(n1141) );
  ivd1_hd U1673 ( .A(intadd_21_SUM_20_), .Y(n1139) );
  ivd1_hd U1674 ( .A(intadd_21_SUM_21_), .Y(n1138) );
  ivd1_hd U1675 ( .A(intadd_21_SUM_22_), .Y(n1137) );
  ivd1_hd U1676 ( .A(intadd_21_SUM_23_), .Y(n1135) );
  ivd1_hd U1677 ( .A(intadd_26_SUM_15_), .Y(n1134) );
  ivd1_hd U1678 ( .A(intadd_30_SUM_0_), .Y(n1133) );
  ivd1_hd U1679 ( .A(intadd_21_SUM_24_), .Y(n1132) );
  ivd1_hd U1680 ( .A(intadd_26_SUM_16_), .Y(n1130) );
  ivd1_hd U1681 ( .A(intadd_26_n1), .Y(n1129) );
  ivd1_hd U1682 ( .A(intadd_41_SUM_2_), .Y(n1128) );
  ivd1_hd U1683 ( .A(intadd_41_n1), .Y(n1127) );
  ivd1_hd U1684 ( .A(intadd_27_SUM_13_), .Y(n1126) );
  ivd1_hd U1685 ( .A(intadd_27_n1), .Y(n1125) );
  ivd1_hd U1686 ( .A(n1004), .Y(n1106) );
endmodule


module iir_lpf ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   r_add_AB_STB, w_add_AB_ACK, w_add_Z_STB, r_add_Z_ACK, w_mult_1_AB_ACK,
         w_mult_2_AB_ACK, w_mult_1_Z_STB, w_mult_2_Z_STB, r_mult_AB_STB,
         r_mult_Z_ACK, N18, N814, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n162, n164,
         n165, n166, n168, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n580, n811, n816, n1195, n1, n161, n163, n167, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n533, n534, n573, n574, n575, n576,
         n577, n578, n579, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721;
  wire   [31:0] r_add_A;
  wire   [31:0] r_add_B;
  wire   [31:0] w_add_Z;
  wire   [29:0] r_mult_1_A;
  wire   [31:0] r_mult_1_B;
  wire   [31:0] w_mult_1_Z;
  wire   [31:0] r_mult_2_A;
  wire   [31:0] r_mult_2_B;
  wire   [31:0] w_mult_2_Z;
  wire   [95:0] r_x_data;
  wire   [63:0] r_y_data;

  float_adder_3 add ( .i_A(r_add_A), .i_B(r_add_B), .i_AB_STB(r_add_AB_STB), 
        .o_AB_ACK(w_add_AB_ACK), .o_Z(w_add_Z), .o_Z_STB(w_add_Z_STB), 
        .i_Z_ACK(r_add_Z_ACK), .i_CLK(i_CLK), .i_RST(N18) );
  float_multiplier_1 mult_1 ( .i_A({1'b0, 1'b0, r_mult_1_A[29:22], 1'b0, 
        r_mult_1_A[20:19], 1'b0, r_mult_1_A[17:14], 1'b0, r_mult_1_A[12:0]}), 
        .i_B(r_mult_1_B), .i_AB_STB(r_mult_AB_STB), .o_AB_ACK(w_mult_1_AB_ACK), 
        .o_Z(w_mult_1_Z), .o_Z_STB(w_mult_1_Z_STB), .i_Z_ACK(r_mult_Z_ACK), 
        .i_CLK(i_CLK), .i_RST(N18) );
  float_multiplier_0 mult_2 ( .i_A({r_mult_2_A[31], 1'b0, r_mult_2_A[29:24], 
        1'b0, r_mult_2_A[22:19], 1'b0, r_mult_2_A[17:16], 1'b0, 
        r_mult_2_A[14:13], 1'b0, r_mult_2_A[11:10], 1'b0, r_mult_2_A[8:0]}), 
        .i_B(r_mult_2_B), .i_AB_STB(r_mult_AB_STB), .o_AB_ACK(w_mult_2_AB_ACK), 
        .o_Z(w_mult_2_Z), .o_Z_STB(w_mult_2_Z_STB), .i_Z_ACK(r_mult_Z_ACK), 
        .i_CLK(i_CLK), .i_RST(N18) );
  ivd1_hd U578 ( .A(i_RSTN), .Y(N18) );
  fd2qd1_hd r_mult_2_A_reg_22_ ( .D(n392), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[22]) );
  fd2qd1_hd r_mult_2_A_reg_19_ ( .D(n395), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[19]) );
  fd2qd1_hd r_mult_2_A_reg_2_ ( .D(n408), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[2]) );
  fd2qd1_hd r_mult_2_A_reg_1_ ( .D(n409), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_19_ ( .D(n420), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[19]) );
  fd2qd1_hd r_mult_1_A_reg_16_ ( .D(n422), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[16]) );
  fd2qd1_hd r_mult_1_A_reg_2_ ( .D(n435), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[2]) );
  fd2qd1_hd r_mult_1_A_reg_1_ ( .D(n436), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_0_ ( .D(n437), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[0]) );
  fd2qd1_hd r_add_B_reg_1_ ( .D(n382), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[1])
         );
  fd2qd1_hd r_add_B_reg_2_ ( .D(n381), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[2])
         );
  fd2qd1_hd r_add_B_reg_3_ ( .D(n380), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[3])
         );
  fd2qd1_hd r_add_B_reg_4_ ( .D(n379), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[4])
         );
  fd2qd1_hd r_add_B_reg_5_ ( .D(n378), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[5])
         );
  fd2qd1_hd r_add_B_reg_6_ ( .D(n377), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[6])
         );
  fd2qd1_hd r_add_B_reg_7_ ( .D(n376), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[7])
         );
  fd2qd1_hd r_add_B_reg_8_ ( .D(n375), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[8])
         );
  fd2qd1_hd r_add_B_reg_9_ ( .D(n374), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[9])
         );
  fd2qd1_hd r_add_B_reg_10_ ( .D(n373), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[10]) );
  fd2qd1_hd r_add_B_reg_11_ ( .D(n372), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[11]) );
  fd2qd1_hd r_add_B_reg_12_ ( .D(n371), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[12]) );
  fd2qd1_hd r_add_B_reg_13_ ( .D(n370), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[13]) );
  fd2qd1_hd r_add_B_reg_14_ ( .D(n369), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[14]) );
  fd2qd1_hd r_add_B_reg_15_ ( .D(n368), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[15]) );
  fd2qd1_hd r_add_B_reg_16_ ( .D(n367), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[16]) );
  fd2qd1_hd r_add_B_reg_17_ ( .D(n366), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[17]) );
  fd2qd1_hd r_add_B_reg_18_ ( .D(n365), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[18]) );
  fd2qd1_hd r_add_B_reg_19_ ( .D(n364), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[19]) );
  fd2qd1_hd r_add_B_reg_20_ ( .D(n363), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[20]) );
  fd2qd1_hd r_add_B_reg_21_ ( .D(n362), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[21]) );
  fd2qd1_hd r_add_B_reg_22_ ( .D(n361), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[22]) );
  fd2qd1_hd r_add_B_reg_23_ ( .D(n360), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[23]) );
  fd2qd1_hd r_add_B_reg_24_ ( .D(n359), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[24]) );
  fd2qd1_hd r_add_B_reg_25_ ( .D(n358), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[25]) );
  fd2qd1_hd r_add_B_reg_26_ ( .D(n357), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[26]) );
  fd2qd1_hd r_add_B_reg_27_ ( .D(n356), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[27]) );
  fd2qd1_hd r_add_B_reg_28_ ( .D(n355), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[28]) );
  fd2qd1_hd r_add_B_reg_29_ ( .D(n354), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[29]) );
  fd2qd1_hd r_add_B_reg_30_ ( .D(n353), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[30]) );
  fd2qd1_hd r_add_B_reg_31_ ( .D(n352), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[31]) );
  fd2qd1_hd r_add_B_reg_0_ ( .D(n383), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[0])
         );
  fd2qd1_hd r_x_data_reg_64_ ( .D(n95), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[64]) );
  fd2qd1_hd r_mult_2_A_reg_31_ ( .D(n385), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[31]) );
  fd2qd1_hd r_mult_2_A_reg_25_ ( .D(n390), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[25]) );
  fd2qd1_hd r_mult_2_A_reg_24_ ( .D(n391), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[24]) );
  fd2qd1_hd r_mult_2_A_reg_21_ ( .D(n393), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[21]) );
  fd2qd1_hd r_mult_2_A_reg_14_ ( .D(n398), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[14]) );
  fd2qd1_hd r_mult_2_A_reg_13_ ( .D(n399), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[13]) );
  fd2qd1_hd r_mult_2_A_reg_8_ ( .D(n402), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[8]) );
  fd2qd1_hd r_mult_2_A_reg_4_ ( .D(n406), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[4]) );
  fd2qd1_hd r_mult_1_A_reg_25_ ( .D(n415), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[25]) );
  fd2qd1_hd r_mult_1_A_reg_24_ ( .D(n416), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[24]) );
  fd2qd1_hd r_mult_1_A_reg_15_ ( .D(n423), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[15]) );
  fd2qd1_hd r_mult_1_A_reg_14_ ( .D(n424), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[14]) );
  fd2qd1_hd r_mult_1_A_reg_12_ ( .D(n425), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[12]) );
  fd2qd1_hd r_mult_1_A_reg_9_ ( .D(n428), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[9]) );
  fd2qd1_hd r_mult_1_A_reg_8_ ( .D(n429), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[8]) );
  fd2qd1_hd r_mult_1_A_reg_4_ ( .D(n433), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[4]) );
  fd2qd1_hd r_x_data_reg_65_ ( .D(n94), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[65]) );
  fd2qd1_hd r_x_data_reg_66_ ( .D(n93), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[66]) );
  fd2qd1_hd r_x_data_reg_67_ ( .D(n92), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[67]) );
  fd2qd1_hd r_x_data_reg_68_ ( .D(n91), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[68]) );
  fd2qd1_hd r_x_data_reg_69_ ( .D(n90), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[69]) );
  fd2qd1_hd r_x_data_reg_70_ ( .D(n89), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[70]) );
  fd2qd1_hd r_x_data_reg_71_ ( .D(n88), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[71]) );
  fd2qd1_hd r_x_data_reg_72_ ( .D(n87), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[72]) );
  fd2qd1_hd r_x_data_reg_73_ ( .D(n86), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[73]) );
  fd2qd1_hd r_x_data_reg_74_ ( .D(n85), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[74]) );
  fd2qd1_hd r_x_data_reg_75_ ( .D(n84), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[75]) );
  fd2qd1_hd r_x_data_reg_76_ ( .D(n83), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[76]) );
  fd2qd1_hd r_x_data_reg_77_ ( .D(n82), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[77]) );
  fd2qd1_hd r_x_data_reg_78_ ( .D(n81), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[78]) );
  fd2qd1_hd r_x_data_reg_79_ ( .D(n80), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[79]) );
  fd2qd1_hd r_x_data_reg_80_ ( .D(n79), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[80]) );
  fd2qd1_hd r_x_data_reg_81_ ( .D(n78), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[81]) );
  fd2qd1_hd r_x_data_reg_82_ ( .D(n77), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[82]) );
  fd2qd1_hd r_x_data_reg_83_ ( .D(n76), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[83]) );
  fd2qd1_hd r_x_data_reg_84_ ( .D(n75), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[84]) );
  fd2qd1_hd r_x_data_reg_85_ ( .D(n74), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[85]) );
  fd2qd1_hd r_x_data_reg_86_ ( .D(n73), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[86]) );
  fd2qd1_hd r_x_data_reg_87_ ( .D(n72), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[87]) );
  fd2qd1_hd r_x_data_reg_88_ ( .D(n71), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[88]) );
  fd2qd1_hd r_x_data_reg_89_ ( .D(n70), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[89]) );
  fd2qd1_hd r_x_data_reg_90_ ( .D(n69), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[90]) );
  fd2qd1_hd r_x_data_reg_91_ ( .D(n68), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[91]) );
  fd2qd1_hd r_x_data_reg_92_ ( .D(n67), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[92]) );
  fd2qd1_hd r_x_data_reg_93_ ( .D(n66), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[93]) );
  fd2qd1_hd r_x_data_reg_94_ ( .D(n65), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[94]) );
  fd2qd1_hd r_x_data_reg_95_ ( .D(n64), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[95]) );
  fd2qd1_hd r_mult_2_A_reg_29_ ( .D(n386), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[29]) );
  fd2qd1_hd r_mult_2_A_reg_28_ ( .D(n387), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[28]) );
  fd2qd1_hd r_mult_2_A_reg_27_ ( .D(n388), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[27]) );
  fd2qd1_hd r_mult_2_A_reg_26_ ( .D(n389), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[26]) );
  fd2qd1_hd r_mult_2_A_reg_20_ ( .D(n394), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[20]) );
  fd2qd1_hd r_mult_2_A_reg_17_ ( .D(n396), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[17]) );
  fd2qd1_hd r_mult_2_A_reg_16_ ( .D(n397), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[16]) );
  fd2qd1_hd r_mult_2_A_reg_11_ ( .D(n400), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[11]) );
  fd2qd1_hd r_mult_2_A_reg_10_ ( .D(n401), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[10]) );
  fd2qd1_hd r_mult_2_A_reg_7_ ( .D(n403), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[7]) );
  fd2qd1_hd r_mult_2_A_reg_6_ ( .D(n404), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[6]) );
  fd2qd1_hd r_mult_2_A_reg_5_ ( .D(n405), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[5]) );
  fd2qd1_hd r_mult_2_A_reg_3_ ( .D(n407), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[3]) );
  fd2qd1_hd r_mult_2_A_reg_0_ ( .D(n410), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[0]) );
  fd2qd1_hd r_mult_1_A_reg_29_ ( .D(n411), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_28_ ( .D(n412), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[28]) );
  fd2qd1_hd r_mult_1_A_reg_27_ ( .D(n413), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[27]) );
  fd2qd1_hd r_mult_1_A_reg_26_ ( .D(n414), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[26]) );
  fd2qd1_hd r_mult_1_A_reg_23_ ( .D(n417), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[23]) );
  fd2qd1_hd r_mult_1_A_reg_22_ ( .D(n418), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[22]) );
  fd2qd1_hd r_mult_1_A_reg_20_ ( .D(n419), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[20]) );
  fd2qd1_hd r_mult_1_A_reg_17_ ( .D(n421), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[17]) );
  fd2qd1_hd r_mult_1_A_reg_11_ ( .D(n426), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[11]) );
  fd2qd1_hd r_mult_1_A_reg_10_ ( .D(n427), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[10]) );
  fd2qd1_hd r_mult_1_A_reg_7_ ( .D(n430), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[7]) );
  fd2qd1_hd r_mult_1_A_reg_6_ ( .D(n431), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[6]) );
  fd2qd1_hd r_mult_1_A_reg_5_ ( .D(n432), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[5]) );
  fd2qd1_hd r_mult_1_A_reg_3_ ( .D(n434), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[3]) );
  fd2qd1_hd r_add_A_reg_0_ ( .D(n571), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[0])
         );
  fd2qd1_hd r_mult_2_B_reg_31_ ( .D(n536), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[31]) );
  fd2qd1_hd r_mult_2_B_reg_30_ ( .D(n439), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_30_ ( .D(n470), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[30]) );
  fd2qd1_hd r_mult_2_B_reg_29_ ( .D(n440), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[29]) );
  fd2qd1_hd r_mult_1_B_reg_29_ ( .D(n471), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[29]) );
  fd2qd1_hd r_mult_2_B_reg_28_ ( .D(n441), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[28]) );
  fd2qd1_hd r_mult_1_B_reg_28_ ( .D(n472), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[28]) );
  fd2qd1_hd r_mult_2_B_reg_27_ ( .D(n442), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[27]) );
  fd2qd1_hd r_mult_1_B_reg_27_ ( .D(n473), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[27]) );
  fd2qd1_hd r_mult_2_B_reg_26_ ( .D(n443), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[26]) );
  fd2qd1_hd r_mult_1_B_reg_26_ ( .D(n474), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[26]) );
  fd2qd1_hd r_mult_2_B_reg_25_ ( .D(n444), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[25]) );
  fd2qd1_hd r_mult_1_B_reg_25_ ( .D(n475), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[25]) );
  fd2qd1_hd r_mult_2_B_reg_24_ ( .D(n445), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[24]) );
  fd2qd1_hd r_mult_1_B_reg_24_ ( .D(n476), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[24]) );
  fd2qd1_hd r_mult_2_B_reg_23_ ( .D(n446), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[23]) );
  fd2qd1_hd r_mult_1_B_reg_23_ ( .D(n477), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[23]) );
  fd2qd1_hd r_mult_2_B_reg_22_ ( .D(n447), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[22]) );
  fd2qd1_hd r_mult_1_B_reg_22_ ( .D(n478), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[22]) );
  fd2qd1_hd r_mult_2_B_reg_21_ ( .D(n448), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[21]) );
  fd2qd1_hd r_mult_1_B_reg_21_ ( .D(n479), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[21]) );
  fd2qd1_hd r_mult_2_B_reg_20_ ( .D(n449), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[20]) );
  fd2qd1_hd r_mult_1_B_reg_20_ ( .D(n480), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[20]) );
  fd2qd1_hd r_mult_2_B_reg_19_ ( .D(n450), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[19]) );
  fd2qd1_hd r_mult_1_B_reg_19_ ( .D(n481), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[19]) );
  fd2qd1_hd r_mult_2_B_reg_18_ ( .D(n451), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[18]) );
  fd2qd1_hd r_mult_1_B_reg_18_ ( .D(n482), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[18]) );
  fd2qd1_hd r_mult_2_B_reg_17_ ( .D(n452), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[17]) );
  fd2qd1_hd r_mult_1_B_reg_17_ ( .D(n483), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[17]) );
  fd2qd1_hd r_mult_2_B_reg_16_ ( .D(n453), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[16]) );
  fd2qd1_hd r_mult_1_B_reg_16_ ( .D(n484), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[16]) );
  fd2qd1_hd r_mult_2_B_reg_15_ ( .D(n454), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[15]) );
  fd2qd1_hd r_mult_1_B_reg_15_ ( .D(n485), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[15]) );
  fd2qd1_hd r_mult_2_B_reg_14_ ( .D(n455), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[14]) );
  fd2qd1_hd r_mult_1_B_reg_14_ ( .D(n486), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[14]) );
  fd2qd1_hd r_mult_2_B_reg_13_ ( .D(n456), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[13]) );
  fd2qd1_hd r_mult_1_B_reg_13_ ( .D(n487), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[13]) );
  fd2qd1_hd r_mult_2_B_reg_12_ ( .D(n457), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[12]) );
  fd2qd1_hd r_mult_1_B_reg_12_ ( .D(n488), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[12]) );
  fd2qd1_hd r_mult_2_B_reg_11_ ( .D(n458), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[11]) );
  fd2qd1_hd r_mult_1_B_reg_11_ ( .D(n489), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[11]) );
  fd2qd1_hd r_mult_2_B_reg_10_ ( .D(n459), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[10]) );
  fd2qd1_hd r_mult_1_B_reg_10_ ( .D(n490), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[10]) );
  fd2qd1_hd r_mult_2_B_reg_9_ ( .D(n460), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[9]) );
  fd2qd1_hd r_mult_1_B_reg_9_ ( .D(n491), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[9]) );
  fd2qd1_hd r_mult_2_B_reg_8_ ( .D(n461), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[8]) );
  fd2qd1_hd r_mult_1_B_reg_8_ ( .D(n492), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[8]) );
  fd2qd1_hd r_mult_2_B_reg_7_ ( .D(n462), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[7]) );
  fd2qd1_hd r_mult_1_B_reg_7_ ( .D(n493), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[7]) );
  fd2qd1_hd r_mult_2_B_reg_6_ ( .D(n463), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[6]) );
  fd2qd1_hd r_mult_1_B_reg_6_ ( .D(n494), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[6]) );
  fd2qd1_hd r_mult_2_B_reg_5_ ( .D(n464), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[5]) );
  fd2qd1_hd r_mult_1_B_reg_5_ ( .D(n495), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[5]) );
  fd2qd1_hd r_mult_2_B_reg_4_ ( .D(n465), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[4]) );
  fd2qd1_hd r_mult_1_B_reg_4_ ( .D(n496), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[4]) );
  fd2qd1_hd r_mult_2_B_reg_3_ ( .D(n466), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[3]) );
  fd2qd1_hd r_mult_1_B_reg_3_ ( .D(n497), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[3]) );
  fd2qd1_hd r_mult_2_B_reg_2_ ( .D(n467), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[2]) );
  fd2qd1_hd r_mult_1_B_reg_2_ ( .D(n498), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[2]) );
  fd2qd1_hd r_mult_2_B_reg_1_ ( .D(n468), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[1]) );
  fd2qd1_hd r_mult_1_B_reg_1_ ( .D(n499), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[1]) );
  fd2qd1_hd r_mult_2_B_reg_0_ ( .D(n469), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[0]) );
  fd2qd1_hd r_mult_1_B_reg_0_ ( .D(n500), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[0]) );
  fd2qd1_hd r_add_A_reg_1_ ( .D(n530), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[1])
         );
  fd2qd1_hd r_add_A_reg_2_ ( .D(n529), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[2])
         );
  fd2qd1_hd r_add_A_reg_3_ ( .D(n528), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[3])
         );
  fd2qd1_hd r_add_A_reg_4_ ( .D(n527), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[4])
         );
  fd2qd1_hd r_add_A_reg_5_ ( .D(n526), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[5])
         );
  fd2qd1_hd r_add_A_reg_6_ ( .D(n525), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[6])
         );
  fd2qd1_hd r_add_A_reg_7_ ( .D(n524), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[7])
         );
  fd2qd1_hd r_add_A_reg_8_ ( .D(n523), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[8])
         );
  fd2qd1_hd r_add_A_reg_9_ ( .D(n522), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[9])
         );
  fd2qd1_hd r_add_A_reg_10_ ( .D(n521), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[10]) );
  fd2qd1_hd r_add_A_reg_11_ ( .D(n520), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[11]) );
  fd2qd1_hd r_add_A_reg_12_ ( .D(n519), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[12]) );
  fd2qd1_hd r_add_A_reg_13_ ( .D(n518), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[13]) );
  fd2qd1_hd r_add_A_reg_14_ ( .D(n517), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[14]) );
  fd2qd1_hd r_add_A_reg_15_ ( .D(n516), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[15]) );
  fd2qd1_hd r_add_A_reg_16_ ( .D(n515), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[16]) );
  fd2qd1_hd r_add_A_reg_17_ ( .D(n514), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[17]) );
  fd2qd1_hd r_add_A_reg_18_ ( .D(n513), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[18]) );
  fd2qd1_hd r_add_A_reg_19_ ( .D(n512), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[19]) );
  fd2qd1_hd r_add_A_reg_20_ ( .D(n511), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[20]) );
  fd2qd1_hd r_add_A_reg_21_ ( .D(n510), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[21]) );
  fd2qd1_hd r_add_A_reg_22_ ( .D(n509), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[22]) );
  fd2qd1_hd r_add_A_reg_23_ ( .D(n508), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[23]) );
  fd2qd1_hd r_add_A_reg_24_ ( .D(n507), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[24]) );
  fd2qd1_hd r_add_A_reg_25_ ( .D(n506), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[25]) );
  fd2qd1_hd r_add_A_reg_26_ ( .D(n505), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[26]) );
  fd2qd1_hd r_add_A_reg_27_ ( .D(n504), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[27]) );
  fd2qd1_hd r_add_A_reg_28_ ( .D(n503), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[28]) );
  fd2qd1_hd r_add_A_reg_29_ ( .D(n502), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[29]) );
  fd2qd1_hd r_add_A_reg_30_ ( .D(n501), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[30]) );
  fd2qd1_hd r_mult_1_B_reg_31_ ( .D(n568), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[31]) );
  fd2qd1_hd r_add_A_reg_31_ ( .D(n570), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[31]) );
  fd2qd1_hd r_y_data_reg_62_ ( .D(n62), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[62]) );
  fd2qd1_hd r_y_data_reg_61_ ( .D(n60), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[61]) );
  fd2qd1_hd r_y_data_reg_60_ ( .D(n58), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[60]) );
  fd2qd1_hd r_y_data_reg_59_ ( .D(n56), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[59]) );
  fd2qd1_hd r_y_data_reg_58_ ( .D(n54), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[58]) );
  fd2qd1_hd r_y_data_reg_57_ ( .D(n52), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[57]) );
  fd2qd1_hd r_y_data_reg_56_ ( .D(n50), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[56]) );
  fd2qd1_hd r_y_data_reg_55_ ( .D(n48), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[55]) );
  fd2qd1_hd r_y_data_reg_54_ ( .D(n46), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[54]) );
  fd2qd1_hd r_y_data_reg_53_ ( .D(n44), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[53]) );
  fd2qd1_hd r_y_data_reg_52_ ( .D(n42), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[52]) );
  fd2qd1_hd r_y_data_reg_51_ ( .D(n40), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[51]) );
  fd2qd1_hd r_y_data_reg_50_ ( .D(n38), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[50]) );
  fd2qd1_hd r_y_data_reg_49_ ( .D(n36), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[49]) );
  fd2qd1_hd r_y_data_reg_48_ ( .D(n34), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[48]) );
  fd2qd1_hd r_y_data_reg_47_ ( .D(n32), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[47]) );
  fd2qd1_hd r_y_data_reg_46_ ( .D(n30), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[46]) );
  fd2qd1_hd r_y_data_reg_45_ ( .D(n28), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[45]) );
  fd2qd1_hd r_y_data_reg_44_ ( .D(n26), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[44]) );
  fd2qd1_hd r_y_data_reg_43_ ( .D(n24), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[43]) );
  fd2qd1_hd r_y_data_reg_42_ ( .D(n22), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[42]) );
  fd2qd1_hd r_y_data_reg_41_ ( .D(n20), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[41]) );
  fd2qd1_hd r_y_data_reg_40_ ( .D(n18), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[40]) );
  fd2qd1_hd r_y_data_reg_39_ ( .D(n16), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[39]) );
  fd2qd1_hd r_y_data_reg_38_ ( .D(n14), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[38]) );
  fd2qd1_hd r_y_data_reg_37_ ( .D(n12), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[37]) );
  fd2qd1_hd r_y_data_reg_36_ ( .D(n10), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[36]) );
  fd2qd1_hd r_y_data_reg_35_ ( .D(n8), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[35]) );
  fd2qd1_hd r_y_data_reg_34_ ( .D(n6), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[34]) );
  fd2qd1_hd r_y_data_reg_33_ ( .D(n4), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[33]) );
  fd2qd1_hd r_y_data_reg_32_ ( .D(n2), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[32]) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(n569), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[31]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(n537), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(n538), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(n539), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(n540), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(n541), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(n542), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(n543), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(n544), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(n545), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(n546), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(n547), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(n548), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(n549), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(n550), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(n551), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(n552), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(n553), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(n554), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(n555), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(n556), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(n557), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(n558), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[9]) );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(n559), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[8]) );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(n560), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[7]) );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(n561), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[6]) );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(n562), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[5]) );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(n563), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[4]) );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(n564), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[3]) );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(n565), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[2]) );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(n566), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[1]) );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(n567), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[0]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(n165), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(n63), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(n61), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(n59), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(n57), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(n55), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(n53), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(n51), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(n49), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(n47), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(n45), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(n43), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(n41), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(n39), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(n37), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(n35), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(n33), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(n31), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(n29), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(n27), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(n25), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(n23), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(n21), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(n19), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(n17), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(n15), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(n13), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(n11), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(n9), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[3])
         );
  fd2qd1_hd r_y_data_reg_2_ ( .D(n7), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[2])
         );
  fd2qd1_hd r_y_data_reg_1_ ( .D(n5), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[1])
         );
  fd2qd1_hd r_y_data_reg_0_ ( .D(n3), .CK(i_CLK), .RN(i_RSTN), .Q(r_y_data[0])
         );
  fd2qd1_hd r_add_Z_ACK_reg ( .D(n531), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_Z_ACK) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n384), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA_VALID) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n163), .E(N814), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_mult_Z_ACK_reg ( .D(n532), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_Z_ACK) );
  fd2qd1_hd r_mult_AB_STB_reg ( .D(n438), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_AB_STB) );
  fd2qd1_hd r_add_AB_STB_reg ( .D(n535), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_AB_STB) );
  fd3d1_hd r_pstate_reg_1_ ( .D(n160), .CK(i_CLK), .SN(i_RSTN), .QN(n580) );
  fd3d1_hd r_pstate_reg_0_ ( .D(n168), .CK(i_CLK), .SN(i_RSTN), .Q(n199), .QN(
        n1195) );
  fd3d1_hd r_counter_reg_0_ ( .D(n162), .CK(i_CLK), .SN(i_RSTN), .Q(n200), 
        .QN(n811) );
  fd3d1_hd r_counter_reg_1_ ( .D(n166), .CK(i_CLK), .SN(i_RSTN), .Q(n170), 
        .QN(n816) );
  fd2d1_hd r_x_data_reg_41_ ( .D(n118), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[41]), .QN(n189) );
  fd2d1_hd r_x_data_reg_39_ ( .D(n120), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[39]), .QN(n191) );
  fd2d1_hd r_x_data_reg_37_ ( .D(n122), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[37]), .QN(n193) );
  fd2d1_hd r_x_data_reg_36_ ( .D(n123), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[36]), .QN(n194) );
  fd2d1_hd r_x_data_reg_34_ ( .D(n125), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[34]), .QN(n196) );
  fd2d1_hd r_x_data_reg_33_ ( .D(n126), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[33]), .QN(n197) );
  fd2d1_hd r_x_data_reg_32_ ( .D(n127), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[32]), .QN(n198) );
  fd2d1_hd r_x_data_reg_59_ ( .D(n100), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[59]), .QN(n171) );
  fd2d1_hd r_x_data_reg_58_ ( .D(n101), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[58]), .QN(n172) );
  fd2d1_hd r_x_data_reg_57_ ( .D(n102), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[57]), .QN(n173) );
  fd2d1_hd r_x_data_reg_54_ ( .D(n105), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[54]), .QN(n176) );
  fd2d1_hd r_x_data_reg_51_ ( .D(n108), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[51]), .QN(n179) );
  fd2d1_hd r_x_data_reg_50_ ( .D(n109), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[50]), .QN(n180) );
  fd2d1_hd r_x_data_reg_48_ ( .D(n111), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[48]), .QN(n182) );
  fd2d1_hd r_x_data_reg_45_ ( .D(n114), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[45]), .QN(n185) );
  fd2d1_hd r_x_data_reg_44_ ( .D(n115), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[44]), .QN(n186) );
  fd2d1_hd r_x_data_reg_40_ ( .D(n119), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[40]), .QN(n190) );
  fd2d1_hd r_x_data_reg_38_ ( .D(n121), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[38]), .QN(n192) );
  fd2d1_hd r_x_data_reg_35_ ( .D(n124), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[35]), .QN(n195) );
  fd2d1_hd r_x_data_reg_56_ ( .D(n103), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[56]), .QN(n174) );
  fd2d1_hd r_x_data_reg_55_ ( .D(n104), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[55]), .QN(n175) );
  fd2d1_hd r_x_data_reg_53_ ( .D(n106), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[53]), .QN(n177) );
  fd2d1_hd r_x_data_reg_52_ ( .D(n107), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[52]), .QN(n178) );
  fd2d1_hd r_x_data_reg_49_ ( .D(n110), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[49]), .QN(n181) );
  fd2d1_hd r_x_data_reg_47_ ( .D(n112), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[47]), .QN(n183) );
  fd2d1_hd r_x_data_reg_46_ ( .D(n113), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[46]), .QN(n184) );
  fd2d1_hd r_x_data_reg_43_ ( .D(n116), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[43]), .QN(n187) );
  fd2d1_hd r_x_data_reg_42_ ( .D(n117), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[42]), .QN(n188) );
  fd2d1_hd r_x_data_reg_27_ ( .D(n132), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[27]), .QN(n201) );
  fd2d1_hd r_x_data_reg_26_ ( .D(n133), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[26]), .QN(n202) );
  fd2d1_hd r_x_data_reg_25_ ( .D(n134), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[25]), .QN(n203) );
  fd2d1_hd r_x_data_reg_24_ ( .D(n135), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[24]), .QN(n204) );
  fd2d1_hd r_x_data_reg_23_ ( .D(n136), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[23]), .QN(n205) );
  fd2d1_hd r_x_data_reg_22_ ( .D(n137), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[22]), .QN(n206) );
  fd2d1_hd r_x_data_reg_21_ ( .D(n138), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[21]), .QN(n207) );
  fd2d1_hd r_x_data_reg_20_ ( .D(n139), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[20]), .QN(n208) );
  fd2d1_hd r_x_data_reg_19_ ( .D(n140), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[19]), .QN(n209) );
  fd2d1_hd r_x_data_reg_18_ ( .D(n141), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[18]), .QN(n210) );
  fd2d1_hd r_x_data_reg_17_ ( .D(n142), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[17]), .QN(n211) );
  fd2d1_hd r_x_data_reg_16_ ( .D(n143), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[16]), .QN(n212) );
  fd2d1_hd r_x_data_reg_15_ ( .D(n144), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[15]), .QN(n213) );
  fd2d1_hd r_x_data_reg_14_ ( .D(n145), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[14]), .QN(n214) );
  fd2d1_hd r_x_data_reg_13_ ( .D(n146), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[13]), .QN(n215) );
  fd2d1_hd r_x_data_reg_12_ ( .D(n147), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[12]), .QN(n216) );
  fd2d1_hd r_x_data_reg_11_ ( .D(n148), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[11]), .QN(n217) );
  fd2d1_hd r_x_data_reg_10_ ( .D(n149), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[10]), .QN(n218) );
  fd2d1_hd r_x_data_reg_9_ ( .D(n150), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[9]), .QN(n219) );
  fd2d1_hd r_x_data_reg_8_ ( .D(n151), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[8]), .QN(n220) );
  fd2d1_hd r_x_data_reg_7_ ( .D(n152), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[7]), .QN(n221) );
  fd2d1_hd r_x_data_reg_6_ ( .D(n153), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[6]), .QN(n222) );
  fd2d1_hd r_x_data_reg_5_ ( .D(n154), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[5]), .QN(n223) );
  fd2d1_hd r_x_data_reg_4_ ( .D(n155), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[4]), .QN(n224) );
  fd2d1_hd r_x_data_reg_3_ ( .D(n156), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[3]), .QN(n225) );
  fd2d1_hd r_x_data_reg_2_ ( .D(n157), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[2]), .QN(n226) );
  fd2d1_hd r_x_data_reg_1_ ( .D(n158), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[1]), .QN(n227) );
  fd2d1_hd r_x_data_reg_0_ ( .D(n159), .CK(i_CLK), .RN(i_RSTN), .Q(r_x_data[0]), .QN(n228) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(n96), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[63]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(n97), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(n98), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_y_data_reg_63_ ( .D(n164), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[63]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(n130), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(n99), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(n128), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[31]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(n129), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(n131), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[28]) );
  clknd2d1_hd U590 ( .A(w_add_Z_STB), .B(n274), .Y(n637) );
  clknd2d1_hd U591 ( .A(n170), .B(n811), .Y(n642) );
  clknd2d1_hd U592 ( .A(n275), .B(n634), .Y(n278) );
  clknd2d1_hd U593 ( .A(n283), .B(n270), .Y(n282) );
  clknd2d1_hd U594 ( .A(n199), .B(n580), .Y(n641) );
  nd2d2_hd U595 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(n572) );
  clknd2d1_hd U596 ( .A(n637), .B(n638), .Y(n631) );
  nid2_hd U597 ( .A(n707), .Y(n229) );
  clknd2d4_hd U598 ( .A(n274), .B(n275), .Y(n721) );
  clknd2d1_hd U599 ( .A(n1), .B(i_X_DATA[0]), .Y(n263) );
  clknd2d1_hd U600 ( .A(n1), .B(i_X_DATA[1]), .Y(n262) );
  clknd2d1_hd U601 ( .A(n1), .B(i_X_DATA[2]), .Y(n261) );
  clknd2d1_hd U602 ( .A(n1), .B(i_X_DATA[3]), .Y(n260) );
  clknd2d1_hd U603 ( .A(n1), .B(i_X_DATA[4]), .Y(n259) );
  clknd2d1_hd U604 ( .A(n1), .B(i_X_DATA[5]), .Y(n258) );
  clknd2d1_hd U605 ( .A(n1), .B(i_X_DATA[6]), .Y(n257) );
  clknd2d1_hd U606 ( .A(n1), .B(i_X_DATA[7]), .Y(n256) );
  clknd2d1_hd U607 ( .A(n1), .B(i_X_DATA[8]), .Y(n255) );
  clknd2d1_hd U608 ( .A(n1), .B(i_X_DATA[9]), .Y(n254) );
  clknd2d1_hd U609 ( .A(n1), .B(i_X_DATA[10]), .Y(n253) );
  clknd2d1_hd U610 ( .A(n1), .B(i_X_DATA[11]), .Y(n252) );
  clknd2d1_hd U611 ( .A(n1), .B(i_X_DATA[12]), .Y(n251) );
  clknd2d1_hd U612 ( .A(n1), .B(i_X_DATA[13]), .Y(n250) );
  clknd2d1_hd U613 ( .A(n1), .B(i_X_DATA[14]), .Y(n249) );
  clknd2d1_hd U614 ( .A(n1), .B(i_X_DATA[15]), .Y(n248) );
  clknd2d1_hd U615 ( .A(n1), .B(i_X_DATA[16]), .Y(n247) );
  clknd2d1_hd U616 ( .A(n1), .B(i_X_DATA[17]), .Y(n246) );
  clknd2d1_hd U617 ( .A(n1), .B(i_X_DATA[18]), .Y(n245) );
  clknd2d1_hd U618 ( .A(n1), .B(i_X_DATA[19]), .Y(n244) );
  clknd2d1_hd U619 ( .A(n1), .B(i_X_DATA[20]), .Y(n243) );
  clknd2d1_hd U620 ( .A(n1), .B(i_X_DATA[21]), .Y(n242) );
  clknd2d1_hd U621 ( .A(n1), .B(i_X_DATA[22]), .Y(n241) );
  clknd2d1_hd U622 ( .A(n1), .B(i_X_DATA[23]), .Y(n240) );
  clknd2d1_hd U623 ( .A(n1), .B(i_X_DATA[24]), .Y(n239) );
  clknd2d1_hd U624 ( .A(n1), .B(i_X_DATA[25]), .Y(n238) );
  clknd2d1_hd U625 ( .A(n1), .B(i_X_DATA[26]), .Y(n237) );
  clknd2d1_hd U626 ( .A(n1), .B(i_X_DATA[27]), .Y(n236) );
  clknd2d1_hd U627 ( .A(w_mult_2_Z_STB), .B(w_mult_1_Z_STB), .Y(n264) );
  clknd2d1_hd U628 ( .A(n639), .B(r_mult_AB_STB), .Y(n287) );
  clknd2d1_hd U629 ( .A(n281), .B(n280), .Y(n384) );
  nid6_hd U630 ( .A(n715), .Y(n232) );
  ivd3_hd U631 ( .A(n163), .Y(n235) );
  ivd3_hd U632 ( .A(n572), .Y(n161) );
  ivd6_hd U633 ( .A(n572), .Y(n1) );
  nid6_hd U634 ( .A(n572), .Y(n163) );
  nr2d4_hd U635 ( .A(n232), .B(n350), .Y(n286) );
  nid6_hd U636 ( .A(n705), .Y(n169) );
  ad2d2_hd U637 ( .A(n285), .B(n284), .Y(n350) );
  scg2d1_hd U638 ( .A(n235), .B(i_X_DATA[30]), .C(r_x_data[30]), .D(n572), .Y(
        n129) );
  scg2d1_hd U639 ( .A(n235), .B(i_X_DATA[31]), .C(r_x_data[31]), .D(n572), .Y(
        n128) );
  or2bd2_hd U640 ( .B(n716), .AN(n721), .Y(n279) );
  nid4_hd U641 ( .A(n717), .Y(n234) );
  nid4_hd U642 ( .A(n714), .Y(n231) );
  ivd3_hd U643 ( .A(n643), .Y(n710) );
  ivd3_hd U644 ( .A(n350), .Y(n167) );
  scg10d1_hd U645 ( .A(n635), .B(r_mult_Z_ACK), .C(n634), .D(n633), .Y(n532)
         );
  nr2d4_hd U646 ( .A(n277), .B(n639), .Y(n715) );
  scg2d1_hd U647 ( .A(n235), .B(i_X_DATA[28]), .C(r_x_data[28]), .D(n163), .Y(
        n131) );
  scg10d1_hd U648 ( .A(n163), .B(o_Y_DATA[12]), .C(r_y_data[12]), .D(n1), .Y(
        n27) );
  scg10d1_hd U649 ( .A(n163), .B(r_x_data[30]), .C(r_x_data[62]), .D(n1), .Y(
        n97) );
  scg10d1_hd U650 ( .A(n163), .B(o_Y_DATA[5]), .C(r_y_data[5]), .D(n1), .Y(n13) );
  scg10d1_hd U651 ( .A(n163), .B(r_x_data[63]), .C(r_x_data[95]), .D(n161), 
        .Y(n64) );
  scg10d1_hd U652 ( .A(n163), .B(o_Y_DATA[6]), .C(r_y_data[6]), .D(n1), .Y(n15) );
  scg2d1_hd U653 ( .A(n1), .B(i_X_DATA[29]), .C(r_x_data[29]), .D(n163), .Y(
        n130) );
  scg10d1_hd U654 ( .A(n163), .B(r_x_data[31]), .C(r_x_data[63]), .D(n1), .Y(
        n96) );
  scg10d1_hd U655 ( .A(n163), .B(r_x_data[28]), .C(r_x_data[60]), .D(n161), 
        .Y(n99) );
  scg10d1_hd U656 ( .A(n163), .B(r_x_data[47]), .C(r_x_data[79]), .D(n161), 
        .Y(n80) );
  scg10d1_hd U657 ( .A(n163), .B(o_Y_DATA[7]), .C(r_y_data[7]), .D(n1), .Y(n17) );
  scg10d1_hd U658 ( .A(n163), .B(r_x_data[49]), .C(r_x_data[81]), .D(n161), 
        .Y(n78) );
  scg10d1_hd U659 ( .A(n163), .B(o_Y_DATA[14]), .C(r_y_data[14]), .D(n1), .Y(
        n31) );
  scg10d1_hd U660 ( .A(n163), .B(o_Y_DATA[11]), .C(r_y_data[11]), .D(n1), .Y(
        n25) );
  scg10d1_hd U661 ( .A(n163), .B(r_y_data[31]), .C(r_y_data[63]), .D(n1), .Y(
        n164) );
  scg10d1_hd U662 ( .A(n163), .B(o_Y_DATA[8]), .C(r_y_data[8]), .D(n1), .Y(n19) );
  scg10d1_hd U663 ( .A(n163), .B(o_Y_DATA[13]), .C(r_y_data[13]), .D(n1), .Y(
        n29) );
  scg10d1_hd U664 ( .A(n163), .B(r_x_data[48]), .C(r_x_data[80]), .D(n161), 
        .Y(n79) );
  scg10d1_hd U665 ( .A(n163), .B(o_Y_DATA[9]), .C(r_y_data[9]), .D(n1), .Y(n21) );
  scg10d1_hd U666 ( .A(n163), .B(r_x_data[50]), .C(r_x_data[82]), .D(n161), 
        .Y(n77) );
  scg10d1_hd U667 ( .A(n163), .B(o_Y_DATA[10]), .C(r_y_data[10]), .D(n1), .Y(
        n23) );
  scg10d1_hd U668 ( .A(n163), .B(r_x_data[58]), .C(r_x_data[90]), .D(n161), 
        .Y(n69) );
  scg10d1_hd U669 ( .A(n163), .B(r_x_data[57]), .C(r_x_data[89]), .D(n161), 
        .Y(n70) );
  scg10d1_hd U670 ( .A(n163), .B(r_x_data[59]), .C(r_x_data[91]), .D(n161), 
        .Y(n68) );
  scg10d1_hd U671 ( .A(n163), .B(r_x_data[56]), .C(r_x_data[88]), .D(n161), 
        .Y(n71) );
  scg10d1_hd U672 ( .A(n163), .B(o_Y_DATA[31]), .C(r_y_data[31]), .D(n1), .Y(
        n165) );
  scg10d1_hd U673 ( .A(n163), .B(r_x_data[55]), .C(r_x_data[87]), .D(n161), 
        .Y(n72) );
  scg10d1_hd U674 ( .A(n163), .B(r_x_data[54]), .C(r_x_data[86]), .D(n161), 
        .Y(n73) );
  scg10d1_hd U675 ( .A(n163), .B(r_x_data[53]), .C(r_x_data[85]), .D(n161), 
        .Y(n74) );
  scg10d1_hd U676 ( .A(n163), .B(r_x_data[60]), .C(r_x_data[92]), .D(n161), 
        .Y(n67) );
  scg10d1_hd U677 ( .A(n163), .B(r_x_data[61]), .C(r_x_data[93]), .D(n161), 
        .Y(n66) );
  scg10d1_hd U678 ( .A(n163), .B(r_x_data[62]), .C(r_x_data[94]), .D(n161), 
        .Y(n65) );
  scg10d1_hd U679 ( .A(n163), .B(o_Y_DATA[0]), .C(r_y_data[0]), .D(n1), .Y(n3)
         );
  scg10d1_hd U680 ( .A(n163), .B(r_x_data[29]), .C(r_x_data[61]), .D(n1), .Y(
        n98) );
  scg10d1_hd U681 ( .A(n163), .B(o_Y_DATA[1]), .C(r_y_data[1]), .D(n161), .Y(
        n5) );
  scg10d1_hd U682 ( .A(n163), .B(o_Y_DATA[2]), .C(r_y_data[2]), .D(n161), .Y(
        n7) );
  scg10d1_hd U683 ( .A(n163), .B(r_x_data[52]), .C(r_x_data[84]), .D(n161), 
        .Y(n75) );
  scg10d1_hd U684 ( .A(n163), .B(o_Y_DATA[3]), .C(r_y_data[3]), .D(n1), .Y(n9)
         );
  scg10d1_hd U685 ( .A(n163), .B(o_Y_DATA[4]), .C(r_y_data[4]), .D(n1), .Y(n11) );
  scg10d1_hd U686 ( .A(n163), .B(r_x_data[51]), .C(r_x_data[83]), .D(n161), 
        .Y(n76) );
  scg10d1_hd U687 ( .A(n163), .B(r_y_data[7]), .C(r_y_data[39]), .D(n1), .Y(
        n16) );
  scg10d1_hd U688 ( .A(n163), .B(r_y_data[8]), .C(r_y_data[40]), .D(n1), .Y(
        n18) );
  scg10d1_hd U689 ( .A(n163), .B(o_Y_DATA[29]), .C(r_y_data[29]), .D(n161), 
        .Y(n61) );
  scg10d1_hd U690 ( .A(n163), .B(r_y_data[9]), .C(r_y_data[41]), .D(n1), .Y(
        n20) );
  scg10d1_hd U691 ( .A(n163), .B(r_y_data[10]), .C(r_y_data[42]), .D(n1), .Y(
        n22) );
  scg10d1_hd U692 ( .A(n163), .B(o_Y_DATA[25]), .C(r_y_data[25]), .D(n161), 
        .Y(n53) );
  scg10d1_hd U693 ( .A(n163), .B(r_y_data[11]), .C(r_y_data[43]), .D(n1), .Y(
        n24) );
  scg10d1_hd U694 ( .A(n163), .B(r_y_data[12]), .C(r_y_data[44]), .D(n1), .Y(
        n26) );
  scg10d1_hd U695 ( .A(n163), .B(r_y_data[13]), .C(r_y_data[45]), .D(n1), .Y(
        n28) );
  scg10d1_hd U696 ( .A(n163), .B(r_x_data[38]), .C(r_x_data[70]), .D(n1), .Y(
        n89) );
  scg10d1_hd U697 ( .A(n163), .B(r_y_data[14]), .C(r_y_data[46]), .D(n1), .Y(
        n30) );
  scg10d1_hd U698 ( .A(n163), .B(r_y_data[15]), .C(r_y_data[47]), .D(n1), .Y(
        n32) );
  scg10d1_hd U699 ( .A(n163), .B(r_y_data[16]), .C(r_y_data[48]), .D(n1), .Y(
        n34) );
  scg10d1_hd U700 ( .A(n163), .B(r_y_data[17]), .C(r_y_data[49]), .D(n1), .Y(
        n36) );
  scg10d1_hd U701 ( .A(n163), .B(r_y_data[18]), .C(r_y_data[50]), .D(n1), .Y(
        n38) );
  scg10d1_hd U702 ( .A(n163), .B(r_y_data[19]), .C(r_y_data[51]), .D(n1), .Y(
        n40) );
  scg10d1_hd U703 ( .A(n163), .B(r_y_data[20]), .C(r_y_data[52]), .D(n1), .Y(
        n42) );
  scg10d1_hd U704 ( .A(n163), .B(r_y_data[21]), .C(r_y_data[53]), .D(n1), .Y(
        n44) );
  scg10d1_hd U705 ( .A(n163), .B(r_x_data[39]), .C(r_x_data[71]), .D(n1), .Y(
        n88) );
  scg10d1_hd U706 ( .A(n163), .B(o_Y_DATA[24]), .C(r_y_data[24]), .D(n161), 
        .Y(n51) );
  scg10d1_hd U707 ( .A(n163), .B(r_y_data[22]), .C(r_y_data[54]), .D(n161), 
        .Y(n46) );
  scg10d1_hd U708 ( .A(n163), .B(o_Y_DATA[30]), .C(r_y_data[30]), .D(n161), 
        .Y(n63) );
  scg10d1_hd U709 ( .A(n163), .B(r_y_data[23]), .C(r_y_data[55]), .D(n161), 
        .Y(n48) );
  scg10d1_hd U710 ( .A(n163), .B(r_y_data[24]), .C(r_y_data[56]), .D(n161), 
        .Y(n50) );
  scg10d1_hd U711 ( .A(n163), .B(r_y_data[25]), .C(r_y_data[57]), .D(n161), 
        .Y(n52) );
  scg10d1_hd U712 ( .A(n163), .B(r_y_data[26]), .C(r_y_data[58]), .D(n1), .Y(
        n54) );
  scg10d1_hd U713 ( .A(n163), .B(r_y_data[27]), .C(r_y_data[59]), .D(n161), 
        .Y(n56) );
  scg10d1_hd U714 ( .A(n163), .B(r_y_data[28]), .C(r_y_data[60]), .D(n161), 
        .Y(n58) );
  scg10d1_hd U715 ( .A(n163), .B(r_y_data[29]), .C(r_y_data[61]), .D(n161), 
        .Y(n60) );
  scg10d1_hd U716 ( .A(n163), .B(o_Y_DATA[23]), .C(r_y_data[23]), .D(n161), 
        .Y(n49) );
  scg10d1_hd U717 ( .A(n163), .B(r_y_data[30]), .C(r_y_data[62]), .D(n161), 
        .Y(n62) );
  scg10d1_hd U718 ( .A(n163), .B(r_y_data[6]), .C(r_y_data[38]), .D(n1), .Y(
        n14) );
  scg10d1_hd U719 ( .A(n163), .B(r_x_data[33]), .C(r_x_data[65]), .D(n1), .Y(
        n94) );
  scg10d1_hd U720 ( .A(n163), .B(o_Y_DATA[28]), .C(r_y_data[28]), .D(n161), 
        .Y(n59) );
  scg10d1_hd U721 ( .A(n163), .B(r_x_data[34]), .C(r_x_data[66]), .D(n1), .Y(
        n93) );
  scg10d1_hd U722 ( .A(n163), .B(r_x_data[32]), .C(r_x_data[64]), .D(n1), .Y(
        n95) );
  scg10d1_hd U723 ( .A(n163), .B(o_Y_DATA[27]), .C(r_y_data[27]), .D(n161), 
        .Y(n57) );
  scg10d1_hd U724 ( .A(n163), .B(r_x_data[35]), .C(r_x_data[67]), .D(n1), .Y(
        n92) );
  scg10d1_hd U725 ( .A(n163), .B(r_x_data[36]), .C(r_x_data[68]), .D(n1), .Y(
        n91) );
  scg10d1_hd U726 ( .A(n163), .B(r_y_data[0]), .C(r_y_data[32]), .D(n1), .Y(n2) );
  scg10d1_hd U727 ( .A(n163), .B(r_y_data[1]), .C(r_y_data[33]), .D(n1), .Y(n4) );
  scg10d1_hd U728 ( .A(n163), .B(o_Y_DATA[26]), .C(r_y_data[26]), .D(n161), 
        .Y(n55) );
  scg10d1_hd U729 ( .A(n163), .B(r_y_data[2]), .C(r_y_data[34]), .D(n161), .Y(
        n6) );
  scg10d1_hd U730 ( .A(n163), .B(r_y_data[3]), .C(r_y_data[35]), .D(n161), .Y(
        n8) );
  scg10d1_hd U731 ( .A(n163), .B(r_y_data[4]), .C(r_y_data[36]), .D(n161), .Y(
        n10) );
  scg10d1_hd U732 ( .A(n163), .B(r_y_data[5]), .C(r_y_data[37]), .D(n1), .Y(
        n12) );
  scg10d1_hd U733 ( .A(n163), .B(r_x_data[37]), .C(r_x_data[69]), .D(n1), .Y(
        n90) );
  scg10d1_hd U734 ( .A(n163), .B(r_x_data[40]), .C(r_x_data[72]), .D(n161), 
        .Y(n87) );
  scg10d1_hd U735 ( .A(n163), .B(r_x_data[41]), .C(r_x_data[73]), .D(n161), 
        .Y(n86) );
  scg10d1_hd U736 ( .A(n163), .B(o_Y_DATA[21]), .C(r_y_data[21]), .D(n161), 
        .Y(n45) );
  scg10d1_hd U737 ( .A(n163), .B(o_Y_DATA[20]), .C(r_y_data[20]), .D(n1), .Y(
        n43) );
  scg10d1_hd U738 ( .A(n163), .B(r_x_data[43]), .C(r_x_data[75]), .D(n161), 
        .Y(n84) );
  scg10d1_hd U739 ( .A(n163), .B(o_Y_DATA[22]), .C(r_y_data[22]), .D(n161), 
        .Y(n47) );
  scg10d1_hd U740 ( .A(n163), .B(o_Y_DATA[19]), .C(r_y_data[19]), .D(n1), .Y(
        n41) );
  scg10d1_hd U741 ( .A(n163), .B(o_Y_DATA[18]), .C(r_y_data[18]), .D(n1), .Y(
        n39) );
  scg10d1_hd U742 ( .A(n163), .B(r_x_data[44]), .C(r_x_data[76]), .D(n161), 
        .Y(n83) );
  scg10d1_hd U743 ( .A(n163), .B(o_Y_DATA[17]), .C(r_y_data[17]), .D(n1), .Y(
        n37) );
  scg10d1_hd U744 ( .A(n163), .B(r_x_data[45]), .C(r_x_data[77]), .D(n161), 
        .Y(n82) );
  scg10d1_hd U745 ( .A(n163), .B(r_x_data[42]), .C(r_x_data[74]), .D(n161), 
        .Y(n85) );
  scg10d1_hd U746 ( .A(n163), .B(o_Y_DATA[15]), .C(r_y_data[15]), .D(n1), .Y(
        n33) );
  scg10d1_hd U747 ( .A(n163), .B(o_Y_DATA[16]), .C(r_y_data[16]), .D(n1), .Y(
        n35) );
  scg10d1_hd U748 ( .A(n163), .B(r_x_data[46]), .C(r_x_data[78]), .D(n161), 
        .Y(n81) );
  ivd1_hd U749 ( .A(n641), .Y(n634) );
  nid2_hd U750 ( .A(n716), .Y(n233) );
  ivd1_hd U751 ( .A(n276), .Y(n639) );
  ivd1_hd U752 ( .A(n283), .Y(n632) );
  nid2_hd U753 ( .A(n708), .Y(n230) );
  nr2d1_hd U754 ( .A(n200), .B(n637), .Y(n708) );
  ivd1_hd U755 ( .A(n638), .Y(n285) );
  nr2d1_hd U756 ( .A(n278), .B(n642), .Y(n716) );
  nr2d1_hd U757 ( .A(n278), .B(n277), .Y(n717) );
  ivd1_hd U758 ( .A(n284), .Y(n277) );
  ivd1_hd U759 ( .A(n635), .Y(n633) );
  nr3d1_hd U760 ( .A(n643), .B(n642), .C(n641), .Y(n707) );
  nr2d1_hd U761 ( .A(n708), .B(n640), .Y(n643) );
  oa211d1_hd U762 ( .A(n285), .B(n283), .C(n284), .D(n282), .Y(n705) );
  oa211d1_hd U763 ( .A(n284), .B(n632), .C(n275), .D(n282), .Y(n714) );
  nr2d1_hd U764 ( .A(n632), .B(n270), .Y(n276) );
  nr2d1_hd U765 ( .A(n811), .B(n816), .Y(n284) );
  nr2d1_hd U766 ( .A(n199), .B(n580), .Y(n283) );
  nd4d1_hd U767 ( .A(n634), .B(w_add_Z_STB), .C(w_mult_2_Z_STB), .D(
        w_mult_1_Z_STB), .Y(n638) );
  ivd1_hd U768 ( .A(n281), .Y(n272) );
  scg6d1_hd U769 ( .A(r_mult_1_A[14]), .B(n169), .C(n715), .Y(n424) );
  scg6d1_hd U770 ( .A(r_mult_1_A[15]), .B(n169), .C(n715), .Y(n423) );
  scg6d1_hd U771 ( .A(r_mult_1_A[25]), .B(n169), .C(n715), .Y(n415) );
  scg6d1_hd U772 ( .A(r_mult_2_A[4]), .B(n169), .C(n715), .Y(n406) );
  scg6d1_hd U773 ( .A(r_mult_1_A[24]), .B(n169), .C(n715), .Y(n416) );
  scg6d1_hd U774 ( .A(r_mult_2_A[8]), .B(n169), .C(n715), .Y(n402) );
  scg6d1_hd U775 ( .A(r_mult_1_A[12]), .B(n169), .C(n715), .Y(n425) );
  scg6d1_hd U776 ( .A(r_mult_1_A[9]), .B(n169), .C(n715), .Y(n428) );
  scg6d1_hd U777 ( .A(r_mult_2_A[13]), .B(n169), .C(n715), .Y(n399) );
  scg6d1_hd U778 ( .A(r_mult_2_A[14]), .B(n169), .C(n715), .Y(n398) );
  scg6d1_hd U779 ( .A(r_mult_2_A[24]), .B(n169), .C(n715), .Y(n391) );
  scg6d1_hd U780 ( .A(r_mult_2_A[21]), .B(n169), .C(n715), .Y(n393) );
  scg6d1_hd U781 ( .A(r_mult_2_A[31]), .B(n169), .C(n232), .Y(n385) );
  scg6d1_hd U782 ( .A(r_mult_2_A[25]), .B(n169), .C(n232), .Y(n390) );
  scg6d1_hd U783 ( .A(r_mult_1_A[4]), .B(n169), .C(n232), .Y(n433) );
  scg6d1_hd U784 ( .A(r_mult_1_A[8]), .B(n169), .C(n232), .Y(n429) );
  scg14d1_hd U785 ( .A(w_add_Z[27]), .B(n350), .C(n291), .Y(n442) );
  scg14d1_hd U786 ( .A(w_add_Z[26]), .B(n350), .C(n292), .Y(n443) );
  scg14d1_hd U787 ( .A(w_add_Z[28]), .B(n350), .C(n290), .Y(n441) );
  scg14d1_hd U788 ( .A(w_add_Z[25]), .B(n350), .C(n293), .Y(n444) );
  scg14d1_hd U789 ( .A(w_add_Z[23]), .B(n350), .C(n295), .Y(n446) );
  scg14d1_hd U790 ( .A(w_add_Z[24]), .B(n350), .C(n294), .Y(n445) );
  ao21d1_hd U791 ( .A(n639), .B(n638), .C(n642), .Y(n640) );
  scg14d1_hd U792 ( .A(r_mult_2_A[22]), .B(n169), .C(n167), .Y(n392) );
  scg14d1_hd U793 ( .A(r_mult_1_A[0]), .B(n169), .C(n167), .Y(n437) );
  scg14d1_hd U794 ( .A(r_mult_2_A[2]), .B(n169), .C(n167), .Y(n408) );
  scg14d1_hd U795 ( .A(r_mult_1_A[2]), .B(n169), .C(n167), .Y(n435) );
  scg14d1_hd U796 ( .A(r_mult_1_A[1]), .B(n169), .C(n167), .Y(n436) );
  scg14d1_hd U797 ( .A(r_mult_2_A[19]), .B(n169), .C(n167), .Y(n395) );
  scg14d1_hd U798 ( .A(r_mult_2_A[1]), .B(n169), .C(n167), .Y(n409) );
  scg4d1_hd U799 ( .A(n279), .B(w_add_Z[17]), .C(n231), .D(r_add_B[17]), .E(
        r_x_data[81]), .F(n715), .G(n234), .H(w_mult_2_Z[17]), .Y(n366) );
  scg4d1_hd U800 ( .A(n279), .B(w_add_Z[19]), .C(n231), .D(r_add_B[19]), .E(
        r_x_data[83]), .F(n715), .G(n234), .H(w_mult_2_Z[19]), .Y(n364) );
  scg4d1_hd U801 ( .A(n279), .B(w_add_Z[13]), .C(n231), .D(r_add_B[13]), .E(
        r_x_data[77]), .F(n715), .G(n234), .H(w_mult_2_Z[13]), .Y(n370) );
  scg14d1_hd U802 ( .A(w_add_Z[22]), .B(n350), .C(n296), .Y(n447) );
  scg14d1_hd U803 ( .A(w_add_Z[19]), .B(n350), .C(n299), .Y(n450) );
  scg14d1_hd U804 ( .A(w_add_Z[21]), .B(n350), .C(n297), .Y(n448) );
  scg14d1_hd U805 ( .A(w_add_Z[13]), .B(n350), .C(n305), .Y(n456) );
  scg14d1_hd U806 ( .A(w_add_Z[17]), .B(n350), .C(n301), .Y(n452) );
  scg14d1_hd U807 ( .A(w_add_Z[15]), .B(n350), .C(n303), .Y(n454) );
  scg14d1_hd U808 ( .A(w_add_Z[20]), .B(n350), .C(n298), .Y(n449) );
  scg14d1_hd U809 ( .A(w_add_Z[16]), .B(n350), .C(n302), .Y(n453) );
  scg14d1_hd U810 ( .A(w_add_Z[12]), .B(n350), .C(n306), .Y(n457) );
  scg14d1_hd U811 ( .A(w_add_Z[14]), .B(n350), .C(n304), .Y(n455) );
  scg14d1_hd U812 ( .A(w_add_Z[18]), .B(n350), .C(n300), .Y(n451) );
  ivd1_hd U813 ( .A(o_Y_DATA[6]), .Y(n693) );
  ivd1_hd U814 ( .A(o_Y_DATA[4]), .Y(n697) );
  ivd1_hd U815 ( .A(o_Y_DATA[5]), .Y(n695) );
  ivd1_hd U816 ( .A(o_Y_DATA[2]), .Y(n701) );
  ivd1_hd U817 ( .A(o_Y_DATA[7]), .Y(n691) );
  ivd1_hd U818 ( .A(o_Y_DATA[8]), .Y(n689) );
  ivd1_hd U819 ( .A(o_Y_DATA[3]), .Y(n699) );
  ivd1_hd U820 ( .A(o_Y_DATA[1]), .Y(n703) );
  ivd1_hd U821 ( .A(o_Y_DATA[20]), .Y(n665) );
  scg14d1_hd U822 ( .A(n350), .B(r_x_data[61]), .C(n320), .Y(n471) );
  scg14d1_hd U823 ( .A(n350), .B(r_x_data[62]), .C(n319), .Y(n470) );
  scg14d1_hd U824 ( .A(n350), .B(r_x_data[60]), .C(n321), .Y(n472) );
  scg4d1_hd U825 ( .A(n279), .B(w_add_Z[11]), .C(n231), .D(r_add_B[11]), .E(
        r_x_data[75]), .F(n715), .G(n234), .H(w_mult_2_Z[11]), .Y(n372) );
  scg4d1_hd U826 ( .A(n279), .B(w_add_Z[26]), .C(n231), .D(r_add_B[26]), .E(
        r_x_data[90]), .F(n715), .G(n234), .H(w_mult_2_Z[26]), .Y(n357) );
  scg4d1_hd U827 ( .A(n279), .B(w_add_Z[28]), .C(n231), .D(r_add_B[28]), .E(
        r_x_data[92]), .F(n715), .G(n234), .H(w_mult_2_Z[28]), .Y(n355) );
  scg4d1_hd U828 ( .A(n279), .B(w_add_Z[22]), .C(n231), .D(r_add_B[22]), .E(
        r_x_data[86]), .F(n715), .G(n234), .H(w_mult_2_Z[22]), .Y(n361) );
  scg4d1_hd U829 ( .A(n279), .B(w_add_Z[12]), .C(n231), .D(r_add_B[12]), .E(
        r_x_data[76]), .F(n715), .G(n234), .H(w_mult_2_Z[12]), .Y(n371) );
  scg4d1_hd U830 ( .A(n279), .B(w_add_Z[24]), .C(n231), .D(r_add_B[24]), .E(
        r_x_data[88]), .F(n715), .G(n234), .H(w_mult_2_Z[24]), .Y(n359) );
  ivd1_hd U831 ( .A(o_Y_DATA[31]), .Y(n713) );
  ivd1_hd U832 ( .A(o_Y_DATA[26]), .Y(n653) );
  ivd1_hd U833 ( .A(o_Y_DATA[23]), .Y(n659) );
  ivd1_hd U834 ( .A(o_Y_DATA[22]), .Y(n661) );
  ivd1_hd U835 ( .A(o_Y_DATA[25]), .Y(n655) );
  ivd1_hd U836 ( .A(o_Y_DATA[28]), .Y(n649) );
  ivd1_hd U837 ( .A(o_Y_DATA[29]), .Y(n647) );
  ivd1_hd U838 ( .A(o_Y_DATA[21]), .Y(n663) );
  ivd1_hd U839 ( .A(o_Y_DATA[27]), .Y(n651) );
  ivd1_hd U840 ( .A(o_Y_DATA[24]), .Y(n657) );
  scg14d1_hd U841 ( .A(w_add_Z[11]), .B(n350), .C(n307), .Y(n458) );
  ivd1_hd U842 ( .A(o_Y_DATA[0]), .Y(n720) );
  ivd1_hd U843 ( .A(o_Y_DATA[9]), .Y(n687) );
  ivd1_hd U844 ( .A(o_Y_DATA[19]), .Y(n667) );
  ivd1_hd U845 ( .A(o_Y_DATA[16]), .Y(n673) );
  ivd1_hd U846 ( .A(o_Y_DATA[30]), .Y(n645) );
  ivd1_hd U847 ( .A(o_Y_DATA[14]), .Y(n677) );
  ivd1_hd U848 ( .A(o_Y_DATA[13]), .Y(n679) );
  ivd1_hd U849 ( .A(o_Y_DATA[15]), .Y(n675) );
  ivd1_hd U850 ( .A(o_Y_DATA[17]), .Y(n671) );
  ivd1_hd U851 ( .A(o_Y_DATA[18]), .Y(n669) );
  ivd1_hd U852 ( .A(o_Y_DATA[10]), .Y(n685) );
  ivd1_hd U853 ( .A(o_Y_DATA[12]), .Y(n681) );
  nd3d1_hd U854 ( .A(w_mult_2_AB_ACK), .B(w_add_AB_ACK), .C(w_mult_1_AB_ACK), 
        .Y(n270) );
  ivd1_hd U855 ( .A(o_Y_DATA[11]), .Y(n683) );
  oa21d1_hd U856 ( .A(n637), .B(n811), .C(n633), .Y(n275) );
  nr2d1_hd U857 ( .A(n641), .B(n170), .Y(n274) );
  nr2d1_hd U858 ( .A(n1195), .B(n580), .Y(n273) );
  nd2bd1_hd U859 ( .AN(r_mult_1_A[29]), .B(n286), .Y(n411) );
  nd2bd1_hd U860 ( .AN(r_mult_1_A[27]), .B(n286), .Y(n413) );
  nd2bd1_hd U861 ( .AN(r_mult_2_A[0]), .B(n286), .Y(n410) );
  nd2bd1_hd U862 ( .AN(r_mult_1_A[26]), .B(n286), .Y(n414) );
  nd2bd1_hd U863 ( .AN(r_mult_1_A[28]), .B(n286), .Y(n412) );
  nd2bd1_hd U864 ( .AN(r_mult_2_A[17]), .B(n286), .Y(n396) );
  nd2bd1_hd U865 ( .AN(r_mult_2_A[28]), .B(n286), .Y(n387) );
  nd2bd1_hd U866 ( .AN(r_mult_2_A[20]), .B(n286), .Y(n394) );
  nd2bd1_hd U867 ( .AN(r_mult_2_A[6]), .B(n286), .Y(n404) );
  nd2bd1_hd U868 ( .AN(r_mult_2_A[16]), .B(n286), .Y(n397) );
  nd2bd1_hd U869 ( .AN(r_mult_2_A[11]), .B(n286), .Y(n400) );
  nd2bd1_hd U870 ( .AN(r_mult_2_A[10]), .B(n286), .Y(n401) );
  nd2bd1_hd U871 ( .AN(r_mult_2_A[7]), .B(n286), .Y(n403) );
  nd2bd1_hd U872 ( .AN(r_mult_1_A[3]), .B(n286), .Y(n434) );
  nd2bd1_hd U873 ( .AN(r_mult_2_A[27]), .B(n286), .Y(n388) );
  nd2bd1_hd U874 ( .AN(r_mult_1_A[22]), .B(n286), .Y(n418) );
  nd2bd1_hd U875 ( .AN(r_mult_2_A[29]), .B(n286), .Y(n386) );
  nd2bd1_hd U876 ( .AN(r_mult_1_A[20]), .B(n286), .Y(n419) );
  nd2bd1_hd U877 ( .AN(r_mult_1_A[17]), .B(n286), .Y(n421) );
  nd2bd1_hd U878 ( .AN(r_mult_2_A[26]), .B(n286), .Y(n389) );
  nd2bd1_hd U879 ( .AN(r_mult_1_A[7]), .B(n286), .Y(n430) );
  oa21d1_hd U880 ( .A(n816), .B(n638), .C(n632), .Y(n635) );
  nd2bd1_hd U881 ( .AN(r_mult_1_A[23]), .B(n286), .Y(n417) );
  nd2bd1_hd U882 ( .AN(r_mult_1_A[10]), .B(n286), .Y(n427) );
  nd2bd1_hd U883 ( .AN(r_mult_2_A[3]), .B(n286), .Y(n407) );
  nd2bd1_hd U884 ( .AN(r_mult_2_A[5]), .B(n286), .Y(n405) );
  nd2bd1_hd U885 ( .AN(r_mult_1_A[6]), .B(n286), .Y(n431) );
  nd2bd1_hd U886 ( .AN(r_mult_1_A[5]), .B(n286), .Y(n432) );
  nd2bd1_hd U887 ( .AN(r_mult_1_A[11]), .B(n286), .Y(n426) );
  nr2bd1_hd U888 ( .AN(n273), .B(N18), .Y(N814) );
  ao22d1_hd U889 ( .A(n235), .B(n201), .C(n171), .D(n163), .Y(n100) );
  ao22d1_hd U890 ( .A(n235), .B(n202), .C(n172), .D(n572), .Y(n101) );
  ao22d1_hd U891 ( .A(n235), .B(n203), .C(n173), .D(n572), .Y(n102) );
  ao22d1_hd U892 ( .A(n235), .B(n204), .C(n174), .D(n163), .Y(n103) );
  ao22d1_hd U893 ( .A(n235), .B(n205), .C(n175), .D(n163), .Y(n104) );
  ao22d1_hd U894 ( .A(n235), .B(n206), .C(n176), .D(n163), .Y(n105) );
  ao22d1_hd U895 ( .A(n235), .B(n207), .C(n177), .D(n163), .Y(n106) );
  ao22d1_hd U896 ( .A(n235), .B(n208), .C(n178), .D(n163), .Y(n107) );
  ao22d1_hd U897 ( .A(n235), .B(n209), .C(n179), .D(n163), .Y(n108) );
  ao22d1_hd U898 ( .A(n235), .B(n210), .C(n180), .D(n572), .Y(n109) );
  ao22d1_hd U899 ( .A(n235), .B(n211), .C(n181), .D(n572), .Y(n110) );
  ao22d1_hd U900 ( .A(n235), .B(n212), .C(n182), .D(n572), .Y(n111) );
  ao22d1_hd U901 ( .A(n235), .B(n213), .C(n183), .D(n572), .Y(n112) );
  ao22d1_hd U902 ( .A(n235), .B(n214), .C(n184), .D(n572), .Y(n113) );
  ao22d1_hd U903 ( .A(n235), .B(n215), .C(n185), .D(n572), .Y(n114) );
  ao22d1_hd U904 ( .A(n235), .B(n216), .C(n186), .D(n572), .Y(n115) );
  ao22d1_hd U905 ( .A(n235), .B(n217), .C(n187), .D(n572), .Y(n116) );
  ao22d1_hd U906 ( .A(n235), .B(n218), .C(n188), .D(n572), .Y(n117) );
  ao22d1_hd U907 ( .A(n235), .B(n219), .C(n189), .D(n572), .Y(n118) );
  ao22d1_hd U908 ( .A(n235), .B(n220), .C(n190), .D(n572), .Y(n119) );
  ao22d1_hd U909 ( .A(n235), .B(n221), .C(n191), .D(n572), .Y(n120) );
  ao22d1_hd U910 ( .A(n235), .B(n222), .C(n192), .D(n572), .Y(n121) );
  ao22d1_hd U911 ( .A(n235), .B(n223), .C(n193), .D(n572), .Y(n122) );
  ao22d1_hd U912 ( .A(n235), .B(n224), .C(n194), .D(n572), .Y(n123) );
  ao22d1_hd U913 ( .A(n235), .B(n225), .C(n195), .D(n572), .Y(n124) );
  ao22d1_hd U914 ( .A(n235), .B(n226), .C(n196), .D(n572), .Y(n125) );
  ao22d1_hd U915 ( .A(n235), .B(n227), .C(n197), .D(n572), .Y(n126) );
  ao22d1_hd U916 ( .A(n235), .B(n228), .C(n198), .D(n572), .Y(n127) );
  oa21d1_hd U917 ( .A(n201), .B(n1), .C(n236), .Y(n132) );
  oa21d1_hd U918 ( .A(n202), .B(n1), .C(n237), .Y(n133) );
  oa21d1_hd U919 ( .A(n203), .B(n1), .C(n238), .Y(n134) );
  oa21d1_hd U920 ( .A(n204), .B(n1), .C(n239), .Y(n135) );
  oa21d1_hd U921 ( .A(n205), .B(n1), .C(n240), .Y(n136) );
  oa21d1_hd U922 ( .A(n206), .B(n1), .C(n241), .Y(n137) );
  oa21d1_hd U923 ( .A(n207), .B(n1), .C(n242), .Y(n138) );
  oa21d1_hd U924 ( .A(n208), .B(n1), .C(n243), .Y(n139) );
  oa21d1_hd U925 ( .A(n209), .B(n1), .C(n244), .Y(n140) );
  oa21d1_hd U926 ( .A(n210), .B(n1), .C(n245), .Y(n141) );
  oa21d1_hd U927 ( .A(n211), .B(n1), .C(n246), .Y(n142) );
  oa21d1_hd U928 ( .A(n212), .B(n1), .C(n247), .Y(n143) );
  oa21d1_hd U929 ( .A(n213), .B(n1), .C(n248), .Y(n144) );
  oa21d1_hd U930 ( .A(n214), .B(n1), .C(n249), .Y(n145) );
  oa21d1_hd U931 ( .A(n215), .B(n1), .C(n250), .Y(n146) );
  oa21d1_hd U932 ( .A(n216), .B(n1), .C(n251), .Y(n147) );
  oa21d1_hd U933 ( .A(n217), .B(n1), .C(n252), .Y(n148) );
  oa21d1_hd U934 ( .A(n218), .B(n235), .C(n253), .Y(n149) );
  oa21d1_hd U935 ( .A(n219), .B(n235), .C(n254), .Y(n150) );
  oa21d1_hd U936 ( .A(n220), .B(n235), .C(n255), .Y(n151) );
  oa21d1_hd U937 ( .A(n221), .B(n235), .C(n256), .Y(n152) );
  oa21d1_hd U938 ( .A(n222), .B(n235), .C(n257), .Y(n153) );
  oa21d1_hd U939 ( .A(n223), .B(n1), .C(n258), .Y(n154) );
  oa21d1_hd U940 ( .A(n224), .B(n1), .C(n259), .Y(n155) );
  oa21d1_hd U941 ( .A(n225), .B(n1), .C(n260), .Y(n156) );
  oa21d1_hd U942 ( .A(n226), .B(n1), .C(n261), .Y(n157) );
  oa21d1_hd U943 ( .A(n227), .B(n1), .C(n262), .Y(n158) );
  oa21d1_hd U944 ( .A(n228), .B(n1), .C(n263), .Y(n159) );
  nr2d1_hd U945 ( .A(n200), .B(n170), .Y(n266) );
  scg17d1_hd U946 ( .A(n170), .B(n264), .C(n266), .D(w_add_Z_STB), .Y(n265) );
  scg15d1_hd U947 ( .A(o_Y_DATA_VALID), .B(i_Y_ACK), .C(n1195), .D(n580), .Y(
        n281) );
  ao211d1_hd U948 ( .A(n634), .B(n265), .C(n272), .D(n276), .Y(n160) );
  nr2d1_hd U949 ( .A(n273), .B(n631), .Y(n268) );
  ao22d1_hd U950 ( .A(n811), .B(n268), .C(n631), .D(n200), .Y(n162) );
  nr2d1_hd U951 ( .A(n268), .B(n200), .Y(n269) );
  nr2d1_hd U952 ( .A(n266), .B(n641), .Y(n267) );
  oa22d1_hd U953 ( .A(n816), .B(n269), .C(n268), .D(n267), .Y(n166) );
  nd2bd1_hd U954 ( .AN(n631), .B(n282), .Y(n271) );
  ao211d1_hd U955 ( .A(n273), .B(n1), .C(n272), .D(n271), .Y(n168) );
  scg4d1_hd U956 ( .A(n279), .B(w_add_Z[31]), .C(n231), .D(r_add_B[31]), .E(
        r_x_data[95]), .F(n715), .G(n234), .H(w_mult_2_Z[31]), .Y(n352) );
  scg4d1_hd U957 ( .A(n279), .B(w_add_Z[30]), .C(n231), .D(r_add_B[30]), .E(
        r_x_data[94]), .F(n715), .G(n234), .H(w_mult_2_Z[30]), .Y(n353) );
  scg4d1_hd U958 ( .A(n279), .B(w_add_Z[29]), .C(n231), .D(r_add_B[29]), .E(
        r_x_data[93]), .F(n715), .G(n234), .H(w_mult_2_Z[29]), .Y(n354) );
  scg4d1_hd U959 ( .A(n279), .B(w_add_Z[27]), .C(n231), .D(r_add_B[27]), .E(
        r_x_data[91]), .F(n715), .G(n234), .H(w_mult_2_Z[27]), .Y(n356) );
  scg4d1_hd U960 ( .A(n279), .B(w_add_Z[25]), .C(n231), .D(r_add_B[25]), .E(
        r_x_data[89]), .F(n715), .G(n234), .H(w_mult_2_Z[25]), .Y(n358) );
  scg4d1_hd U961 ( .A(n279), .B(w_add_Z[23]), .C(n231), .D(r_add_B[23]), .E(
        r_x_data[87]), .F(n715), .G(n234), .H(w_mult_2_Z[23]), .Y(n360) );
  scg4d1_hd U962 ( .A(n279), .B(w_add_Z[21]), .C(n231), .D(r_add_B[21]), .E(
        r_x_data[85]), .F(n715), .G(n234), .H(w_mult_2_Z[21]), .Y(n362) );
  scg4d1_hd U963 ( .A(n279), .B(w_add_Z[20]), .C(n231), .D(r_add_B[20]), .E(
        r_x_data[84]), .F(n715), .G(n234), .H(w_mult_2_Z[20]), .Y(n363) );
  scg4d1_hd U964 ( .A(n279), .B(w_add_Z[18]), .C(n231), .D(r_add_B[18]), .E(
        r_x_data[82]), .F(n715), .G(n234), .H(w_mult_2_Z[18]), .Y(n365) );
  scg4d1_hd U965 ( .A(n279), .B(w_add_Z[16]), .C(n231), .D(r_add_B[16]), .E(
        r_x_data[80]), .F(n715), .G(n234), .H(w_mult_2_Z[16]), .Y(n367) );
  scg4d1_hd U966 ( .A(n279), .B(w_add_Z[15]), .C(n714), .D(r_add_B[15]), .E(
        r_x_data[79]), .F(n715), .G(n234), .H(w_mult_2_Z[15]), .Y(n368) );
  scg4d1_hd U967 ( .A(n279), .B(w_add_Z[14]), .C(n714), .D(r_add_B[14]), .E(
        r_x_data[78]), .F(n715), .G(n234), .H(w_mult_2_Z[14]), .Y(n369) );
  scg4d1_hd U968 ( .A(n279), .B(w_add_Z[10]), .C(n231), .D(r_add_B[10]), .E(
        r_x_data[74]), .F(n715), .G(n234), .H(w_mult_2_Z[10]), .Y(n373) );
  scg4d1_hd U969 ( .A(n279), .B(w_add_Z[9]), .C(n231), .D(r_add_B[9]), .E(
        r_x_data[73]), .F(n715), .G(n234), .H(w_mult_2_Z[9]), .Y(n374) );
  scg4d1_hd U970 ( .A(n279), .B(w_add_Z[8]), .C(n231), .D(r_add_B[8]), .E(
        r_x_data[72]), .F(n715), .G(n234), .H(w_mult_2_Z[8]), .Y(n375) );
  scg4d1_hd U971 ( .A(n279), .B(w_add_Z[7]), .C(n231), .D(r_add_B[7]), .E(
        r_x_data[71]), .F(n715), .G(n234), .H(w_mult_2_Z[7]), .Y(n376) );
  scg4d1_hd U972 ( .A(n279), .B(w_add_Z[6]), .C(n231), .D(r_add_B[6]), .E(
        r_x_data[70]), .F(n715), .G(n234), .H(w_mult_2_Z[6]), .Y(n377) );
  scg4d1_hd U973 ( .A(n279), .B(w_add_Z[5]), .C(n231), .D(r_add_B[5]), .E(
        r_x_data[69]), .F(n715), .G(n234), .H(w_mult_2_Z[5]), .Y(n378) );
  scg4d1_hd U974 ( .A(n279), .B(w_add_Z[4]), .C(n231), .D(r_add_B[4]), .E(
        r_x_data[68]), .F(n715), .G(n234), .H(w_mult_2_Z[4]), .Y(n379) );
  scg4d1_hd U975 ( .A(n279), .B(w_add_Z[3]), .C(n231), .D(r_add_B[3]), .E(
        r_x_data[67]), .F(n715), .G(n234), .H(w_mult_2_Z[3]), .Y(n380) );
  scg4d1_hd U976 ( .A(n279), .B(w_add_Z[2]), .C(n231), .D(r_add_B[2]), .E(
        r_x_data[66]), .F(n715), .G(n234), .H(w_mult_2_Z[2]), .Y(n381) );
  scg4d1_hd U977 ( .A(n279), .B(w_add_Z[1]), .C(n231), .D(r_add_B[1]), .E(
        r_x_data[65]), .F(n715), .G(n234), .H(w_mult_2_Z[1]), .Y(n382) );
  scg4d1_hd U978 ( .A(n279), .B(w_add_Z[0]), .C(n231), .D(r_add_B[0]), .E(
        r_x_data[64]), .F(n715), .G(n234), .H(w_mult_2_Z[0]), .Y(n383) );
  oa21d1_hd U979 ( .A(n283), .B(n634), .C(o_Y_DATA_VALID), .Y(n280) );
  scg14d1_hd U980 ( .A(r_mult_1_A[19]), .B(n705), .C(n167), .Y(n420) );
  scg14d1_hd U981 ( .A(r_mult_1_A[16]), .B(n705), .C(n167), .Y(n422) );
  oa22d1_hd U982 ( .A(n634), .B(n287), .C(n816), .D(n639), .Y(n438) );
  ao22d1_hd U983 ( .A(n232), .B(r_y_data[62]), .C(r_mult_2_B[30]), .D(n169), 
        .Y(n288) );
  scg14d1_hd U984 ( .A(w_add_Z[30]), .B(n350), .C(n288), .Y(n439) );
  ao22d1_hd U985 ( .A(n232), .B(r_y_data[61]), .C(r_mult_2_B[29]), .D(n169), 
        .Y(n289) );
  scg14d1_hd U986 ( .A(w_add_Z[29]), .B(n350), .C(n289), .Y(n440) );
  ao22d1_hd U987 ( .A(n232), .B(r_y_data[60]), .C(r_mult_2_B[28]), .D(n169), 
        .Y(n290) );
  ao22d1_hd U988 ( .A(n232), .B(r_y_data[59]), .C(r_mult_2_B[27]), .D(n169), 
        .Y(n291) );
  ao22d1_hd U989 ( .A(n232), .B(r_y_data[58]), .C(r_mult_2_B[26]), .D(n169), 
        .Y(n292) );
  ao22d1_hd U990 ( .A(n232), .B(r_y_data[57]), .C(r_mult_2_B[25]), .D(n169), 
        .Y(n293) );
  ao22d1_hd U991 ( .A(n232), .B(r_y_data[56]), .C(r_mult_2_B[24]), .D(n169), 
        .Y(n294) );
  ao22d1_hd U992 ( .A(n232), .B(r_y_data[55]), .C(r_mult_2_B[23]), .D(n169), 
        .Y(n295) );
  ao22d1_hd U993 ( .A(n232), .B(r_y_data[54]), .C(r_mult_2_B[22]), .D(n169), 
        .Y(n296) );
  ao22d1_hd U994 ( .A(n232), .B(r_y_data[53]), .C(r_mult_2_B[21]), .D(n169), 
        .Y(n297) );
  ao22d1_hd U995 ( .A(n232), .B(r_y_data[52]), .C(r_mult_2_B[20]), .D(n169), 
        .Y(n298) );
  ao22d1_hd U996 ( .A(n232), .B(r_y_data[51]), .C(r_mult_2_B[19]), .D(n169), 
        .Y(n299) );
  ao22d1_hd U997 ( .A(n232), .B(r_y_data[50]), .C(r_mult_2_B[18]), .D(n169), 
        .Y(n300) );
  ao22d1_hd U998 ( .A(n232), .B(r_y_data[49]), .C(r_mult_2_B[17]), .D(n169), 
        .Y(n301) );
  ao22d1_hd U999 ( .A(n232), .B(r_y_data[48]), .C(r_mult_2_B[16]), .D(n169), 
        .Y(n302) );
  ao22d1_hd U1000 ( .A(n232), .B(r_y_data[47]), .C(r_mult_2_B[15]), .D(n169), 
        .Y(n303) );
  ao22d1_hd U1001 ( .A(n232), .B(r_y_data[46]), .C(r_mult_2_B[14]), .D(n169), 
        .Y(n304) );
  ao22d1_hd U1002 ( .A(n232), .B(r_y_data[45]), .C(r_mult_2_B[13]), .D(n169), 
        .Y(n305) );
  ao22d1_hd U1003 ( .A(n232), .B(r_y_data[44]), .C(r_mult_2_B[12]), .D(n169), 
        .Y(n306) );
  ao22d1_hd U1004 ( .A(n232), .B(r_y_data[43]), .C(r_mult_2_B[11]), .D(n705), 
        .Y(n307) );
  ao22d1_hd U1005 ( .A(n232), .B(r_y_data[42]), .C(r_mult_2_B[10]), .D(n169), 
        .Y(n308) );
  scg14d1_hd U1006 ( .A(w_add_Z[10]), .B(n350), .C(n308), .Y(n459) );
  ao22d1_hd U1007 ( .A(n232), .B(r_y_data[41]), .C(r_mult_2_B[9]), .D(n169), 
        .Y(n309) );
  scg14d1_hd U1008 ( .A(w_add_Z[9]), .B(n350), .C(n309), .Y(n460) );
  ao22d1_hd U1009 ( .A(n232), .B(r_y_data[40]), .C(r_mult_2_B[8]), .D(n169), 
        .Y(n310) );
  scg14d1_hd U1010 ( .A(w_add_Z[8]), .B(n350), .C(n310), .Y(n461) );
  ao22d1_hd U1011 ( .A(n232), .B(r_y_data[39]), .C(r_mult_2_B[7]), .D(n169), 
        .Y(n311) );
  scg14d1_hd U1012 ( .A(w_add_Z[7]), .B(n350), .C(n311), .Y(n462) );
  ao22d1_hd U1013 ( .A(n232), .B(r_y_data[38]), .C(r_mult_2_B[6]), .D(n169), 
        .Y(n312) );
  scg14d1_hd U1014 ( .A(w_add_Z[6]), .B(n350), .C(n312), .Y(n463) );
  ao22d1_hd U1015 ( .A(n232), .B(r_y_data[37]), .C(r_mult_2_B[5]), .D(n169), 
        .Y(n313) );
  scg14d1_hd U1016 ( .A(w_add_Z[5]), .B(n350), .C(n313), .Y(n464) );
  ao22d1_hd U1017 ( .A(n232), .B(r_y_data[36]), .C(r_mult_2_B[4]), .D(n169), 
        .Y(n314) );
  scg14d1_hd U1018 ( .A(w_add_Z[4]), .B(n350), .C(n314), .Y(n465) );
  ao22d1_hd U1019 ( .A(n232), .B(r_y_data[35]), .C(r_mult_2_B[3]), .D(n169), 
        .Y(n315) );
  scg14d1_hd U1020 ( .A(w_add_Z[3]), .B(n350), .C(n315), .Y(n466) );
  ao22d1_hd U1021 ( .A(n232), .B(r_y_data[34]), .C(r_mult_2_B[2]), .D(n169), 
        .Y(n316) );
  scg14d1_hd U1022 ( .A(w_add_Z[2]), .B(n350), .C(n316), .Y(n467) );
  ao22d1_hd U1023 ( .A(n232), .B(r_y_data[33]), .C(r_mult_2_B[1]), .D(n169), 
        .Y(n317) );
  scg14d1_hd U1024 ( .A(w_add_Z[1]), .B(n350), .C(n317), .Y(n468) );
  ao22d1_hd U1025 ( .A(n232), .B(r_y_data[32]), .C(r_mult_2_B[0]), .D(n169), 
        .Y(n318) );
  scg14d1_hd U1026 ( .A(w_add_Z[0]), .B(n350), .C(n318), .Y(n469) );
  ao22d1_hd U1027 ( .A(n232), .B(r_y_data[30]), .C(r_mult_1_B[30]), .D(n169), 
        .Y(n319) );
  ao22d1_hd U1028 ( .A(n232), .B(r_y_data[29]), .C(r_mult_1_B[29]), .D(n169), 
        .Y(n320) );
  ao22d1_hd U1029 ( .A(n232), .B(r_y_data[28]), .C(r_mult_1_B[28]), .D(n169), 
        .Y(n321) );
  ao22d1_hd U1030 ( .A(n232), .B(r_y_data[27]), .C(r_mult_1_B[27]), .D(n169), 
        .Y(n322) );
  oa21d1_hd U1031 ( .A(n167), .B(n171), .C(n322), .Y(n473) );
  ao22d1_hd U1032 ( .A(n232), .B(r_y_data[26]), .C(r_mult_1_B[26]), .D(n169), 
        .Y(n323) );
  oa21d1_hd U1033 ( .A(n167), .B(n172), .C(n323), .Y(n474) );
  ao22d1_hd U1034 ( .A(n232), .B(r_y_data[25]), .C(r_mult_1_B[25]), .D(n169), 
        .Y(n324) );
  oa21d1_hd U1035 ( .A(n167), .B(n173), .C(n324), .Y(n475) );
  ao22d1_hd U1036 ( .A(n232), .B(r_y_data[24]), .C(r_mult_1_B[24]), .D(n169), 
        .Y(n325) );
  oa21d1_hd U1037 ( .A(n167), .B(n174), .C(n325), .Y(n476) );
  ao22d1_hd U1038 ( .A(n232), .B(r_y_data[23]), .C(r_mult_1_B[23]), .D(n169), 
        .Y(n326) );
  oa21d1_hd U1039 ( .A(n167), .B(n175), .C(n326), .Y(n477) );
  ao22d1_hd U1040 ( .A(n232), .B(r_y_data[22]), .C(r_mult_1_B[22]), .D(n169), 
        .Y(n327) );
  oa21d1_hd U1041 ( .A(n167), .B(n176), .C(n327), .Y(n478) );
  ao22d1_hd U1042 ( .A(n232), .B(r_y_data[21]), .C(r_mult_1_B[21]), .D(n169), 
        .Y(n328) );
  oa21d1_hd U1043 ( .A(n167), .B(n177), .C(n328), .Y(n479) );
  ao22d1_hd U1044 ( .A(n232), .B(r_y_data[20]), .C(r_mult_1_B[20]), .D(n169), 
        .Y(n329) );
  oa21d1_hd U1045 ( .A(n167), .B(n178), .C(n329), .Y(n480) );
  ao22d1_hd U1046 ( .A(n232), .B(r_y_data[19]), .C(r_mult_1_B[19]), .D(n169), 
        .Y(n330) );
  oa21d1_hd U1047 ( .A(n167), .B(n179), .C(n330), .Y(n481) );
  ao22d1_hd U1048 ( .A(n232), .B(r_y_data[18]), .C(r_mult_1_B[18]), .D(n169), 
        .Y(n331) );
  oa21d1_hd U1049 ( .A(n167), .B(n180), .C(n331), .Y(n482) );
  ao22d1_hd U1050 ( .A(n232), .B(r_y_data[17]), .C(r_mult_1_B[17]), .D(n169), 
        .Y(n332) );
  oa21d1_hd U1051 ( .A(n167), .B(n181), .C(n332), .Y(n483) );
  ao22d1_hd U1052 ( .A(n232), .B(r_y_data[16]), .C(r_mult_1_B[16]), .D(n169), 
        .Y(n333) );
  oa21d1_hd U1053 ( .A(n167), .B(n182), .C(n333), .Y(n484) );
  ao22d1_hd U1054 ( .A(n232), .B(r_y_data[15]), .C(r_mult_1_B[15]), .D(n169), 
        .Y(n334) );
  oa21d1_hd U1055 ( .A(n167), .B(n183), .C(n334), .Y(n485) );
  ao22d1_hd U1056 ( .A(n232), .B(r_y_data[14]), .C(r_mult_1_B[14]), .D(n169), 
        .Y(n335) );
  oa21d1_hd U1057 ( .A(n167), .B(n184), .C(n335), .Y(n486) );
  ao22d1_hd U1058 ( .A(n232), .B(r_y_data[13]), .C(r_mult_1_B[13]), .D(n169), 
        .Y(n336) );
  oa21d1_hd U1059 ( .A(n167), .B(n185), .C(n336), .Y(n487) );
  ao22d1_hd U1060 ( .A(n232), .B(r_y_data[12]), .C(r_mult_1_B[12]), .D(n169), 
        .Y(n337) );
  oa21d1_hd U1061 ( .A(n167), .B(n186), .C(n337), .Y(n488) );
  ao22d1_hd U1062 ( .A(n232), .B(r_y_data[11]), .C(r_mult_1_B[11]), .D(n169), 
        .Y(n338) );
  oa21d1_hd U1063 ( .A(n167), .B(n187), .C(n338), .Y(n489) );
  ao22d1_hd U1064 ( .A(n232), .B(r_y_data[10]), .C(r_mult_1_B[10]), .D(n169), 
        .Y(n339) );
  oa21d1_hd U1065 ( .A(n167), .B(n188), .C(n339), .Y(n490) );
  ao22d1_hd U1066 ( .A(n232), .B(r_y_data[9]), .C(r_mult_1_B[9]), .D(n169), 
        .Y(n340) );
  oa21d1_hd U1067 ( .A(n167), .B(n189), .C(n340), .Y(n491) );
  ao22d1_hd U1068 ( .A(n232), .B(r_y_data[8]), .C(r_mult_1_B[8]), .D(n169), 
        .Y(n341) );
  oa21d1_hd U1069 ( .A(n167), .B(n190), .C(n341), .Y(n492) );
  ao22d1_hd U1070 ( .A(n232), .B(r_y_data[7]), .C(r_mult_1_B[7]), .D(n169), 
        .Y(n342) );
  oa21d1_hd U1071 ( .A(n167), .B(n191), .C(n342), .Y(n493) );
  ao22d1_hd U1072 ( .A(n232), .B(r_y_data[6]), .C(r_mult_1_B[6]), .D(n169), 
        .Y(n343) );
  oa21d1_hd U1073 ( .A(n167), .B(n192), .C(n343), .Y(n494) );
  ao22d1_hd U1074 ( .A(n232), .B(r_y_data[5]), .C(r_mult_1_B[5]), .D(n169), 
        .Y(n344) );
  oa21d1_hd U1075 ( .A(n167), .B(n193), .C(n344), .Y(n495) );
  ao22d1_hd U1076 ( .A(n232), .B(r_y_data[4]), .C(r_mult_1_B[4]), .D(n169), 
        .Y(n345) );
  oa21d1_hd U1077 ( .A(n167), .B(n194), .C(n345), .Y(n496) );
  ao22d1_hd U1078 ( .A(n232), .B(r_y_data[3]), .C(r_mult_1_B[3]), .D(n169), 
        .Y(n346) );
  oa21d1_hd U1079 ( .A(n167), .B(n195), .C(n346), .Y(n497) );
  ao22d1_hd U1080 ( .A(n232), .B(r_y_data[2]), .C(r_mult_1_B[2]), .D(n169), 
        .Y(n347) );
  oa21d1_hd U1081 ( .A(n167), .B(n196), .C(n347), .Y(n498) );
  ao22d1_hd U1082 ( .A(n232), .B(r_y_data[1]), .C(r_mult_1_B[1]), .D(n169), 
        .Y(n348) );
  oa21d1_hd U1083 ( .A(n167), .B(n197), .C(n348), .Y(n499) );
  ao22d1_hd U1084 ( .A(n232), .B(r_y_data[0]), .C(r_mult_1_B[0]), .D(n169), 
        .Y(n349) );
  oa21d1_hd U1085 ( .A(n167), .B(n198), .C(n349), .Y(n500) );
  ao22d1_hd U1086 ( .A(n232), .B(r_x_data[30]), .C(r_add_A[30]), .D(n231), .Y(
        n533) );
  ao22d1_hd U1087 ( .A(n234), .B(w_mult_1_Z[30]), .C(n233), .D(w_mult_2_Z[30]), 
        .Y(n351) );
  oa211d1_hd U1088 ( .A(n721), .B(n645), .C(n533), .D(n351), .Y(n501) );
  ao22d1_hd U1089 ( .A(n232), .B(r_x_data[29]), .C(r_add_A[29]), .D(n231), .Y(
        n573) );
  ao22d1_hd U1090 ( .A(n234), .B(w_mult_1_Z[29]), .C(n233), .D(w_mult_2_Z[29]), 
        .Y(n534) );
  oa211d1_hd U1091 ( .A(n721), .B(n647), .C(n573), .D(n534), .Y(n502) );
  ao22d1_hd U1092 ( .A(n232), .B(r_x_data[28]), .C(r_add_A[28]), .D(n231), .Y(
        n575) );
  ao22d1_hd U1093 ( .A(n234), .B(w_mult_1_Z[28]), .C(n233), .D(w_mult_2_Z[28]), 
        .Y(n574) );
  oa211d1_hd U1094 ( .A(n721), .B(n649), .C(n575), .D(n574), .Y(n503) );
  ao22d1_hd U1095 ( .A(n232), .B(r_x_data[27]), .C(r_add_A[27]), .D(n231), .Y(
        n577) );
  ao22d1_hd U1096 ( .A(n234), .B(w_mult_1_Z[27]), .C(n233), .D(w_mult_2_Z[27]), 
        .Y(n576) );
  oa211d1_hd U1097 ( .A(n721), .B(n651), .C(n577), .D(n576), .Y(n504) );
  ao22d1_hd U1098 ( .A(n232), .B(r_x_data[26]), .C(r_add_A[26]), .D(n231), .Y(
        n579) );
  ao22d1_hd U1099 ( .A(n234), .B(w_mult_1_Z[26]), .C(n233), .D(w_mult_2_Z[26]), 
        .Y(n578) );
  oa211d1_hd U1100 ( .A(n721), .B(n653), .C(n579), .D(n578), .Y(n505) );
  ao22d1_hd U1101 ( .A(n232), .B(r_x_data[25]), .C(r_add_A[25]), .D(n231), .Y(
        n582) );
  ao22d1_hd U1102 ( .A(n234), .B(w_mult_1_Z[25]), .C(n233), .D(w_mult_2_Z[25]), 
        .Y(n581) );
  oa211d1_hd U1103 ( .A(n721), .B(n655), .C(n582), .D(n581), .Y(n506) );
  ao22d1_hd U1104 ( .A(n232), .B(r_x_data[24]), .C(r_add_A[24]), .D(n231), .Y(
        n584) );
  ao22d1_hd U1105 ( .A(n234), .B(w_mult_1_Z[24]), .C(n233), .D(w_mult_2_Z[24]), 
        .Y(n583) );
  oa211d1_hd U1106 ( .A(n721), .B(n657), .C(n584), .D(n583), .Y(n507) );
  ao22d1_hd U1107 ( .A(n232), .B(r_x_data[23]), .C(r_add_A[23]), .D(n231), .Y(
        n586) );
  ao22d1_hd U1108 ( .A(n234), .B(w_mult_1_Z[23]), .C(n233), .D(w_mult_2_Z[23]), 
        .Y(n585) );
  oa211d1_hd U1109 ( .A(n721), .B(n659), .C(n586), .D(n585), .Y(n508) );
  ao22d1_hd U1110 ( .A(n232), .B(r_x_data[22]), .C(r_add_A[22]), .D(n231), .Y(
        n588) );
  ao22d1_hd U1111 ( .A(n234), .B(w_mult_1_Z[22]), .C(n233), .D(w_mult_2_Z[22]), 
        .Y(n587) );
  oa211d1_hd U1112 ( .A(n721), .B(n661), .C(n588), .D(n587), .Y(n509) );
  ao22d1_hd U1113 ( .A(n232), .B(r_x_data[21]), .C(r_add_A[21]), .D(n231), .Y(
        n590) );
  ao22d1_hd U1114 ( .A(n234), .B(w_mult_1_Z[21]), .C(n233), .D(w_mult_2_Z[21]), 
        .Y(n589) );
  oa211d1_hd U1115 ( .A(n721), .B(n663), .C(n590), .D(n589), .Y(n510) );
  ao22d1_hd U1116 ( .A(n232), .B(r_x_data[20]), .C(r_add_A[20]), .D(n231), .Y(
        n592) );
  ao22d1_hd U1117 ( .A(n234), .B(w_mult_1_Z[20]), .C(n233), .D(w_mult_2_Z[20]), 
        .Y(n591) );
  oa211d1_hd U1118 ( .A(n721), .B(n665), .C(n592), .D(n591), .Y(n511) );
  ao22d1_hd U1119 ( .A(n232), .B(r_x_data[19]), .C(r_add_A[19]), .D(n231), .Y(
        n594) );
  ao22d1_hd U1120 ( .A(n234), .B(w_mult_1_Z[19]), .C(n233), .D(w_mult_2_Z[19]), 
        .Y(n593) );
  oa211d1_hd U1121 ( .A(n721), .B(n667), .C(n594), .D(n593), .Y(n512) );
  ao22d1_hd U1122 ( .A(n232), .B(r_x_data[18]), .C(r_add_A[18]), .D(n231), .Y(
        n596) );
  ao22d1_hd U1123 ( .A(n234), .B(w_mult_1_Z[18]), .C(n233), .D(w_mult_2_Z[18]), 
        .Y(n595) );
  oa211d1_hd U1124 ( .A(n721), .B(n669), .C(n596), .D(n595), .Y(n513) );
  ao22d1_hd U1125 ( .A(n232), .B(r_x_data[17]), .C(r_add_A[17]), .D(n231), .Y(
        n598) );
  ao22d1_hd U1126 ( .A(n717), .B(w_mult_1_Z[17]), .C(n233), .D(w_mult_2_Z[17]), 
        .Y(n597) );
  oa211d1_hd U1127 ( .A(n721), .B(n671), .C(n598), .D(n597), .Y(n514) );
  ao22d1_hd U1128 ( .A(n232), .B(r_x_data[16]), .C(r_add_A[16]), .D(n231), .Y(
        n600) );
  ao22d1_hd U1129 ( .A(n717), .B(w_mult_1_Z[16]), .C(n233), .D(w_mult_2_Z[16]), 
        .Y(n599) );
  oa211d1_hd U1130 ( .A(n721), .B(n673), .C(n600), .D(n599), .Y(n515) );
  ao22d1_hd U1131 ( .A(n232), .B(r_x_data[15]), .C(r_add_A[15]), .D(n231), .Y(
        n602) );
  ao22d1_hd U1132 ( .A(n717), .B(w_mult_1_Z[15]), .C(n233), .D(w_mult_2_Z[15]), 
        .Y(n601) );
  oa211d1_hd U1133 ( .A(n721), .B(n675), .C(n602), .D(n601), .Y(n516) );
  ao22d1_hd U1134 ( .A(n232), .B(r_x_data[14]), .C(r_add_A[14]), .D(n231), .Y(
        n604) );
  ao22d1_hd U1135 ( .A(n717), .B(w_mult_1_Z[14]), .C(n233), .D(w_mult_2_Z[14]), 
        .Y(n603) );
  oa211d1_hd U1136 ( .A(n721), .B(n677), .C(n604), .D(n603), .Y(n517) );
  ao22d1_hd U1137 ( .A(n232), .B(r_x_data[13]), .C(r_add_A[13]), .D(n231), .Y(
        n606) );
  ao22d1_hd U1138 ( .A(n234), .B(w_mult_1_Z[13]), .C(n716), .D(w_mult_2_Z[13]), 
        .Y(n605) );
  oa211d1_hd U1139 ( .A(n721), .B(n679), .C(n606), .D(n605), .Y(n518) );
  ao22d1_hd U1140 ( .A(n232), .B(r_x_data[12]), .C(r_add_A[12]), .D(n714), .Y(
        n608) );
  ao22d1_hd U1141 ( .A(n234), .B(w_mult_1_Z[12]), .C(n716), .D(w_mult_2_Z[12]), 
        .Y(n607) );
  oa211d1_hd U1142 ( .A(n721), .B(n681), .C(n608), .D(n607), .Y(n519) );
  ao22d1_hd U1143 ( .A(n232), .B(r_x_data[11]), .C(r_add_A[11]), .D(n714), .Y(
        n610) );
  ao22d1_hd U1144 ( .A(n234), .B(w_mult_1_Z[11]), .C(n716), .D(w_mult_2_Z[11]), 
        .Y(n609) );
  oa211d1_hd U1145 ( .A(n721), .B(n683), .C(n610), .D(n609), .Y(n520) );
  ao22d1_hd U1146 ( .A(n232), .B(r_x_data[10]), .C(r_add_A[10]), .D(n714), .Y(
        n612) );
  ao22d1_hd U1147 ( .A(n717), .B(w_mult_1_Z[10]), .C(n233), .D(w_mult_2_Z[10]), 
        .Y(n611) );
  oa211d1_hd U1148 ( .A(n721), .B(n685), .C(n612), .D(n611), .Y(n521) );
  ao22d1_hd U1149 ( .A(n232), .B(r_x_data[9]), .C(r_add_A[9]), .D(n231), .Y(
        n614) );
  ao22d1_hd U1150 ( .A(n234), .B(w_mult_1_Z[9]), .C(n233), .D(w_mult_2_Z[9]), 
        .Y(n613) );
  oa211d1_hd U1151 ( .A(n721), .B(n687), .C(n614), .D(n613), .Y(n522) );
  ao22d1_hd U1152 ( .A(n232), .B(r_x_data[8]), .C(r_add_A[8]), .D(n231), .Y(
        n616) );
  ao22d1_hd U1153 ( .A(n234), .B(w_mult_1_Z[8]), .C(n233), .D(w_mult_2_Z[8]), 
        .Y(n615) );
  oa211d1_hd U1154 ( .A(n721), .B(n689), .C(n616), .D(n615), .Y(n523) );
  ao22d1_hd U1155 ( .A(n232), .B(r_x_data[7]), .C(r_add_A[7]), .D(n231), .Y(
        n618) );
  ao22d1_hd U1156 ( .A(n234), .B(w_mult_1_Z[7]), .C(n716), .D(w_mult_2_Z[7]), 
        .Y(n617) );
  oa211d1_hd U1157 ( .A(n721), .B(n691), .C(n618), .D(n617), .Y(n524) );
  ao22d1_hd U1158 ( .A(n232), .B(r_x_data[6]), .C(r_add_A[6]), .D(n231), .Y(
        n620) );
  ao22d1_hd U1159 ( .A(n234), .B(w_mult_1_Z[6]), .C(n233), .D(w_mult_2_Z[6]), 
        .Y(n619) );
  oa211d1_hd U1160 ( .A(n721), .B(n693), .C(n620), .D(n619), .Y(n525) );
  ao22d1_hd U1161 ( .A(n232), .B(r_x_data[5]), .C(r_add_A[5]), .D(n231), .Y(
        n622) );
  ao22d1_hd U1162 ( .A(n234), .B(w_mult_1_Z[5]), .C(n233), .D(w_mult_2_Z[5]), 
        .Y(n621) );
  oa211d1_hd U1163 ( .A(n721), .B(n695), .C(n622), .D(n621), .Y(n526) );
  ao22d1_hd U1164 ( .A(n232), .B(r_x_data[4]), .C(r_add_A[4]), .D(n231), .Y(
        n624) );
  ao22d1_hd U1165 ( .A(n234), .B(w_mult_1_Z[4]), .C(n233), .D(w_mult_2_Z[4]), 
        .Y(n623) );
  oa211d1_hd U1166 ( .A(n721), .B(n697), .C(n624), .D(n623), .Y(n527) );
  ao22d1_hd U1167 ( .A(n232), .B(r_x_data[3]), .C(r_add_A[3]), .D(n231), .Y(
        n626) );
  ao22d1_hd U1168 ( .A(n234), .B(w_mult_1_Z[3]), .C(n233), .D(w_mult_2_Z[3]), 
        .Y(n625) );
  oa211d1_hd U1169 ( .A(n721), .B(n699), .C(n626), .D(n625), .Y(n528) );
  ao22d1_hd U1170 ( .A(n232), .B(r_x_data[2]), .C(r_add_A[2]), .D(n231), .Y(
        n628) );
  ao22d1_hd U1171 ( .A(n234), .B(w_mult_1_Z[2]), .C(n233), .D(w_mult_2_Z[2]), 
        .Y(n627) );
  oa211d1_hd U1172 ( .A(n721), .B(n701), .C(n628), .D(n627), .Y(n529) );
  ao22d1_hd U1173 ( .A(n232), .B(r_x_data[1]), .C(r_add_A[1]), .D(n231), .Y(
        n630) );
  ao22d1_hd U1174 ( .A(n234), .B(w_mult_1_Z[1]), .C(n233), .D(w_mult_2_Z[1]), 
        .Y(n629) );
  oa211d1_hd U1175 ( .A(n721), .B(n703), .C(n630), .D(n629), .Y(n530) );
  scg6d1_hd U1176 ( .A(r_add_Z_ACK), .B(n632), .C(n631), .Y(n531) );
  scg14d1_hd U1177 ( .A(r_add_AB_STB), .B(n641), .C(n639), .Y(n535) );
  ao22d1_hd U1178 ( .A(n232), .B(r_y_data[63]), .C(r_mult_2_B[31]), .D(n169), 
        .Y(n636) );
  scg14d1_hd U1179 ( .A(w_add_Z[31]), .B(n350), .C(n636), .Y(n536) );
  ao22d1_hd U1180 ( .A(w_add_Z[30]), .B(n230), .C(w_mult_1_Z[30]), .D(n229), 
        .Y(n644) );
  oa21d1_hd U1181 ( .A(n645), .B(n710), .C(n644), .Y(n537) );
  ao22d1_hd U1182 ( .A(w_add_Z[29]), .B(n230), .C(w_mult_1_Z[29]), .D(n229), 
        .Y(n646) );
  oa21d1_hd U1183 ( .A(n647), .B(n710), .C(n646), .Y(n538) );
  ao22d1_hd U1184 ( .A(w_add_Z[28]), .B(n230), .C(w_mult_1_Z[28]), .D(n229), 
        .Y(n648) );
  oa21d1_hd U1185 ( .A(n649), .B(n710), .C(n648), .Y(n539) );
  ao22d1_hd U1186 ( .A(w_add_Z[27]), .B(n230), .C(w_mult_1_Z[27]), .D(n229), 
        .Y(n650) );
  oa21d1_hd U1187 ( .A(n651), .B(n710), .C(n650), .Y(n540) );
  ao22d1_hd U1188 ( .A(w_add_Z[26]), .B(n230), .C(w_mult_1_Z[26]), .D(n229), 
        .Y(n652) );
  oa21d1_hd U1189 ( .A(n653), .B(n710), .C(n652), .Y(n541) );
  ao22d1_hd U1190 ( .A(w_add_Z[25]), .B(n230), .C(w_mult_1_Z[25]), .D(n229), 
        .Y(n654) );
  oa21d1_hd U1191 ( .A(n655), .B(n710), .C(n654), .Y(n542) );
  ao22d1_hd U1192 ( .A(w_add_Z[24]), .B(n230), .C(w_mult_1_Z[24]), .D(n229), 
        .Y(n656) );
  oa21d1_hd U1193 ( .A(n657), .B(n710), .C(n656), .Y(n543) );
  ao22d1_hd U1194 ( .A(w_add_Z[23]), .B(n708), .C(w_mult_1_Z[23]), .D(n229), 
        .Y(n658) );
  oa21d1_hd U1195 ( .A(n659), .B(n710), .C(n658), .Y(n544) );
  ao22d1_hd U1196 ( .A(w_add_Z[22]), .B(n708), .C(w_mult_1_Z[22]), .D(n229), 
        .Y(n660) );
  oa21d1_hd U1197 ( .A(n661), .B(n710), .C(n660), .Y(n545) );
  ao22d1_hd U1198 ( .A(w_add_Z[21]), .B(n230), .C(w_mult_1_Z[21]), .D(n229), 
        .Y(n662) );
  oa21d1_hd U1199 ( .A(n663), .B(n710), .C(n662), .Y(n546) );
  ao22d1_hd U1200 ( .A(w_add_Z[20]), .B(n230), .C(w_mult_1_Z[20]), .D(n229), 
        .Y(n664) );
  oa21d1_hd U1201 ( .A(n665), .B(n710), .C(n664), .Y(n547) );
  ao22d1_hd U1202 ( .A(w_add_Z[19]), .B(n230), .C(w_mult_1_Z[19]), .D(n707), 
        .Y(n666) );
  oa21d1_hd U1203 ( .A(n667), .B(n710), .C(n666), .Y(n548) );
  ao22d1_hd U1204 ( .A(w_add_Z[18]), .B(n230), .C(w_mult_1_Z[18]), .D(n707), 
        .Y(n668) );
  oa21d1_hd U1205 ( .A(n669), .B(n710), .C(n668), .Y(n549) );
  ao22d1_hd U1206 ( .A(w_add_Z[17]), .B(n230), .C(w_mult_1_Z[17]), .D(n707), 
        .Y(n670) );
  oa21d1_hd U1207 ( .A(n671), .B(n710), .C(n670), .Y(n550) );
  ao22d1_hd U1208 ( .A(w_add_Z[16]), .B(n230), .C(w_mult_1_Z[16]), .D(n229), 
        .Y(n672) );
  oa21d1_hd U1209 ( .A(n673), .B(n710), .C(n672), .Y(n551) );
  ao22d1_hd U1210 ( .A(w_add_Z[15]), .B(n230), .C(w_mult_1_Z[15]), .D(n229), 
        .Y(n674) );
  oa21d1_hd U1211 ( .A(n675), .B(n710), .C(n674), .Y(n552) );
  ao22d1_hd U1212 ( .A(w_add_Z[14]), .B(n230), .C(w_mult_1_Z[14]), .D(n229), 
        .Y(n676) );
  oa21d1_hd U1213 ( .A(n677), .B(n710), .C(n676), .Y(n553) );
  ao22d1_hd U1214 ( .A(w_add_Z[13]), .B(n230), .C(w_mult_1_Z[13]), .D(n229), 
        .Y(n678) );
  oa21d1_hd U1215 ( .A(n679), .B(n710), .C(n678), .Y(n554) );
  ao22d1_hd U1216 ( .A(w_add_Z[12]), .B(n230), .C(w_mult_1_Z[12]), .D(n229), 
        .Y(n680) );
  oa21d1_hd U1217 ( .A(n681), .B(n710), .C(n680), .Y(n555) );
  ao22d1_hd U1218 ( .A(w_add_Z[11]), .B(n708), .C(w_mult_1_Z[11]), .D(n229), 
        .Y(n682) );
  oa21d1_hd U1219 ( .A(n683), .B(n710), .C(n682), .Y(n556) );
  ao22d1_hd U1220 ( .A(w_add_Z[10]), .B(n708), .C(w_mult_1_Z[10]), .D(n229), 
        .Y(n684) );
  oa21d1_hd U1221 ( .A(n685), .B(n710), .C(n684), .Y(n557) );
  ao22d1_hd U1222 ( .A(w_add_Z[9]), .B(n230), .C(w_mult_1_Z[9]), .D(n229), .Y(
        n686) );
  oa21d1_hd U1223 ( .A(n687), .B(n710), .C(n686), .Y(n558) );
  ao22d1_hd U1224 ( .A(w_add_Z[8]), .B(n230), .C(w_mult_1_Z[8]), .D(n229), .Y(
        n688) );
  oa21d1_hd U1225 ( .A(n689), .B(n710), .C(n688), .Y(n559) );
  ao22d1_hd U1226 ( .A(w_add_Z[7]), .B(n230), .C(w_mult_1_Z[7]), .D(n229), .Y(
        n690) );
  oa21d1_hd U1227 ( .A(n691), .B(n710), .C(n690), .Y(n560) );
  ao22d1_hd U1228 ( .A(w_add_Z[6]), .B(n230), .C(w_mult_1_Z[6]), .D(n229), .Y(
        n692) );
  oa21d1_hd U1229 ( .A(n693), .B(n710), .C(n692), .Y(n561) );
  ao22d1_hd U1230 ( .A(w_add_Z[5]), .B(n230), .C(w_mult_1_Z[5]), .D(n229), .Y(
        n694) );
  oa21d1_hd U1231 ( .A(n695), .B(n710), .C(n694), .Y(n562) );
  ao22d1_hd U1232 ( .A(w_add_Z[4]), .B(n230), .C(w_mult_1_Z[4]), .D(n229), .Y(
        n696) );
  oa21d1_hd U1233 ( .A(n697), .B(n710), .C(n696), .Y(n563) );
  ao22d1_hd U1234 ( .A(w_add_Z[3]), .B(n230), .C(w_mult_1_Z[3]), .D(n229), .Y(
        n698) );
  oa21d1_hd U1235 ( .A(n699), .B(n710), .C(n698), .Y(n564) );
  ao22d1_hd U1236 ( .A(w_add_Z[2]), .B(n230), .C(w_mult_1_Z[2]), .D(n229), .Y(
        n700) );
  oa21d1_hd U1237 ( .A(n701), .B(n710), .C(n700), .Y(n565) );
  ao22d1_hd U1238 ( .A(w_add_Z[1]), .B(n230), .C(w_mult_1_Z[1]), .D(n229), .Y(
        n702) );
  oa21d1_hd U1239 ( .A(n703), .B(n710), .C(n702), .Y(n566) );
  ao22d1_hd U1240 ( .A(w_add_Z[0]), .B(n230), .C(w_mult_1_Z[0]), .D(n229), .Y(
        n704) );
  oa21d1_hd U1241 ( .A(n720), .B(n710), .C(n704), .Y(n567) );
  ao22d1_hd U1242 ( .A(n232), .B(r_y_data[31]), .C(r_mult_1_B[31]), .D(n169), 
        .Y(n706) );
  scg14d1_hd U1243 ( .A(n350), .B(r_x_data[63]), .C(n706), .Y(n568) );
  ao22d1_hd U1244 ( .A(w_add_Z[31]), .B(n230), .C(w_mult_1_Z[31]), .D(n229), 
        .Y(n709) );
  oa21d1_hd U1245 ( .A(n713), .B(n710), .C(n709), .Y(n569) );
  ao22d1_hd U1246 ( .A(n232), .B(r_x_data[31]), .C(r_add_A[31]), .D(n231), .Y(
        n712) );
  ao22d1_hd U1247 ( .A(n234), .B(w_mult_1_Z[31]), .C(w_mult_2_Z[31]), .D(n233), 
        .Y(n711) );
  oa211d1_hd U1248 ( .A(n721), .B(n713), .C(n712), .D(n711), .Y(n570) );
  ao22d1_hd U1249 ( .A(n232), .B(r_x_data[0]), .C(r_add_A[0]), .D(n231), .Y(
        n719) );
  ao22d1_hd U1250 ( .A(n234), .B(w_mult_1_Z[0]), .C(n233), .D(w_mult_2_Z[0]), 
        .Y(n718) );
  oa211d1_hd U1251 ( .A(n721), .B(n720), .C(n719), .D(n718), .Y(n571) );
endmodule


module float_adder_1 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3, C91_DATA2_4,
         C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8, n1, n2, n27, n266,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n509, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23, C2_Z_22,
         C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16, C2_Z_15,
         C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8, C2_Z_7,
         C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_43J4_124_6938_n58, DP_OP_43J4_124_6938_n57,
         DP_OP_43J4_124_6938_n56, DP_OP_43J4_124_6938_n55,
         DP_OP_43J4_124_6938_n54, DP_OP_43J4_124_6938_n53,
         DP_OP_43J4_124_6938_n52, DP_OP_43J4_124_6938_n51,
         DP_OP_43J4_124_6938_n50, DP_OP_43J4_124_6938_n49,
         DP_OP_43J4_124_6938_n48, DP_OP_43J4_124_6938_n47,
         DP_OP_43J4_124_6938_n46, DP_OP_43J4_124_6938_n45,
         DP_OP_43J4_124_6938_n44, DP_OP_43J4_124_6938_n43,
         DP_OP_43J4_124_6938_n42, DP_OP_43J4_124_6938_n41,
         DP_OP_43J4_124_6938_n40, DP_OP_43J4_124_6938_n39,
         DP_OP_43J4_124_6938_n38, DP_OP_43J4_124_6938_n37,
         DP_OP_43J4_124_6938_n36, DP_OP_43J4_124_6938_n35,
         DP_OP_43J4_124_6938_n34, DP_OP_43J4_124_6938_n33,
         DP_OP_43J4_124_6938_n32, DP_OP_43J4_124_6938_n27,
         DP_OP_43J4_124_6938_n26, DP_OP_43J4_124_6938_n25,
         DP_OP_43J4_124_6938_n24, DP_OP_43J4_124_6938_n23,
         DP_OP_43J4_124_6938_n22, DP_OP_43J4_124_6938_n21,
         DP_OP_43J4_124_6938_n20, DP_OP_43J4_124_6938_n19,
         DP_OP_43J4_124_6938_n18, DP_OP_43J4_124_6938_n17,
         DP_OP_43J4_124_6938_n16, DP_OP_43J4_124_6938_n15,
         DP_OP_43J4_124_6938_n14, DP_OP_43J4_124_6938_n13,
         DP_OP_43J4_124_6938_n12, DP_OP_43J4_124_6938_n11,
         DP_OP_43J4_124_6938_n10, DP_OP_43J4_124_6938_n9,
         DP_OP_43J4_124_6938_n8, DP_OP_43J4_124_6938_n7,
         DP_OP_43J4_124_6938_n6, DP_OP_43J4_124_6938_n5,
         DP_OP_43J4_124_6938_n4, DP_OP_43J4_124_6938_n3,
         DP_OP_43J4_124_6938_n2, DP_OP_43J4_124_6938_n1,
         DP_OP_154J4_137_6175_n9, DP_OP_154J4_137_6175_n8,
         DP_OP_154J4_137_6175_n7, DP_OP_154J4_137_6175_n6,
         DP_OP_154J4_137_6175_n5, DP_OP_154J4_137_6175_n4,
         DP_OP_154J4_137_6175_n3, DP_OP_154J4_137_6175_n2, n1895, n1222, n1284,
         n1285, n1291, n1891, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J4_137_6175_U10 ( .A(n1291), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J4_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J4_137_6175_U9 ( .A(n1291), .B(z_e[2]), .CI(
        DP_OP_154J4_137_6175_n9), .CO(DP_OP_154J4_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J4_137_6175_U8 ( .A(n1291), .B(z_e[3]), .CI(
        DP_OP_154J4_137_6175_n8), .CO(DP_OP_154J4_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J4_137_6175_U7 ( .A(n1291), .B(z_e[4]), .CI(
        DP_OP_154J4_137_6175_n7), .CO(DP_OP_154J4_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J4_137_6175_U6 ( .A(n1291), .B(z_e[5]), .CI(
        DP_OP_154J4_137_6175_n6), .CO(DP_OP_154J4_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J4_137_6175_U5 ( .A(n1291), .B(z_e[6]), .CI(
        DP_OP_154J4_137_6175_n5), .CO(DP_OP_154J4_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J4_137_6175_U4 ( .A(n1291), .B(z_e[7]), .CI(
        DP_OP_154J4_137_6175_n4), .CO(DP_OP_154J4_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J4_137_6175_U3 ( .A(n1291), .B(z_e[8]), .CI(
        DP_OP_154J4_137_6175_n3), .CO(DP_OP_154J4_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n2281), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n2281), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n509), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n2281), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n2281), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n2281), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n2281), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n2281), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n509), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n509), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n509), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n509), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n2281), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n2281), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n2281), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n2281), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n2281), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n2281), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n2281), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n2281), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n2281), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n509), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n2281), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n2281), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n2281), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n2281), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n2281), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n2281), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n2281), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n2281), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n2281), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n2282), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n2282), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n2282), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n2282), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n2268), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n2268), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n2282), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n2282), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n2282), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n2282), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n2282), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n27), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n2282), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n2282), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n2282), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n27), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n27), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n27), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n27), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n27), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n27), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n2282), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n27), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n2282), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n2282), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n27), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n27), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n2282), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n2282), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n2282), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n2282), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n2282), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n2282), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n2282), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n2282), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n2282), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n2282), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n2282), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n2282), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n2282), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n2282), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n2282), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n2282), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n2282), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n2282), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n2282), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n2282), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n2282), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n2282), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n2282), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n2282), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n2282), .CK(i_CLK), .Q(b[22]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n2268), .CK(i_CLK), .Q(sum[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n2268), .CK(i_CLK), .Q(sum[2]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n2268), .CK(i_CLK), .Q(sum[26]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n2268), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n2268), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n2268), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n2268), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n2268), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n2268), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n2268), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n2268), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n2268), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n2268), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n2268), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n2268), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n2268), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n2268), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n2268), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n2268), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n2268), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n2268), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n2268), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n2268), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n2268), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n2268), .CK(i_CLK), .Q(sum[25]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n2268), .CK(i_CLK), .Q(sum[1]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n2282), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n2282), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n2282), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n2282), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n2268), .CK(i_CLK), .Q(sum[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n2282), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n2282), .CK(i_CLK), .Q(b[28]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n2282), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n2282), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n2282), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n2282), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n2282), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n2282), .CK(i_CLK), .Q(b[26]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n2282), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n2282), .CK(i_CLK), .Q(b[23]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n1222), .CK(i_CLK), .Q(guard) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n2277), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n2277), .CK(i_CLK), .Q(a_s) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n1895), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n1895), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J4_124_6938_U28 ( .A(C2_Z_0), .B(n1891), .CI(
        DP_OP_43J4_124_6938_n58), .CO(DP_OP_43J4_124_6938_n27), .S(N310) );
  fad1_hd DP_OP_43J4_124_6938_U27 ( .A(DP_OP_43J4_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J4_124_6938_n27), .CO(DP_OP_43J4_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J4_124_6938_U26 ( .A(DP_OP_43J4_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J4_124_6938_n26), .CO(DP_OP_43J4_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J4_124_6938_U25 ( .A(DP_OP_43J4_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J4_124_6938_n25), .CO(DP_OP_43J4_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J4_124_6938_U2 ( .A(DP_OP_43J4_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J4_124_6938_n2), .CO(DP_OP_43J4_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J4_124_6938_U16 ( .A(DP_OP_43J4_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J4_124_6938_n16), .CO(DP_OP_43J4_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J4_124_6938_U17 ( .A(DP_OP_43J4_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J4_124_6938_n17), .CO(DP_OP_43J4_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J4_124_6938_U18 ( .A(DP_OP_43J4_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J4_124_6938_n18), .CO(DP_OP_43J4_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J4_124_6938_U19 ( .A(DP_OP_43J4_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J4_124_6938_n19), .CO(DP_OP_43J4_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J4_124_6938_U20 ( .A(DP_OP_43J4_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J4_124_6938_n20), .CO(DP_OP_43J4_124_6938_n19), .S(N318)
         );
  fad1_hd DP_OP_43J4_124_6938_U21 ( .A(DP_OP_43J4_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J4_124_6938_n21), .CO(DP_OP_43J4_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J4_124_6938_U22 ( .A(DP_OP_43J4_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J4_124_6938_n22), .CO(DP_OP_43J4_124_6938_n21), .S(N316)
         );
  fad1_hd DP_OP_43J4_124_6938_U23 ( .A(DP_OP_43J4_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J4_124_6938_n23), .CO(DP_OP_43J4_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J4_124_6938_U24 ( .A(DP_OP_43J4_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J4_124_6938_n24), .CO(DP_OP_43J4_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J4_124_6938_U15 ( .A(DP_OP_43J4_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J4_124_6938_n15), .CO(DP_OP_43J4_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J4_124_6938_U14 ( .A(DP_OP_43J4_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J4_124_6938_n14), .CO(DP_OP_43J4_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J4_124_6938_U13 ( .A(DP_OP_43J4_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J4_124_6938_n13), .CO(DP_OP_43J4_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J4_124_6938_U12 ( .A(DP_OP_43J4_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J4_124_6938_n12), .CO(DP_OP_43J4_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J4_124_6938_U5 ( .A(DP_OP_43J4_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J4_124_6938_n5), .CO(DP_OP_43J4_124_6938_n4), .S(N333) );
  fad1_hd DP_OP_43J4_124_6938_U4 ( .A(DP_OP_43J4_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J4_124_6938_n4), .CO(DP_OP_43J4_124_6938_n3), .S(N334) );
  fad1_hd DP_OP_43J4_124_6938_U3 ( .A(DP_OP_43J4_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J4_124_6938_n3), .CO(DP_OP_43J4_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J4_124_6938_U11 ( .A(DP_OP_43J4_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J4_124_6938_n11), .CO(DP_OP_43J4_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J4_124_6938_U10 ( .A(DP_OP_43J4_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J4_124_6938_n10), .CO(DP_OP_43J4_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J4_124_6938_U9 ( .A(DP_OP_43J4_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J4_124_6938_n9), .CO(DP_OP_43J4_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J4_124_6938_U8 ( .A(DP_OP_43J4_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J4_124_6938_n8), .CO(DP_OP_43J4_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J4_124_6938_U7 ( .A(DP_OP_43J4_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J4_124_6938_n7), .CO(DP_OP_43J4_124_6938_n6), .S(N331) );
  fad1_hd DP_OP_43J4_124_6938_U6 ( .A(DP_OP_43J4_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J4_124_6938_n6), .CO(DP_OP_43J4_124_6938_n5), .S(N332) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  clknd2d1_hd U523 ( .A(a_m[24]), .B(n2698), .Y(n2321) );
  clknd2d1_hd U524 ( .A(a_m[7]), .B(n2732), .Y(n2291) );
  clknd2d1_hd U525 ( .A(a_m[11]), .B(n2724), .Y(n2298) );
  clknd2d1_hd U526 ( .A(a_e[3]), .B(n2898), .Y(n2391) );
  clknd2d1_hd U527 ( .A(b_e[6]), .B(n2803), .Y(n2394) );
  clknd2d1_hd U528 ( .A(b_m[19]), .B(n2756), .Y(n2311) );
  clknd2d1_hd U529 ( .A(a_m[18]), .B(n2710), .Y(n2309) );
  clknd2d1_hd U530 ( .A(n2381), .B(n2394), .Y(n2387) );
  clknd2d1_hd U531 ( .A(z_e[7]), .B(z_e[8]), .Y(n2501) );
  clknd2d1_hd U532 ( .A(b_e[0]), .B(n2838), .Y(n2382) );
  clknd2d1_hd U533 ( .A(b_e[4]), .B(n2888), .Y(n2864) );
  clknd2d1_hd U534 ( .A(b_e[6]), .B(b_e[5]), .Y(n2865) );
  clknd2d1_hd U535 ( .A(n2889), .B(n2406), .Y(n2928) );
  ad2bd1_hd U536 ( .B(n2514), .AN(n1222), .Y(n2635) );
  clknd2d1_hd U537 ( .A(n2657), .B(n2512), .Y(n2513) );
  clknd2d1_hd U538 ( .A(n2415), .B(n2413), .Y(n2434) );
  clknd2d1_hd U539 ( .A(n2427), .B(n2472), .Y(n2502) );
  clknd2d1_hd U540 ( .A(n2863), .B(n2412), .Y(n2410) );
  clknd2d1_hd U541 ( .A(n2797), .B(n2414), .Y(n2450) );
  clknd2d1_hd U542 ( .A(n2947), .B(n2942), .Y(n2667) );
  clknd2d1_hd U543 ( .A(a_e[2]), .B(n2841), .Y(n2801) );
  clknd2d1_hd U544 ( .A(state[0]), .B(n2942), .Y(n2926) );
  clknd2d1_hd U545 ( .A(z_m[19]), .B(z_m[20]), .Y(n2669) );
  clknd2d1_hd U546 ( .A(n2275), .B(n2889), .Y(n2742) );
  clknd2d1_hd U547 ( .A(n2273), .B(n2889), .Y(n2790) );
  clknd2d1_hd U548 ( .A(n2405), .B(n2947), .Y(n2408) );
  clknd2d1_hd U549 ( .A(n2840), .B(n2838), .Y(n2857) );
  clknd2d1_hd U550 ( .A(b_e[2]), .B(n2908), .Y(n2897) );
  clknd2d1_hd U551 ( .A(n2909), .B(n2898), .Y(n2896) );
  clknd2d1_hd U552 ( .A(n2824), .B(n2800), .Y(n2809) );
  clknd2d1_hd U553 ( .A(n2816), .B(n2812), .Y(n2860) );
  clknd2d1_hd U554 ( .A(n2890), .B(b[28]), .Y(n2883) );
  clknd2d1_hd U555 ( .A(n2405), .B(n2936), .Y(n2940) );
  clknd2d1_hd U556 ( .A(state[2]), .B(n2962), .Y(n2944) );
  clknd2d1_hd U557 ( .A(N41), .B(n2961), .Y(n2963) );
  clknd2d1_hd U558 ( .A(n2660), .B(n2650), .Y(n2641) );
  clknd2d1_hd U559 ( .A(z_m[0]), .B(n2660), .Y(n2633) );
  clknd2d1_hd U560 ( .A(n2646), .B(n2641), .Y(n2636) );
  clknd2d1_hd U561 ( .A(n2609), .B(n2660), .Y(n2616) );
  clknd2d1_hd U562 ( .A(n2585), .B(n2660), .Y(n2592) );
  clknd2d1_hd U563 ( .A(z_m[21]), .B(n2670), .Y(n2662) );
  clknd2d1_hd U564 ( .A(n2676), .B(sum[27]), .Y(n2674) );
  clknd2d1_hd U565 ( .A(n2562), .B(n2660), .Y(n2568) );
  clknd2d1_hd U566 ( .A(n2534), .B(n2660), .Y(n2541) );
  clknd2d1_hd U567 ( .A(z_m[15]), .B(z_m[16]), .Y(n2548) );
  clknd2d1_hd U568 ( .A(n2515), .B(n2530), .Y(n2663) );
  clknd2d1_hd U569 ( .A(n2803), .B(n2874), .Y(n2443) );
  clknd2d1_hd U570 ( .A(a_e[0]), .B(b_e[0]), .Y(n2484) );
  clknd2d1_hd U571 ( .A(n2477), .B(n2472), .Y(n2471) );
  clknd2d1_hd U572 ( .A(n2463), .B(n2459), .Y(n2458) );
  clknd2d1_hd U573 ( .A(a_e[7]), .B(b_e[7]), .Y(n2438) );
  clknd2d1_hd U574 ( .A(n2449), .B(n2445), .Y(n2444) );
  clknd2d1_hd U575 ( .A(n2488), .B(n2435), .Y(n2487) );
  ivd1_hd U576 ( .A(b_m[1]), .Y(n2743) );
  clknd2d1_hd U577 ( .A(n2359), .B(n1891), .Y(n2351) );
  ivd1_hd U578 ( .A(b_m[2]), .Y(n2741) );
  clknd2d1_hd U579 ( .A(n2503), .B(n2428), .Y(n2435) );
  clknd2d1_hd U580 ( .A(n2426), .B(n2425), .Y(n2429) );
  nid1_hd U581 ( .A(n2498), .Y(n2270) );
  ivd2_hd U582 ( .A(n2351), .Y(n2356) );
  ivd2_hd U583 ( .A(n2357), .Y(n1891) );
  clknd2d1_hd U584 ( .A(n2324), .B(a_m[26]), .Y(n2325) );
  nr2d1_hd U585 ( .A(n2324), .B(a_m[26]), .Y(n2326) );
  ivd4_hd U586 ( .A(n2359), .Y(n2269) );
  clknd2d1_hd U587 ( .A(state[1]), .B(n2947), .Y(n2923) );
  clknd2d1_hd U588 ( .A(a[23]), .B(a[24]), .Y(n2851) );
  clknd2d1_hd U589 ( .A(n2839), .B(n2857), .Y(n2849) );
  clknd2d1_hd U590 ( .A(a_e[3]), .B(n2833), .Y(n2831) );
  clknd2d1_hd U591 ( .A(n2842), .B(a[26]), .Y(n2835) );
  clknd2d1_hd U592 ( .A(b[23]), .B(b[24]), .Y(n2914) );
  clknd2d1_hd U593 ( .A(n2909), .B(n2912), .Y(n2910) );
  clknd2d1_hd U594 ( .A(a_e[5]), .B(n2819), .Y(n2818) );
  clknd2d1_hd U595 ( .A(n2839), .B(n2889), .Y(n2859) );
  clknd2d1_hd U596 ( .A(a_e[4]), .B(a_e[3]), .Y(n2799) );
  clknd2d1_hd U597 ( .A(n2826), .B(a[28]), .Y(n2820) );
  clknd2d1_hd U598 ( .A(n2903), .B(b[26]), .Y(n2900) );
  clknd2d1_hd U599 ( .A(n2899), .B(n2896), .Y(n2893) );
  clknd2d1_hd U600 ( .A(n2505), .B(n2504), .Y(n393) );
  clknd2d1_hd U601 ( .A(b[30]), .B(n2868), .Y(n2873) );
  clknd2d1_hd U602 ( .A(a_e[0]), .B(n2855), .Y(n2856) );
  clknd2d1_hd U603 ( .A(n2279), .B(n2806), .Y(n2811) );
  clknd2d1_hd U604 ( .A(b_e[5]), .B(n2874), .Y(n2880) );
  clknd2d1_hd U605 ( .A(n2883), .B(n2875), .Y(n2876) );
  clknd2d1_hd U606 ( .A(n2661), .B(n2641), .Y(n2643) );
  clknd2d1_hd U607 ( .A(n2696), .B(n2695), .Y(n428) );
  clknd2d1_hd U608 ( .A(DP_OP_154J4_137_6175_n2), .B(n2694), .Y(n2692) );
  clknd2d1_hd U609 ( .A(n2653), .B(z_m[14]), .Y(n2557) );
  clknd2d1_hd U610 ( .A(n2675), .B(n2508), .Y(n1222) );
  clknd2d1_hd U611 ( .A(n2653), .B(z_m[15]), .Y(n2550) );
  clknd2d1_hd U612 ( .A(n2486), .B(n2441), .Y(n362) );
  clknd2d1_hd U613 ( .A(n2493), .B(n2492), .Y(n2494) );
  clknd2d1_hd U614 ( .A(n2913), .B(n2910), .Y(n2906) );
  clknd2d1_hd U615 ( .A(n2820), .B(n2813), .Y(n2815) );
  clknd2d1_hd U616 ( .A(n2909), .B(n2888), .Y(n2895) );
  oa22ad1_hd U617 ( .A(n2323), .B(b_m[25]), .C(n2322), .D(a_m[25]), .Y(n2324)
         );
  ivd1_hd U618 ( .A(b_m[23]), .Y(n2700) );
  ivd1_hd U619 ( .A(b_m[3]), .Y(n2740) );
  ivd1_hd U620 ( .A(b_m[21]), .Y(n2704) );
  ivd1_hd U621 ( .A(a_m[24]), .Y(n2746) );
  nr2d1_hd U622 ( .A(n2322), .B(a_m[25]), .Y(n2323) );
  ao22d1_hd U623 ( .A(b_m[24]), .B(n2746), .C(n2321), .D(n2320), .Y(n2322) );
  oa22d1_hd U624 ( .A(a_m[23]), .B(n2700), .C(n2319), .D(n2318), .Y(n2320) );
  nr2d1_hd U625 ( .A(n2317), .B(n2316), .Y(n2319) );
  ao21d1_hd U626 ( .A(n2704), .B(a_m[21]), .C(n2315), .Y(n2316) );
  ivd3_hd U627 ( .A(n1284), .Y(n2268) );
  oa22d2_hd U628 ( .A(n2432), .B(n2416), .C(b_s), .D(a_s), .Y(n2357) );
  xo2d1_hd U629 ( .A(n1891), .B(DP_OP_43J4_124_6938_n1), .Y(N337) );
  oa211d8_hd U630 ( .A(b_m[26]), .B(n2326), .C(n1891), .D(n2325), .Y(n2359) );
  nid4_hd U631 ( .A(n27), .Y(n2282) );
  ad3d1_hd U632 ( .A(n2847), .B(n2841), .C(n2840), .Y(n2845) );
  scg6d1_hd U633 ( .A(b_m[17]), .B(n2310), .C(n2760), .Y(n2308) );
  scg6d1_hd U634 ( .A(b_m[10]), .B(n2299), .C(n2774), .Y(n2297) );
  scg9d1_hd U635 ( .A(n2958), .B(n2515), .C(n2528), .Y(n2519) );
  scg9d1_hd U636 ( .A(n2940), .B(n2406), .C(n2280), .Y(n2951) );
  ad3d1_hd U637 ( .A(n2960), .B(n2276), .C(n2958), .Y(n2964) );
  scg6d1_hd U638 ( .A(b_m[6]), .B(n2292), .C(n2782), .Y(n2290) );
  ivd2_hd U639 ( .A(n2674), .Y(n2648) );
  scg10d1_hd U640 ( .A(n2415), .B(n2414), .C(n2413), .D(n2412), .Y(n2492) );
  ad2d1_hd U641 ( .A(n2930), .B(n2511), .Y(n2507) );
  ivd2_hd U642 ( .A(n1285), .Y(n2280) );
  or2d1_hd U643 ( .A(n2944), .B(n2667), .Y(n1284) );
  or2d1_hd U644 ( .A(state[2]), .B(n2962), .Y(n2922) );
  ivd1_hd U645 ( .A(b_m[0]), .Y(n2744) );
  nr2ad1_hd U646 ( .A(n2958), .B(n2635), .Y(n2660) );
  nr2d2_hd U647 ( .A(n2489), .B(n2924), .Y(n2499) );
  nr2ad1_hd U648 ( .A(n2678), .B(n2690), .Y(n2693) );
  nr2ad1_hd U649 ( .A(n2960), .B(n2635), .Y(n2642) );
  nr2ad1_hd U650 ( .A(n2923), .B(n2944), .Y(n1291) );
  oa22ad1_hd U651 ( .A(n2296), .B(a_m[9]), .C(n2295), .D(b_m[9]), .Y(n2299) );
  oa22ad1_hd U652 ( .A(n2289), .B(a_m[5]), .C(n2288), .D(b_m[5]), .Y(n2292) );
  ivd1_hd U653 ( .A(b_m[4]), .Y(n2738) );
  ivd1_hd U654 ( .A(a_m[4]), .Y(n2786) );
  ivd1_hd U655 ( .A(a_m[3]), .Y(n2788) );
  ad3d1_hd U656 ( .A(n2921), .B(i_AB_STB), .C(o_AB_ACK), .Y(n27) );
  nid2_hd U657 ( .A(n2959), .Y(n2276) );
  ivd1_hd U658 ( .A(n2660), .Y(n2634) );
  ivd1_hd U659 ( .A(n2688), .Y(n2690) );
  ivd1_hd U660 ( .A(n2796), .Y(n2274) );
  ivd1_hd U661 ( .A(n2940), .Y(n2889) );
  ivd1_hd U662 ( .A(b_m[7]), .Y(n2732) );
  ivd1_hd U663 ( .A(b_m[8]), .Y(n2730) );
  nid2_hd U664 ( .A(n2500), .Y(n2271) );
  ivd1_hd U665 ( .A(n2653), .Y(n2661) );
  nr2d1_hd U666 ( .A(n2934), .B(n2635), .Y(n2653) );
  ivd1_hd U667 ( .A(n2677), .Y(n2958) );
  nid2_hd U668 ( .A(n2647), .Y(n2272) );
  ivd1_hd U669 ( .A(n2642), .Y(n2649) );
  ivd1_hd U670 ( .A(n2676), .Y(n2508) );
  ivd1_hd U671 ( .A(n2280), .Y(n2277) );
  ivd2_hd U672 ( .A(n2790), .Y(n2793) );
  nr2d1_hd U673 ( .A(n2922), .B(n2667), .Y(n2677) );
  ivd2_hd U674 ( .A(n2951), .Y(n2275) );
  ivd2_hd U675 ( .A(n2274), .Y(n2273) );
  oa21d1_hd U676 ( .A(n2927), .B(n2928), .C(n2280), .Y(n2796) );
  nr2d1_hd U677 ( .A(n2418), .B(n2925), .Y(n2946) );
  ivd1_hd U678 ( .A(n1895), .Y(n2925) );
  ivd1_hd U679 ( .A(n2280), .Y(n2279) );
  ivd1_hd U680 ( .A(b_m[15]), .Y(n2716) );
  ivd1_hd U681 ( .A(b_m[14]), .Y(n2718) );
  ivd1_hd U682 ( .A(b_m[13]), .Y(n2720) );
  ivd1_hd U683 ( .A(a_m[12]), .Y(n2770) );
  ivd1_hd U684 ( .A(b_m[16]), .Y(n2714) );
  ivd1_hd U685 ( .A(b_m[18]), .Y(n2710) );
  ivd1_hd U686 ( .A(b_m[24]), .Y(n2698) );
  nid2_hd U687 ( .A(n509), .Y(n2281) );
  ivd1_hd U688 ( .A(n2488), .Y(n2924) );
  ivd2_hd U689 ( .A(n2742), .Y(n2949) );
  ivd1_hd U690 ( .A(n2495), .Y(n2479) );
  nr2d1_hd U691 ( .A(n2926), .B(n2922), .Y(n2488) );
  ivd1_hd U692 ( .A(n2511), .Y(n2960) );
  ivd2_hd U693 ( .A(n2280), .Y(n2278) );
  ivd1_hd U694 ( .A(n1291), .Y(n2934) );
  nr2d1_hd U695 ( .A(n2926), .B(n2944), .Y(n2676) );
  nr2bd1_hd U696 ( .AN(n2936), .B(n2944), .Y(n2511) );
  nr2bd1_hd U697 ( .AN(z_e[1]), .B(n2501), .Y(n2503) );
  ivd1_hd U698 ( .A(n2861), .Y(n2853) );
  ivd1_hd U699 ( .A(n2909), .Y(n2954) );
  nr2d1_hd U700 ( .A(n2919), .B(n2940), .Y(n2909) );
  ao21d1_hd U701 ( .A(n2863), .B(n2946), .C(n2275), .Y(n2919) );
  ivd1_hd U702 ( .A(n2855), .Y(n2839) );
  ao21d1_hd U703 ( .A(n2797), .B(n2946), .C(n2273), .Y(n2855) );
  ivd1_hd U704 ( .A(b_e[7]), .Y(n2869) );
  ivd1_hd U705 ( .A(a_e[6]), .Y(n2803) );
  ivd1_hd U706 ( .A(a_e[5]), .Y(n2823) );
  ivd1_hd U707 ( .A(b_e[1]), .Y(n2912) );
  nr2d1_hd U708 ( .A(n2942), .B(n2408), .Y(n1895) );
  ivd1_hd U709 ( .A(b_e[8]), .Y(n2867) );
  ivd1_hd U710 ( .A(n2450), .Y(n2411) );
  ivd1_hd U711 ( .A(n2491), .Y(n2415) );
  ivd1_hd U712 ( .A(a_e[4]), .Y(n2802) );
  ivd1_hd U713 ( .A(a_e[0]), .Y(n2838) );
  nr2d1_hd U714 ( .A(n2947), .B(n2942), .Y(n2936) );
  ivd1_hd U715 ( .A(state[0]), .Y(n2947) );
  nr2bd1_hd U716 ( .AN(n2405), .B(n2926), .Y(n1285) );
  ivd1_hd U717 ( .A(state[1]), .Y(n2942) );
  ivd1_hd U718 ( .A(a_m[23]), .Y(n2748) );
  ivd1_hd U719 ( .A(a_m[22]), .Y(n2750) );
  ivd1_hd U720 ( .A(b_m[19]), .Y(n2708) );
  ivd1_hd U721 ( .A(b_m[20]), .Y(n2706) );
  ivd1_hd U722 ( .A(a_m[20]), .Y(n2754) );
  ivd1_hd U723 ( .A(b_m[22]), .Y(n2702) );
  ivd1_hd U724 ( .A(n2946), .Y(n2407) );
  ivd1_hd U725 ( .A(z_m[1]), .Y(n2650) );
  ivd1_hd U726 ( .A(z_m[14]), .Y(n2567) );
  ivd1_hd U727 ( .A(n2635), .Y(n2656) );
  nr4d1_hd U728 ( .A(n2491), .B(n2411), .C(n2410), .D(n2925), .Y(n2498) );
  oa21d1_hd U729 ( .A(n2935), .B(n2934), .C(n2933), .Y(n2961) );
  nr2d1_hd U730 ( .A(n2923), .B(n2922), .Y(n509) );
  ivd1_hd U731 ( .A(z_m[19]), .Y(n2539) );
  nr2d1_hd U732 ( .A(n2276), .B(n2925), .Y(n2495) );
  ao22d1_hd U733 ( .A(n2489), .B(n2488), .C(n1895), .D(n2434), .Y(n2486) );
  scg20d1_hd U734 ( .A(z_e[7]), .B(z_e[8]), .C(z_e[9]), .Y(n2489) );
  ivd1_hd U735 ( .A(z_m[22]), .Y(n2659) );
  ivd1_hd U736 ( .A(round_bit), .Y(n2512) );
  ivd1_hd U737 ( .A(z_m[0]), .Y(n2657) );
  ivd1_hd U738 ( .A(n2916), .Y(n2956) );
  ivd1_hd U739 ( .A(z_m[12]), .Y(n2578) );
  ivd1_hd U740 ( .A(z_m[11]), .Y(n2590) );
  ivd1_hd U741 ( .A(z_m[7]), .Y(n2614) );
  ivd1_hd U742 ( .A(z_m[8]), .Y(n2602) );
  ivd1_hd U743 ( .A(z_m[3]), .Y(n2640) );
  ivd1_hd U744 ( .A(z_m[4]), .Y(n2626) );
  ivd1_hd U745 ( .A(z_m[23]), .Y(n2670) );
  ivd1_hd U746 ( .A(state[3]), .Y(n2962) );
  ivd1_hd U747 ( .A(z_e[2]), .Y(n2472) );
  ivd1_hd U748 ( .A(z_e[0]), .Y(n2689) );
  nr2d1_hd U749 ( .A(n2919), .B(n2925), .Y(n2916) );
  ivd1_hd U750 ( .A(n2859), .Y(n2840) );
  ivd1_hd U751 ( .A(a_e[7]), .Y(n2807) );
  ivd1_hd U752 ( .A(b_e[3]), .Y(n2898) );
  nr4d1_hd U753 ( .A(n2404), .B(n2386), .C(n2387), .D(n2385), .Y(n2927) );
  ivd1_hd U754 ( .A(a_e[2]), .Y(n2847) );
  nr2d1_hd U755 ( .A(b_e[9]), .B(n2380), .Y(n2404) );
  scg13d1_hd U756 ( .A(n2434), .B(n2411), .C(n2410), .Y(n2418) );
  ivd1_hd U757 ( .A(b_e[0]), .Y(n2911) );
  ivd1_hd U758 ( .A(b_e[5]), .Y(n2886) );
  ivd1_hd U759 ( .A(b_e[6]), .Y(n2874) );
  ivd1_hd U760 ( .A(a_e[3]), .Y(n2832) );
  ivd1_hd U761 ( .A(a_e[9]), .Y(n2380) );
  ivd1_hd U762 ( .A(a_e[8]), .Y(n2805) );
  ivd1_hd U763 ( .A(a_e[1]), .Y(n2798) );
  nr2d1_hd U764 ( .A(state[2]), .B(state[3]), .Y(n2405) );
  ivd1_hd U765 ( .A(a[30]), .Y(n2812) );
  ivd1_hd U766 ( .A(a_m[0]), .Y(n2792) );
  ivd1_hd U767 ( .A(a_m[1]), .Y(n2791) );
  ivd1_hd U768 ( .A(a_m[2]), .Y(n2789) );
  ivd1_hd U769 ( .A(b_m[5]), .Y(n2736) );
  ivd1_hd U770 ( .A(a_m[5]), .Y(n2784) );
  ivd1_hd U771 ( .A(b_m[6]), .Y(n2734) );
  ivd1_hd U772 ( .A(b_m[9]), .Y(n2728) );
  ivd1_hd U773 ( .A(a_m[9]), .Y(n2776) );
  ivd1_hd U774 ( .A(b_m[10]), .Y(n2726) );
  ivd1_hd U775 ( .A(b_m[12]), .Y(n2722) );
  ivd1_hd U776 ( .A(a_m[14]), .Y(n2766) );
  ivd1_hd U777 ( .A(b_m[17]), .Y(n2712) );
  ivd1_hd U778 ( .A(a_m[18]), .Y(n2758) );
  ivd1_hd U779 ( .A(a_m[21]), .Y(n2752) );
  ivd1_hd U780 ( .A(b_m[25]), .Y(n2952) );
  ivd1_hd U781 ( .A(a_m[19]), .Y(n2756) );
  ivd1_hd U782 ( .A(a_m[17]), .Y(n2760) );
  ivd1_hd U783 ( .A(a_m[13]), .Y(n2768) );
  ivd1_hd U784 ( .A(a_m[10]), .Y(n2774) );
  ivd1_hd U785 ( .A(b_m[11]), .Y(n2724) );
  ivd1_hd U786 ( .A(a_m[6]), .Y(n2782) );
  ivd1_hd U787 ( .A(a_m[8]), .Y(n2778) );
  ivd1_hd U788 ( .A(a_m[7]), .Y(n2780) );
  ivd1_hd U789 ( .A(a_m[11]), .Y(n2772) );
  ivd1_hd U790 ( .A(a_m[16]), .Y(n2762) );
  ivd1_hd U791 ( .A(a_m[15]), .Y(n2764) );
  ivd1_hd U792 ( .A(b_s), .Y(n2416) );
  ivd1_hd U793 ( .A(a_s), .Y(n2432) );
  nr2d1_hd U794 ( .A(state[1]), .B(n2408), .Y(n2921) );
  nr2d1_hd U795 ( .A(sum[27]), .B(n2508), .Y(n2647) );
  nd2bd1_hd U796 ( .AN(b[30]), .B(n2877), .Y(n2955) );
  nr2d1_hd U797 ( .A(n2925), .B(n2855), .Y(n2861) );
  nd2bd1_hd U798 ( .AN(n2404), .B(n2403), .Y(n2406) );
  ivd1_hd U799 ( .A(b_e[9]), .Y(n2400) );
  ivd1_hd U800 ( .A(a_m[25]), .Y(n2795) );
  oa22d1_hd U801 ( .A(a_m[21]), .B(n2704), .C(a_m[22]), .D(n2702), .Y(n2317)
         );
  ao22d1_hd U802 ( .A(a_m[20]), .B(n2706), .C(a_m[19]), .D(n2708), .Y(n2314)
         );
  ao22d1_hd U803 ( .A(b_m[15]), .B(n2764), .C(b_m[16]), .D(n2762), .Y(n2307)
         );
  ao22d1_hd U804 ( .A(b_m[11]), .B(n2772), .C(b_m[12]), .D(n2770), .Y(n2302)
         );
  ao22d1_hd U805 ( .A(b_m[7]), .B(n2780), .C(b_m[8]), .D(n2778), .Y(n2294) );
  ao22d1_hd U806 ( .A(b_m[3]), .B(n2788), .C(b_m[4]), .D(n2786), .Y(n2287) );
  ao211d1_hd U807 ( .A(a_m[1]), .B(n2743), .C(a_m[0]), .D(n2744), .Y(n2285) );
  oa22d1_hd U808 ( .A(a_m[1]), .B(n2743), .C(a_m[2]), .D(n2741), .Y(n2284) );
  ao22d1_hd U809 ( .A(a_m[3]), .B(n2740), .C(a_m[2]), .D(n2741), .Y(n2283) );
  oa21d1_hd U810 ( .A(n2285), .B(n2284), .C(n2283), .Y(n2286) );
  ao22d1_hd U811 ( .A(a_m[4]), .B(n2738), .C(n2287), .D(n2286), .Y(n2288) );
  nr2d1_hd U812 ( .A(n2288), .B(b_m[5]), .Y(n2289) );
  oa211d1_hd U813 ( .A(b_m[6]), .B(n2292), .C(n2291), .D(n2290), .Y(n2293) );
  ao22d1_hd U814 ( .A(a_m[8]), .B(n2730), .C(n2294), .D(n2293), .Y(n2295) );
  nr2d1_hd U815 ( .A(n2295), .B(b_m[9]), .Y(n2296) );
  oa211d1_hd U816 ( .A(b_m[10]), .B(n2299), .C(n2298), .D(n2297), .Y(n2301) );
  oa22d1_hd U817 ( .A(b_m[13]), .B(n2768), .C(b_m[12]), .D(n2770), .Y(n2300)
         );
  ao21d1_hd U818 ( .A(n2302), .B(n2301), .C(n2300), .Y(n2305) );
  oa22d1_hd U819 ( .A(a_m[13]), .B(n2720), .C(a_m[14]), .D(n2718), .Y(n2304)
         );
  ao22d1_hd U820 ( .A(a_m[15]), .B(n2716), .C(a_m[14]), .D(n2718), .Y(n2303)
         );
  oa21d1_hd U821 ( .A(n2305), .B(n2304), .C(n2303), .Y(n2306) );
  ao22d1_hd U822 ( .A(a_m[16]), .B(n2714), .C(n2307), .D(n2306), .Y(n2310) );
  oa211d1_hd U823 ( .A(b_m[17]), .B(n2310), .C(n2309), .D(n2308), .Y(n2312) );
  oa211d1_hd U824 ( .A(a_m[18]), .B(n2710), .C(n2312), .D(n2311), .Y(n2313) );
  ao22d1_hd U825 ( .A(b_m[20]), .B(n2754), .C(n2314), .D(n2313), .Y(n2315) );
  oa22d1_hd U826 ( .A(b_m[22]), .B(n2750), .C(b_m[23]), .D(n2748), .Y(n2318)
         );
  ao22d1_hd U827 ( .A(n2269), .B(n2744), .C(n2792), .D(n2359), .Y(C2_Z_0) );
  ao22d1_hd U828 ( .A(n2269), .B(n2743), .C(n2791), .D(n2359), .Y(C2_Z_1) );
  ao22d1_hd U829 ( .A(n2269), .B(n2726), .C(n2774), .D(n2359), .Y(C2_Z_10) );
  ao22d1_hd U830 ( .A(n2269), .B(n2724), .C(n2772), .D(n2359), .Y(C2_Z_11) );
  ao22d1_hd U831 ( .A(n2269), .B(n2722), .C(n2770), .D(n2359), .Y(C2_Z_12) );
  ao22d1_hd U832 ( .A(n2269), .B(n2720), .C(n2768), .D(n2359), .Y(C2_Z_13) );
  ao22d1_hd U833 ( .A(n2269), .B(n2718), .C(n2766), .D(n2359), .Y(C2_Z_14) );
  ao22d1_hd U834 ( .A(n2269), .B(n2716), .C(n2764), .D(n2359), .Y(C2_Z_15) );
  ao22d1_hd U835 ( .A(n2269), .B(n2714), .C(n2762), .D(n2359), .Y(C2_Z_16) );
  ao22d1_hd U836 ( .A(n2269), .B(n2712), .C(n2760), .D(n2359), .Y(C2_Z_17) );
  ao22d1_hd U837 ( .A(n2269), .B(n2710), .C(n2758), .D(n2359), .Y(C2_Z_18) );
  ao22d1_hd U838 ( .A(n2269), .B(n2708), .C(n2756), .D(n2359), .Y(C2_Z_19) );
  ao22d1_hd U839 ( .A(n2269), .B(n2741), .C(n2789), .D(n2359), .Y(C2_Z_2) );
  ao22d1_hd U840 ( .A(n2269), .B(n2706), .C(n2754), .D(n2359), .Y(C2_Z_20) );
  ao22d1_hd U841 ( .A(n2269), .B(n2704), .C(n2752), .D(n2359), .Y(C2_Z_21) );
  ao22d1_hd U842 ( .A(n2269), .B(n2702), .C(n2750), .D(n2359), .Y(C2_Z_22) );
  ao22d1_hd U843 ( .A(n2269), .B(n2700), .C(n2748), .D(n2359), .Y(C2_Z_23) );
  ao22d1_hd U844 ( .A(n2269), .B(n2698), .C(n2746), .D(n2359), .Y(C2_Z_24) );
  ao22d1_hd U845 ( .A(n2269), .B(n2952), .C(n2795), .D(n2359), .Y(C2_Z_25) );
  ivd1_hd U846 ( .A(b_m[26]), .Y(n2328) );
  ivd1_hd U847 ( .A(a_m[26]), .Y(n2327) );
  oa21d1_hd U848 ( .A(n2328), .B(n2357), .C(n2327), .Y(C2_Z_26) );
  ao22d1_hd U849 ( .A(n2269), .B(n2740), .C(n2788), .D(n2359), .Y(C2_Z_3) );
  ao22d1_hd U850 ( .A(n2269), .B(n2738), .C(n2786), .D(n2359), .Y(C2_Z_4) );
  ao22d1_hd U851 ( .A(n2269), .B(n2736), .C(n2784), .D(n2359), .Y(C2_Z_5) );
  ao22d1_hd U852 ( .A(n2269), .B(n2734), .C(n2782), .D(n2359), .Y(C2_Z_6) );
  ao22d1_hd U853 ( .A(n2269), .B(n2732), .C(n2780), .D(n2359), .Y(C2_Z_7) );
  ao22d1_hd U854 ( .A(n2269), .B(n2730), .C(n2778), .D(n2359), .Y(C2_Z_8) );
  ao22d1_hd U855 ( .A(n2269), .B(n2728), .C(n2776), .D(n2359), .Y(C2_Z_9) );
  nr2d1_hd U856 ( .A(n2328), .B(n2327), .Y(n2329) );
  ao22d1_hd U857 ( .A(n1891), .B(n2329), .C(n2328), .D(n2357), .Y(
        DP_OP_43J4_124_6938_n32) );
  ao22d1_hd U858 ( .A(b_m[25]), .B(n2357), .C(n2356), .D(n2952), .Y(n2330) );
  oa21d1_hd U859 ( .A(a_m[25]), .B(n2359), .C(n2330), .Y(
        DP_OP_43J4_124_6938_n33) );
  ao22d1_hd U860 ( .A(n2269), .B(n2746), .C(n2356), .D(n2698), .Y(n2331) );
  oa21d1_hd U861 ( .A(n1891), .B(n2698), .C(n2331), .Y(DP_OP_43J4_124_6938_n34) );
  ao22d1_hd U862 ( .A(n2269), .B(n2748), .C(n2356), .D(n2700), .Y(n2332) );
  oa21d1_hd U863 ( .A(n1891), .B(n2700), .C(n2332), .Y(DP_OP_43J4_124_6938_n35) );
  ao22d1_hd U864 ( .A(n2269), .B(n2750), .C(n2356), .D(n2702), .Y(n2333) );
  oa21d1_hd U865 ( .A(n1891), .B(n2702), .C(n2333), .Y(DP_OP_43J4_124_6938_n36) );
  ao22d1_hd U866 ( .A(b_m[21]), .B(n2357), .C(n2356), .D(n2704), .Y(n2334) );
  oa21d1_hd U867 ( .A(a_m[21]), .B(n2359), .C(n2334), .Y(
        DP_OP_43J4_124_6938_n37) );
  ao22d1_hd U868 ( .A(n2269), .B(n2754), .C(n2356), .D(n2706), .Y(n2335) );
  oa21d1_hd U869 ( .A(n1891), .B(n2706), .C(n2335), .Y(DP_OP_43J4_124_6938_n38) );
  ao22d1_hd U870 ( .A(n2269), .B(n2756), .C(n2356), .D(n2708), .Y(n2336) );
  oa21d1_hd U871 ( .A(n1891), .B(n2708), .C(n2336), .Y(DP_OP_43J4_124_6938_n39) );
  ao22d1_hd U872 ( .A(b_m[18]), .B(n2357), .C(n2356), .D(n2710), .Y(n2337) );
  oa21d1_hd U873 ( .A(a_m[18]), .B(n2359), .C(n2337), .Y(
        DP_OP_43J4_124_6938_n40) );
  ao22d1_hd U874 ( .A(b_m[17]), .B(n2357), .C(n2356), .D(n2712), .Y(n2338) );
  oa21d1_hd U875 ( .A(a_m[17]), .B(n2359), .C(n2338), .Y(
        DP_OP_43J4_124_6938_n41) );
  ao22d1_hd U876 ( .A(n2269), .B(n2762), .C(n2356), .D(n2714), .Y(n2339) );
  oa21d1_hd U877 ( .A(n1891), .B(n2714), .C(n2339), .Y(DP_OP_43J4_124_6938_n42) );
  ao22d1_hd U878 ( .A(n2269), .B(n2764), .C(n2356), .D(n2716), .Y(n2340) );
  oa21d1_hd U879 ( .A(n1891), .B(n2716), .C(n2340), .Y(DP_OP_43J4_124_6938_n43) );
  ao22d1_hd U880 ( .A(b_m[14]), .B(n2357), .C(n2356), .D(n2718), .Y(n2341) );
  oa21d1_hd U881 ( .A(a_m[14]), .B(n2359), .C(n2341), .Y(
        DP_OP_43J4_124_6938_n44) );
  ao22d1_hd U882 ( .A(n2269), .B(n2768), .C(n2356), .D(n2720), .Y(n2342) );
  oa21d1_hd U883 ( .A(n1891), .B(n2720), .C(n2342), .Y(DP_OP_43J4_124_6938_n45) );
  ao22d1_hd U884 ( .A(n2269), .B(n2770), .C(b_m[12]), .D(n2357), .Y(n2343) );
  oa21d1_hd U885 ( .A(b_m[12]), .B(n2351), .C(n2343), .Y(
        DP_OP_43J4_124_6938_n46) );
  ao22d1_hd U886 ( .A(n2269), .B(n2772), .C(n2356), .D(n2724), .Y(n2344) );
  oa21d1_hd U887 ( .A(n1891), .B(n2724), .C(n2344), .Y(DP_OP_43J4_124_6938_n47) );
  ao22d1_hd U888 ( .A(n2269), .B(n2774), .C(b_m[10]), .D(n2357), .Y(n2345) );
  oa21d1_hd U889 ( .A(b_m[10]), .B(n2351), .C(n2345), .Y(
        DP_OP_43J4_124_6938_n48) );
  ao22d1_hd U890 ( .A(n2269), .B(n2776), .C(b_m[9]), .D(n2357), .Y(n2346) );
  oa21d1_hd U891 ( .A(b_m[9]), .B(n2351), .C(n2346), .Y(
        DP_OP_43J4_124_6938_n49) );
  ao22d1_hd U892 ( .A(n2269), .B(n2778), .C(n2356), .D(n2730), .Y(n2347) );
  oa21d1_hd U893 ( .A(n1891), .B(n2730), .C(n2347), .Y(DP_OP_43J4_124_6938_n50) );
  ao22d1_hd U894 ( .A(n2269), .B(n2780), .C(n2356), .D(n2732), .Y(n2348) );
  oa21d1_hd U895 ( .A(n1891), .B(n2732), .C(n2348), .Y(DP_OP_43J4_124_6938_n51) );
  ao22d1_hd U896 ( .A(n2269), .B(n2782), .C(b_m[6]), .D(n2357), .Y(n2349) );
  oa21d1_hd U897 ( .A(b_m[6]), .B(n2351), .C(n2349), .Y(
        DP_OP_43J4_124_6938_n52) );
  ao22d1_hd U898 ( .A(n2269), .B(n2784), .C(b_m[5]), .D(n2357), .Y(n2350) );
  oa21d1_hd U899 ( .A(b_m[5]), .B(n2351), .C(n2350), .Y(
        DP_OP_43J4_124_6938_n53) );
  ao22d1_hd U900 ( .A(n2269), .B(n2786), .C(n2356), .D(n2738), .Y(n2352) );
  oa21d1_hd U901 ( .A(n1891), .B(n2738), .C(n2352), .Y(DP_OP_43J4_124_6938_n54) );
  ao22d1_hd U902 ( .A(n2269), .B(n2788), .C(n2356), .D(n2740), .Y(n2353) );
  oa21d1_hd U903 ( .A(n1891), .B(n2740), .C(n2353), .Y(DP_OP_43J4_124_6938_n55) );
  ao22d1_hd U904 ( .A(b_m[2]), .B(n2357), .C(n2356), .D(n2741), .Y(n2354) );
  oa21d1_hd U905 ( .A(a_m[2]), .B(n2359), .C(n2354), .Y(
        DP_OP_43J4_124_6938_n56) );
  ao22d1_hd U906 ( .A(b_m[1]), .B(n2357), .C(n2356), .D(n2743), .Y(n2355) );
  oa21d1_hd U907 ( .A(a_m[1]), .B(n2359), .C(n2355), .Y(
        DP_OP_43J4_124_6938_n57) );
  ao22d1_hd U908 ( .A(b_m[0]), .B(n2357), .C(n2356), .D(n2744), .Y(n2358) );
  oa21d1_hd U909 ( .A(a_m[0]), .B(n2359), .C(n2358), .Y(
        DP_OP_43J4_124_6938_n58) );
  ao22d1_hd U910 ( .A(n2269), .B(n2416), .C(n2432), .D(n2359), .Y(N338) );
  nr4d1_hd U911 ( .A(a_e[6]), .B(a_e[2]), .C(a_e[1]), .D(a_e[5]), .Y(n2360) );
  nd4d1_hd U912 ( .A(a_e[7]), .B(n2360), .C(n2802), .D(n2832), .Y(n2361) );
  nr4d1_hd U913 ( .A(n2805), .B(n2838), .C(n2380), .D(n2361), .Y(n2797) );
  nr4d1_hd U914 ( .A(a_e[8]), .B(a_e[0]), .C(a_e[9]), .D(n2361), .Y(n2491) );
  nr4d1_hd U915 ( .A(b_e[2]), .B(b_e[1]), .C(b_e[3]), .D(b_e[4]), .Y(n2362) );
  nd4d1_hd U916 ( .A(b_e[7]), .B(n2362), .C(n2874), .D(n2886), .Y(n2371) );
  nr4d1_hd U917 ( .A(b_e[9]), .B(b_e[8]), .C(b_e[0]), .D(n2371), .Y(n2490) );
  ivd1_hd U918 ( .A(n2490), .Y(n2413) );
  nd4d1_hd U919 ( .A(n2748), .B(n2774), .C(n2792), .D(n2789), .Y(n2370) );
  nr4d1_hd U920 ( .A(a_m[25]), .B(a_m[11]), .C(a_m[12]), .D(a_m[26]), .Y(n2363) );
  nd4d1_hd U921 ( .A(n2363), .B(n2746), .C(n2754), .D(n2750), .Y(n2369) );
  nr4d1_hd U922 ( .A(a_m[13]), .B(a_m[14]), .C(a_m[15]), .D(a_m[16]), .Y(n2367) );
  nr4d1_hd U923 ( .A(a_m[21]), .B(a_m[17]), .C(a_m[18]), .D(a_m[19]), .Y(n2366) );
  nr4d1_hd U924 ( .A(a_m[5]), .B(a_m[1]), .C(a_m[3]), .D(a_m[4]), .Y(n2365) );
  nr4d1_hd U925 ( .A(a_m[9]), .B(a_m[6]), .C(a_m[7]), .D(a_m[8]), .Y(n2364) );
  nd4d1_hd U926 ( .A(n2367), .B(n2366), .C(n2365), .D(n2364), .Y(n2368) );
  nr3d1_hd U927 ( .A(n2370), .B(n2369), .C(n2368), .Y(n2414) );
  nr4d1_hd U928 ( .A(n2371), .B(n2867), .C(n2400), .D(n2911), .Y(n2863) );
  nd4d1_hd U929 ( .A(n2698), .B(n2712), .C(n2722), .D(n2714), .Y(n2379) );
  nr4d1_hd U930 ( .A(b_m[0]), .B(b_m[7]), .C(b_m[14]), .D(b_m[26]), .Y(n2372)
         );
  nd4d1_hd U931 ( .A(n2372), .B(n2700), .C(n2743), .D(n2741), .Y(n2378) );
  nr4d1_hd U932 ( .A(b_m[21]), .B(b_m[13]), .C(b_m[19]), .D(b_m[20]), .Y(n2376) );
  nr4d1_hd U933 ( .A(b_m[25]), .B(b_m[10]), .C(b_m[18]), .D(b_m[22]), .Y(n2375) );
  nr4d1_hd U934 ( .A(b_m[3]), .B(b_m[4]), .C(b_m[11]), .D(b_m[15]), .Y(n2374)
         );
  nr4d1_hd U935 ( .A(b_m[9]), .B(b_m[6]), .C(b_m[5]), .D(b_m[8]), .Y(n2373) );
  nd4d1_hd U936 ( .A(n2376), .B(n2375), .C(n2374), .D(n2373), .Y(n2377) );
  nr3d1_hd U937 ( .A(n2379), .B(n2378), .C(n2377), .Y(n2412) );
  nr2d1_hd U938 ( .A(a_e[1]), .B(n2912), .Y(n2386) );
  ao22d1_hd U939 ( .A(b_e[4]), .B(n2802), .C(b_e[5]), .D(n2823), .Y(n2381) );
  ao22d1_hd U940 ( .A(b_e[2]), .B(n2847), .C(b_e[3]), .D(n2832), .Y(n2388) );
  nr2d1_hd U941 ( .A(n2867), .B(a_e[8]), .Y(n2401) );
  ivd1_hd U942 ( .A(n2401), .Y(n2384) );
  nr2d1_hd U943 ( .A(n2869), .B(a_e[7]), .Y(n2397) );
  ivd1_hd U944 ( .A(n2397), .Y(n2383) );
  nd4d1_hd U945 ( .A(n2388), .B(n2384), .C(n2383), .D(n2382), .Y(n2385) );
  ivd1_hd U946 ( .A(n2387), .Y(n2396) );
  ao211d1_hd U947 ( .A(b_e[1]), .B(n2798), .C(b_e[0]), .D(n2838), .Y(n2390) );
  oa22d1_hd U948 ( .A(b_e[2]), .B(n2847), .C(b_e[1]), .D(n2798), .Y(n2389) );
  oa21d1_hd U949 ( .A(n2390), .B(n2389), .C(n2388), .Y(n2392) );
  oa211d1_hd U950 ( .A(b_e[4]), .B(n2802), .C(n2392), .D(n2391), .Y(n2395) );
  oa22d1_hd U951 ( .A(b_e[6]), .B(n2803), .C(b_e[5]), .D(n2823), .Y(n2393) );
  ao22d1_hd U952 ( .A(n2396), .B(n2395), .C(n2394), .D(n2393), .Y(n2398) );
  oa22d1_hd U953 ( .A(b_e[8]), .B(n2805), .C(n2398), .D(n2397), .Y(n2399) );
  ao21d1_hd U954 ( .A(a_e[7]), .B(n2869), .C(n2399), .Y(n2402) );
  oa22d1_hd U955 ( .A(n2402), .B(n2401), .C(a_e[9]), .D(n2400), .Y(n2403) );
  oa21d1_hd U956 ( .A(n2797), .B(n2407), .C(n2274), .Y(n1) );
  oa21d1_hd U957 ( .A(n2863), .B(n2407), .C(n2951), .Y(n2) );
  scg4d1_hd U958 ( .A(n1291), .B(round_bit), .C(z_m[0]), .D(n2511), .E(n2648), 
        .F(sum[3]), .G(n2272), .H(sum[2]), .Y(n266) );
  oa22d1_hd U959 ( .A(n2490), .B(n2415), .C(n2416), .D(n2450), .Y(n2409) );
  ao21d1_hd U960 ( .A(n1895), .B(n2409), .C(n2270), .Y(n2433) );
  ao21d1_hd U961 ( .A(n2411), .B(n2410), .C(n2490), .Y(n2417) );
  oa21d1_hd U962 ( .A(n2417), .B(n2416), .C(n2492), .Y(n2419) );
  ao21d1_hd U963 ( .A(n1895), .B(n2418), .C(n2488), .Y(n2959) );
  ao22d1_hd U964 ( .A(n1895), .B(n2419), .C(n2276), .D(z[31]), .Y(n2431) );
  ivd1_hd U965 ( .A(z_m[15]), .Y(n2555) );
  ivd1_hd U966 ( .A(z_m[16]), .Y(n2546) );
  ivd1_hd U967 ( .A(z_m[2]), .Y(n2632) );
  nd4d1_hd U968 ( .A(n2555), .B(n2546), .C(n2632), .D(n2626), .Y(n2420) );
  nr4d1_hd U969 ( .A(z_m[0]), .B(z_m[22]), .C(z_m[1]), .D(n2420), .Y(n2426) );
  ivd1_hd U970 ( .A(z_m[9]), .Y(n2591) );
  ivd1_hd U971 ( .A(z_m[10]), .Y(n2584) );
  nd4d1_hd U972 ( .A(n2614), .B(n2591), .C(n2584), .D(n2590), .Y(n2424) );
  ivd1_hd U973 ( .A(z_m[5]), .Y(n2615) );
  ivd1_hd U974 ( .A(z_m[6]), .Y(n2608) );
  nd4d1_hd U975 ( .A(n2640), .B(n2615), .C(n2608), .D(n2602), .Y(n2423) );
  ivd1_hd U976 ( .A(z_m[21]), .Y(n2671) );
  ivd1_hd U977 ( .A(z_m[20]), .Y(n2527) );
  ivd1_hd U978 ( .A(z_m[18]), .Y(n2533) );
  nd4d1_hd U979 ( .A(n2671), .B(n2539), .C(n2527), .D(n2533), .Y(n2422) );
  ivd1_hd U980 ( .A(z_m[13]), .Y(n2561) );
  ivd1_hd U981 ( .A(z_m[17]), .Y(n2540) );
  nd4d1_hd U982 ( .A(n2578), .B(n2561), .C(n2567), .D(n2540), .Y(n2421) );
  nr4d1_hd U983 ( .A(n2424), .B(n2423), .C(n2422), .D(n2421), .Y(n2425) );
  ivd1_hd U984 ( .A(z_e[9]), .Y(n2691) );
  nr4d1_hd U985 ( .A(z_e[6]), .B(z_e[4]), .C(z_e[3]), .D(z_e[5]), .Y(n2427) );
  nr4d1_hd U986 ( .A(z_m[23]), .B(z_e[0]), .C(n2691), .D(n2502), .Y(n2428) );
  oa211d1_hd U987 ( .A(n2429), .B(n2435), .C(n2488), .D(z_s), .Y(n2430) );
  oa211d1_hd U988 ( .A(n2433), .B(n2432), .C(n2431), .D(n2430), .Y(n361) );
  nr2d1_hd U989 ( .A(z_e[1]), .B(z_e[0]), .Y(n2477) );
  nr2d1_hd U990 ( .A(z_e[3]), .B(n2471), .Y(n2463) );
  ivd1_hd U991 ( .A(z_e[4]), .Y(n2459) );
  nr2d1_hd U992 ( .A(z_e[5]), .B(n2458), .Y(n2449) );
  ivd1_hd U993 ( .A(z_e[6]), .Y(n2445) );
  nr2d1_hd U994 ( .A(z_e[7]), .B(n2444), .Y(n2436) );
  ao211d1_hd U995 ( .A(z_e[7]), .B(n2444), .C(n2487), .D(n2436), .Y(n2440) );
  nd3d1_hd U996 ( .A(n2798), .B(n2912), .C(n2484), .Y(n2478) );
  nd2bd1_hd U997 ( .AN(b_e[2]), .B(n2847), .Y(n2470) );
  nr2d1_hd U998 ( .A(n2478), .B(n2470), .Y(n2469) );
  nd3d1_hd U999 ( .A(n2469), .B(n2832), .C(n2898), .Y(n2464) );
  nd2bd1_hd U1000 ( .AN(b_e[4]), .B(n2802), .Y(n2457) );
  nr2d1_hd U1001 ( .A(n2464), .B(n2457), .Y(n2456) );
  nd3d1_hd U1002 ( .A(n2456), .B(n2823), .C(n2886), .Y(n2451) );
  nr2d1_hd U1003 ( .A(n2451), .B(n2443), .Y(n2442) );
  nr2d1_hd U1004 ( .A(n2442), .B(n2438), .Y(n2437) );
  ao211d1_hd U1005 ( .A(n2442), .B(n2438), .C(n2479), .D(n2437), .Y(n2439) );
  ao211d1_hd U1006 ( .A(n2276), .B(z[30]), .C(n2440), .D(n2439), .Y(n2441) );
  ao21d1_hd U1007 ( .A(n2451), .B(n2443), .C(n2442), .Y(n2448) );
  ivd1_hd U1008 ( .A(n2487), .Y(n2474) );
  oa21d1_hd U1009 ( .A(n2449), .B(n2445), .C(n2444), .Y(n2446) );
  ao22d1_hd U1010 ( .A(n2276), .B(z[29]), .C(n2474), .D(n2446), .Y(n2447) );
  oa211d1_hd U1011 ( .A(n2448), .B(n2479), .C(n2486), .D(n2447), .Y(n363) );
  ao21d1_hd U1012 ( .A(z_e[5]), .B(n2458), .C(n2449), .Y(n2455) );
  nr3d1_hd U1013 ( .A(n2490), .B(n2450), .C(n2925), .Y(n2500) );
  ao22d1_hd U1014 ( .A(a_e[5]), .B(n2495), .C(b_e[5]), .D(n2271), .Y(n2452) );
  oa22d1_hd U1015 ( .A(n2456), .B(n2452), .C(n2479), .D(n2451), .Y(n2453) );
  ao21d1_hd U1016 ( .A(n2276), .B(z[28]), .C(n2453), .Y(n2454) );
  oa211d1_hd U1017 ( .A(n2455), .B(n2487), .C(n2486), .D(n2454), .Y(n364) );
  ao21d1_hd U1018 ( .A(n2464), .B(n2457), .C(n2456), .Y(n2462) );
  oa21d1_hd U1019 ( .A(n2463), .B(n2459), .C(n2458), .Y(n2460) );
  ao22d1_hd U1020 ( .A(n2276), .B(z[27]), .C(n2474), .D(n2460), .Y(n2461) );
  oa211d1_hd U1021 ( .A(n2462), .B(n2479), .C(n2486), .D(n2461), .Y(n365) );
  ao21d1_hd U1022 ( .A(z_e[3]), .B(n2471), .C(n2463), .Y(n2468) );
  ao22d1_hd U1023 ( .A(a_e[3]), .B(n2495), .C(b_e[3]), .D(n2271), .Y(n2465) );
  oa22d1_hd U1024 ( .A(n2469), .B(n2465), .C(n2479), .D(n2464), .Y(n2466) );
  ao21d1_hd U1025 ( .A(n2276), .B(z[26]), .C(n2466), .Y(n2467) );
  oa211d1_hd U1026 ( .A(n2468), .B(n2487), .C(n2486), .D(n2467), .Y(n366) );
  ao21d1_hd U1027 ( .A(n2478), .B(n2470), .C(n2469), .Y(n2476) );
  oa21d1_hd U1028 ( .A(n2477), .B(n2472), .C(n2471), .Y(n2473) );
  ao22d1_hd U1029 ( .A(n2276), .B(z[25]), .C(n2474), .D(n2473), .Y(n2475) );
  oa211d1_hd U1030 ( .A(n2476), .B(n2479), .C(n2486), .D(n2475), .Y(n367) );
  ao21d1_hd U1031 ( .A(z_e[0]), .B(z_e[1]), .C(n2477), .Y(n2483) );
  ao22d1_hd U1032 ( .A(a_e[1]), .B(n2495), .C(b_e[1]), .D(n2271), .Y(n2480) );
  oa22d1_hd U1033 ( .A(n2480), .B(n2484), .C(n2479), .D(n2478), .Y(n2481) );
  ao21d1_hd U1034 ( .A(n2276), .B(z[24]), .C(n2481), .Y(n2482) );
  oa211d1_hd U1035 ( .A(n2483), .B(n2487), .C(n2486), .D(n2482), .Y(n368) );
  ao22d1_hd U1036 ( .A(n2276), .B(z[23]), .C(n2495), .D(n2484), .Y(n2485) );
  oa211d1_hd U1037 ( .A(z_e[0]), .B(n2487), .C(n2486), .D(n2485), .Y(n369) );
  ao22d1_hd U1038 ( .A(b_m[25]), .B(n2271), .C(z_m[22]), .D(n2499), .Y(n2497)
         );
  nd3d1_hd U1039 ( .A(n2491), .B(n2490), .C(n1891), .Y(n2493) );
  ao22d1_hd U1040 ( .A(n2276), .B(z[22]), .C(n2495), .D(n2494), .Y(n2496) );
  scg15d1_hd U1041 ( .A(a_m[25]), .B(n2270), .C(n2497), .D(n2496), .Y(n370) );
  scg4d1_hd U1042 ( .A(b_m[24]), .B(n2271), .C(z_m[21]), .D(n2499), .E(a_m[24]), .F(n2270), .G(n2276), .H(z[21]), .Y(n371) );
  scg4d1_hd U1043 ( .A(b_m[23]), .B(n2271), .C(z_m[20]), .D(n2499), .E(a_m[23]), .F(n2498), .G(n2276), .H(z[20]), .Y(n372) );
  scg4d1_hd U1044 ( .A(b_m[22]), .B(n2271), .C(z_m[19]), .D(n2499), .E(a_m[22]), .F(n2270), .G(n2276), .H(z[19]), .Y(n373) );
  scg4d1_hd U1045 ( .A(b_m[21]), .B(n2271), .C(z_m[18]), .D(n2499), .E(a_m[21]), .F(n2270), .G(n2276), .H(z[18]), .Y(n374) );
  scg4d1_hd U1046 ( .A(b_m[20]), .B(n2271), .C(z_m[17]), .D(n2499), .E(a_m[20]), .F(n2270), .G(n2276), .H(z[17]), .Y(n375) );
  scg4d1_hd U1047 ( .A(b_m[19]), .B(n2271), .C(z_m[16]), .D(n2499), .E(a_m[19]), .F(n2270), .G(n2276), .H(z[16]), .Y(n376) );
  scg4d1_hd U1048 ( .A(b_m[18]), .B(n2271), .C(z_m[15]), .D(n2499), .E(a_m[18]), .F(n2270), .G(n2276), .H(z[15]), .Y(n377) );
  scg4d1_hd U1049 ( .A(a_m[17]), .B(n2270), .C(z_m[14]), .D(n2499), .E(n2271), 
        .F(b_m[17]), .G(n2276), .H(z[14]), .Y(n378) );
  scg4d1_hd U1050 ( .A(b_m[16]), .B(n2271), .C(z_m[13]), .D(n2499), .E(a_m[16]), .F(n2270), .G(n2276), .H(z[13]), .Y(n379) );
  scg4d1_hd U1051 ( .A(b_m[15]), .B(n2271), .C(z_m[12]), .D(n2499), .E(a_m[15]), .F(n2498), .G(n2276), .H(z[12]), .Y(n380) );
  scg4d1_hd U1052 ( .A(b_m[14]), .B(n2271), .C(z_m[11]), .D(n2499), .E(a_m[14]), .F(n2498), .G(n2276), .H(z[11]), .Y(n381) );
  scg4d1_hd U1053 ( .A(b_m[13]), .B(n2271), .C(z_m[10]), .D(n2499), .E(a_m[13]), .F(n2498), .G(n2276), .H(z[10]), .Y(n382) );
  scg4d1_hd U1054 ( .A(b_m[12]), .B(n2271), .C(z_m[9]), .D(n2499), .E(a_m[12]), 
        .F(n2498), .G(n2276), .H(z[9]), .Y(n383) );
  scg4d1_hd U1055 ( .A(b_m[11]), .B(n2271), .C(z_m[8]), .D(n2499), .E(a_m[11]), 
        .F(n2270), .G(n2276), .H(z[8]), .Y(n384) );
  scg4d1_hd U1056 ( .A(b_m[10]), .B(n2271), .C(z_m[7]), .D(n2499), .E(a_m[10]), 
        .F(n2270), .G(n2276), .H(z[7]), .Y(n385) );
  scg4d1_hd U1057 ( .A(b_m[9]), .B(n2271), .C(z_m[6]), .D(n2499), .E(a_m[9]), 
        .F(n2270), .G(n2276), .H(z[6]), .Y(n386) );
  scg4d1_hd U1058 ( .A(b_m[8]), .B(n2271), .C(z_m[5]), .D(n2499), .E(a_m[8]), 
        .F(n2270), .G(n2276), .H(z[5]), .Y(n387) );
  scg4d1_hd U1059 ( .A(b_m[7]), .B(n2271), .C(z_m[4]), .D(n2499), .E(a_m[7]), 
        .F(n2270), .G(n2276), .H(z[4]), .Y(n388) );
  scg4d1_hd U1060 ( .A(b_m[6]), .B(n2271), .C(z_m[3]), .D(n2499), .E(a_m[6]), 
        .F(n2270), .G(n2276), .H(z[3]), .Y(n389) );
  scg4d1_hd U1061 ( .A(b_m[5]), .B(n2271), .C(z_m[2]), .D(n2499), .E(a_m[5]), 
        .F(n2270), .G(n2276), .H(z[2]), .Y(n390) );
  scg4d1_hd U1062 ( .A(b_m[4]), .B(n2271), .C(z_m[1]), .D(n2499), .E(a_m[4]), 
        .F(n2270), .G(n2276), .H(z[1]), .Y(n391) );
  scg4d1_hd U1063 ( .A(b_m[3]), .B(n2271), .C(z_m[0]), .D(n2499), .E(a_m[3]), 
        .F(n2498), .G(n2276), .H(z[0]), .Y(n392) );
  ao22d1_hd U1064 ( .A(n2676), .B(sum[0]), .C(sticky), .D(n2508), .Y(n2505) );
  scg16d1_hd U1065 ( .A(n2502), .B(n2501), .C(z_e[9]), .Y(n2506) );
  nr2d1_hd U1066 ( .A(n2503), .B(n2506), .Y(n2930) );
  ao22d1_hd U1067 ( .A(n2507), .B(round_bit), .C(n2648), .D(sum[1]), .Y(n2504)
         );
  scg21d1_hd U1068 ( .A(n2506), .B(z_e[0]), .C(z_m[23]), .D(n2930), .Y(n2935)
         );
  ao21d1_hd U1069 ( .A(n2935), .B(n1291), .C(n2507), .Y(n2675) );
  ao22d1_hd U1070 ( .A(n2648), .B(sum[2]), .C(n2272), .D(sum[1]), .Y(n2510) );
  nd3d1_hd U1071 ( .A(n2511), .B(guard), .C(n1222), .Y(n2509) );
  oa211d1_hd U1072 ( .A(n2512), .B(n1222), .C(n2510), .D(n2509), .Y(n394) );
  oa211d1_hd U1073 ( .A(sticky), .B(n2513), .C(guard), .D(n2677), .Y(n2514) );
  ao22d1_hd U1074 ( .A(n2648), .B(sum[26]), .C(n2272), .D(sum[25]), .Y(n2518)
         );
  ivd1_hd U1075 ( .A(n2669), .Y(n2515) );
  nd3d1_hd U1076 ( .A(z_m[0]), .B(z_m[1]), .C(z_m[2]), .Y(n2621) );
  nr3d1_hd U1077 ( .A(n2621), .B(n2626), .C(n2640), .Y(n2609) );
  nd3d1_hd U1078 ( .A(n2609), .B(z_m[5]), .C(z_m[6]), .Y(n2597) );
  nr3d1_hd U1079 ( .A(n2597), .B(n2602), .C(n2614), .Y(n2585) );
  nd3d1_hd U1080 ( .A(n2585), .B(z_m[9]), .C(z_m[10]), .Y(n2573) );
  nr3d1_hd U1081 ( .A(n2573), .B(n2590), .C(n2578), .Y(n2562) );
  nd3d1_hd U1082 ( .A(n2562), .B(z_m[13]), .C(z_m[14]), .Y(n2547) );
  nr2d1_hd U1083 ( .A(n2548), .B(n2547), .Y(n2534) );
  nd3d1_hd U1084 ( .A(n2534), .B(z_m[17]), .C(z_m[18]), .Y(n2668) );
  nr2d1_hd U1085 ( .A(n2668), .B(n2634), .Y(n2530) );
  oa21d1_hd U1086 ( .A(z_m[22]), .B(n2663), .C(n2661), .Y(n2516) );
  ao21d1_hd U1087 ( .A(n2668), .B(n2677), .C(n2635), .Y(n2528) );
  oa21d1_hd U1088 ( .A(z_m[21]), .B(n2634), .C(n2519), .Y(n2658) );
  ao22d1_hd U1089 ( .A(z_m[21]), .B(n2516), .C(z_m[22]), .D(n2658), .Y(n2517)
         );
  oa211d1_hd U1090 ( .A(n2670), .B(n2649), .C(n2518), .D(n2517), .Y(n395) );
  ao22d1_hd U1091 ( .A(n2648), .B(sum[25]), .C(n2272), .D(sum[24]), .Y(n2522)
         );
  ao22d1_hd U1092 ( .A(z_m[21]), .B(n2519), .C(n2663), .D(n2671), .Y(n2520) );
  ao21d1_hd U1093 ( .A(n2653), .B(z_m[20]), .C(n2520), .Y(n2521) );
  oa211d1_hd U1094 ( .A(n2659), .B(n2649), .C(n2522), .D(n2521), .Y(n396) );
  ao21d1_hd U1095 ( .A(n2530), .B(n2527), .C(n2653), .Y(n2526) );
  ao22d1_hd U1096 ( .A(n2648), .B(sum[24]), .C(n2272), .D(sum[23]), .Y(n2525)
         );
  oa21d1_hd U1097 ( .A(z_m[19]), .B(n2634), .C(n2528), .Y(n2523) );
  ao22d1_hd U1098 ( .A(z_m[21]), .B(n2642), .C(z_m[20]), .D(n2523), .Y(n2524)
         );
  oa211d1_hd U1099 ( .A(n2526), .B(n2539), .C(n2525), .D(n2524), .Y(n397) );
  ao22d1_hd U1100 ( .A(n2648), .B(sum[23]), .C(n2272), .D(sum[22]), .Y(n2532)
         );
  oa22d1_hd U1101 ( .A(n2528), .B(n2539), .C(n2527), .D(n2649), .Y(n2529) );
  ao21d1_hd U1102 ( .A(n2530), .B(n2539), .C(n2529), .Y(n2531) );
  oa211d1_hd U1103 ( .A(n2661), .B(n2533), .C(n2532), .D(n2531), .Y(n398) );
  ao22d1_hd U1104 ( .A(n2648), .B(sum[22]), .C(n2272), .D(sum[21]), .Y(n2538)
         );
  oa21d1_hd U1105 ( .A(z_m[18]), .B(n2541), .C(n2661), .Y(n2536) );
  scg20d1_hd U1106 ( .A(n2958), .B(n2534), .C(n2635), .Y(n2542) );
  oa21d1_hd U1107 ( .A(z_m[17]), .B(n2634), .C(n2542), .Y(n2535) );
  ao22d1_hd U1108 ( .A(z_m[17]), .B(n2536), .C(z_m[18]), .D(n2535), .Y(n2537)
         );
  oa211d1_hd U1109 ( .A(n2539), .B(n2649), .C(n2538), .D(n2537), .Y(n399) );
  ao22d1_hd U1110 ( .A(n2648), .B(sum[21]), .C(n2272), .D(sum[20]), .Y(n2545)
         );
  ao22d1_hd U1111 ( .A(z_m[17]), .B(n2542), .C(n2541), .D(n2540), .Y(n2543) );
  ao21d1_hd U1112 ( .A(z_m[18]), .B(n2642), .C(n2543), .Y(n2544) );
  oa211d1_hd U1113 ( .A(n2661), .B(n2546), .C(n2545), .D(n2544), .Y(n400) );
  ao22d1_hd U1114 ( .A(n2648), .B(sum[20]), .C(n2272), .D(sum[19]), .Y(n2553)
         );
  ivd1_hd U1115 ( .A(n2547), .Y(n2556) );
  oa21d1_hd U1116 ( .A(n2556), .B(n2958), .C(n2656), .Y(n2554) );
  ao22d1_hd U1117 ( .A(z_m[16]), .B(n2554), .C(z_m[17]), .D(n2642), .Y(n2552)
         );
  nr2d1_hd U1118 ( .A(n2555), .B(n2547), .Y(n2549) );
  oa211d1_hd U1119 ( .A(z_m[16]), .B(n2549), .C(n2660), .D(n2548), .Y(n2551)
         );
  nd4d1_hd U1120 ( .A(n2553), .B(n2552), .C(n2551), .D(n2550), .Y(n401) );
  ao22d1_hd U1121 ( .A(n2648), .B(sum[19]), .C(n2272), .D(sum[18]), .Y(n2560)
         );
  ao22d1_hd U1122 ( .A(z_m[15]), .B(n2554), .C(z_m[16]), .D(n2642), .Y(n2559)
         );
  nd3d1_hd U1123 ( .A(n2556), .B(n2660), .C(n2555), .Y(n2558) );
  nd4d1_hd U1124 ( .A(n2560), .B(n2559), .C(n2558), .D(n2557), .Y(n402) );
  oa21d1_hd U1125 ( .A(n2562), .B(n2958), .C(n2656), .Y(n2570) );
  ao21d1_hd U1126 ( .A(n2660), .B(n2561), .C(n2570), .Y(n2566) );
  ao22d1_hd U1127 ( .A(n2648), .B(sum[18]), .C(n2272), .D(sum[17]), .Y(n2565)
         );
  oa21d1_hd U1128 ( .A(z_m[14]), .B(n2568), .C(n2661), .Y(n2563) );
  ao22d1_hd U1129 ( .A(z_m[15]), .B(n2642), .C(z_m[13]), .D(n2563), .Y(n2564)
         );
  oa211d1_hd U1130 ( .A(n2566), .B(n2567), .C(n2565), .D(n2564), .Y(n403) );
  ao22d1_hd U1131 ( .A(n2648), .B(sum[17]), .C(n2272), .D(sum[16]), .Y(n2572)
         );
  oa22d1_hd U1132 ( .A(z_m[13]), .B(n2568), .C(n2649), .D(n2567), .Y(n2569) );
  ao21d1_hd U1133 ( .A(z_m[13]), .B(n2570), .C(n2569), .Y(n2571) );
  oa211d1_hd U1134 ( .A(n2661), .B(n2578), .C(n2572), .D(n2571), .Y(n404) );
  nr2d1_hd U1135 ( .A(n2573), .B(n2634), .Y(n2581) );
  ao21d1_hd U1136 ( .A(n2581), .B(n2578), .C(n2653), .Y(n2577) );
  ao22d1_hd U1137 ( .A(n2648), .B(sum[16]), .C(n2272), .D(sum[15]), .Y(n2576)
         );
  ao21d1_hd U1138 ( .A(n2677), .B(n2573), .C(n2635), .Y(n2579) );
  oa21d1_hd U1139 ( .A(z_m[11]), .B(n2634), .C(n2579), .Y(n2574) );
  ao22d1_hd U1140 ( .A(z_m[12]), .B(n2574), .C(z_m[13]), .D(n2642), .Y(n2575)
         );
  oa211d1_hd U1141 ( .A(n2577), .B(n2590), .C(n2576), .D(n2575), .Y(n405) );
  ao22d1_hd U1142 ( .A(n2648), .B(sum[15]), .C(n2272), .D(sum[14]), .Y(n2583)
         );
  oa22d1_hd U1143 ( .A(n2579), .B(n2590), .C(n2578), .D(n2649), .Y(n2580) );
  ao21d1_hd U1144 ( .A(n2581), .B(n2590), .C(n2580), .Y(n2582) );
  oa211d1_hd U1145 ( .A(n2661), .B(n2584), .C(n2583), .D(n2582), .Y(n406) );
  ao22d1_hd U1146 ( .A(n2648), .B(sum[14]), .C(n2272), .D(sum[13]), .Y(n2589)
         );
  oa21d1_hd U1147 ( .A(z_m[10]), .B(n2592), .C(n2661), .Y(n2587) );
  scg20d1_hd U1148 ( .A(n2958), .B(n2585), .C(n2635), .Y(n2593) );
  oa21d1_hd U1149 ( .A(z_m[9]), .B(n2634), .C(n2593), .Y(n2586) );
  ao22d1_hd U1150 ( .A(z_m[9]), .B(n2587), .C(z_m[10]), .D(n2586), .Y(n2588)
         );
  oa211d1_hd U1151 ( .A(n2590), .B(n2649), .C(n2589), .D(n2588), .Y(n407) );
  ao22d1_hd U1152 ( .A(n2648), .B(sum[13]), .C(n2272), .D(sum[12]), .Y(n2596)
         );
  ao22d1_hd U1153 ( .A(z_m[9]), .B(n2593), .C(n2592), .D(n2591), .Y(n2594) );
  ao21d1_hd U1154 ( .A(z_m[10]), .B(n2642), .C(n2594), .Y(n2595) );
  oa211d1_hd U1155 ( .A(n2661), .B(n2602), .C(n2596), .D(n2595), .Y(n408) );
  nr2d1_hd U1156 ( .A(n2597), .B(n2634), .Y(n2605) );
  ao21d1_hd U1157 ( .A(n2605), .B(n2602), .C(n2653), .Y(n2601) );
  ao22d1_hd U1158 ( .A(n2648), .B(sum[12]), .C(n2272), .D(sum[11]), .Y(n2600)
         );
  ao21d1_hd U1159 ( .A(n2677), .B(n2597), .C(n2635), .Y(n2603) );
  oa21d1_hd U1160 ( .A(z_m[7]), .B(n2634), .C(n2603), .Y(n2598) );
  ao22d1_hd U1161 ( .A(z_m[8]), .B(n2598), .C(z_m[9]), .D(n2642), .Y(n2599) );
  oa211d1_hd U1162 ( .A(n2601), .B(n2614), .C(n2600), .D(n2599), .Y(n409) );
  ao22d1_hd U1163 ( .A(n2648), .B(sum[11]), .C(n2272), .D(sum[10]), .Y(n2607)
         );
  oa22d1_hd U1164 ( .A(n2603), .B(n2614), .C(n2602), .D(n2649), .Y(n2604) );
  ao21d1_hd U1165 ( .A(n2605), .B(n2614), .C(n2604), .Y(n2606) );
  oa211d1_hd U1166 ( .A(n2661), .B(n2608), .C(n2607), .D(n2606), .Y(n410) );
  ao22d1_hd U1167 ( .A(n2648), .B(sum[10]), .C(n2272), .D(sum[9]), .Y(n2613)
         );
  oa21d1_hd U1168 ( .A(z_m[6]), .B(n2616), .C(n2661), .Y(n2611) );
  scg20d1_hd U1169 ( .A(n2958), .B(n2609), .C(n2635), .Y(n2617) );
  oa21d1_hd U1170 ( .A(z_m[5]), .B(n2634), .C(n2617), .Y(n2610) );
  ao22d1_hd U1171 ( .A(z_m[5]), .B(n2611), .C(z_m[6]), .D(n2610), .Y(n2612) );
  oa211d1_hd U1172 ( .A(n2614), .B(n2649), .C(n2613), .D(n2612), .Y(n411) );
  ao22d1_hd U1173 ( .A(n2648), .B(sum[9]), .C(n2272), .D(sum[8]), .Y(n2620) );
  ao22d1_hd U1174 ( .A(z_m[5]), .B(n2617), .C(n2616), .D(n2615), .Y(n2618) );
  ao21d1_hd U1175 ( .A(z_m[6]), .B(n2642), .C(n2618), .Y(n2619) );
  oa211d1_hd U1176 ( .A(n2661), .B(n2626), .C(n2620), .D(n2619), .Y(n412) );
  nr2d1_hd U1177 ( .A(n2621), .B(n2634), .Y(n2629) );
  ao21d1_hd U1178 ( .A(n2629), .B(n2626), .C(n2653), .Y(n2625) );
  ao22d1_hd U1179 ( .A(n2648), .B(sum[8]), .C(n2272), .D(sum[7]), .Y(n2624) );
  ao21d1_hd U1180 ( .A(n2677), .B(n2621), .C(n2635), .Y(n2627) );
  oa21d1_hd U1181 ( .A(z_m[3]), .B(n2634), .C(n2627), .Y(n2622) );
  ao22d1_hd U1182 ( .A(z_m[4]), .B(n2622), .C(z_m[5]), .D(n2642), .Y(n2623) );
  oa211d1_hd U1183 ( .A(n2625), .B(n2640), .C(n2624), .D(n2623), .Y(n413) );
  ao22d1_hd U1184 ( .A(n2648), .B(sum[7]), .C(n2272), .D(sum[6]), .Y(n2631) );
  oa22d1_hd U1185 ( .A(n2627), .B(n2640), .C(n2626), .D(n2649), .Y(n2628) );
  ao21d1_hd U1186 ( .A(n2629), .B(n2640), .C(n2628), .Y(n2630) );
  oa211d1_hd U1187 ( .A(n2661), .B(n2632), .C(n2631), .D(n2630), .Y(n414) );
  ao22d1_hd U1188 ( .A(n2648), .B(sum[6]), .C(n2272), .D(sum[5]), .Y(n2639) );
  oa21d1_hd U1189 ( .A(z_m[2]), .B(n2633), .C(n2661), .Y(n2637) );
  nr2d1_hd U1190 ( .A(z_m[0]), .B(n2634), .Y(n2652) );
  nr2d1_hd U1191 ( .A(n2635), .B(n2652), .Y(n2646) );
  ao22d1_hd U1192 ( .A(z_m[1]), .B(n2637), .C(z_m[2]), .D(n2636), .Y(n2638) );
  oa211d1_hd U1193 ( .A(n2640), .B(n2649), .C(n2639), .D(n2638), .Y(n415) );
  ao22d1_hd U1194 ( .A(n2648), .B(sum[5]), .C(n2272), .D(sum[4]), .Y(n2645) );
  ao22d1_hd U1195 ( .A(z_m[0]), .B(n2643), .C(z_m[2]), .D(n2642), .Y(n2644) );
  oa211d1_hd U1196 ( .A(n2646), .B(n2650), .C(n2645), .D(n2644), .Y(n416) );
  ao22d1_hd U1197 ( .A(n2648), .B(sum[4]), .C(n2272), .D(sum[3]), .Y(n2655) );
  nr2d1_hd U1198 ( .A(n2650), .B(n2649), .Y(n2651) );
  ao211d1_hd U1199 ( .A(n2653), .B(guard), .C(n2652), .D(n2651), .Y(n2654) );
  oa211d1_hd U1200 ( .A(n2657), .B(n2656), .C(n2655), .D(n2654), .Y(n417) );
  ao21d1_hd U1201 ( .A(n2660), .B(n2659), .C(n2658), .Y(n2666) );
  oa21d1_hd U1202 ( .A(n2663), .B(n2662), .C(n2661), .Y(n2664) );
  ao22d1_hd U1203 ( .A(n2676), .B(sum[26]), .C(z_m[22]), .D(n2664), .Y(n2665)
         );
  oa211d1_hd U1204 ( .A(n2666), .B(n2670), .C(n2665), .D(n2674), .Y(n418) );
  nr4d1_hd U1205 ( .A(n2671), .B(n2670), .C(n2669), .D(n2668), .Y(n2672) );
  nd4d1_hd U1206 ( .A(n2677), .B(guard), .C(z_m[22]), .D(n2672), .Y(n2673) );
  nd4d1_hd U1207 ( .A(n2675), .B(n1284), .C(n2674), .D(n2673), .Y(n2688) );
  nr3d1_hd U1208 ( .A(n2677), .B(state[1]), .C(n2676), .Y(n2678) );
  ao22d1_hd U1209 ( .A(a_e[8]), .B(n2268), .C(n2693), .D(C91_DATA2_8), .Y(
        n2679) );
  scg14d1_hd U1210 ( .A(z_e[8]), .B(n2690), .C(n2679), .Y(n419) );
  ao22d1_hd U1211 ( .A(z_e[7]), .B(n2690), .C(n2693), .D(C91_DATA2_7), .Y(
        n2680) );
  oa21d1_hd U1212 ( .A(n2807), .B(n1284), .C(n2680), .Y(n420) );
  ao22d1_hd U1213 ( .A(z_e[6]), .B(n2690), .C(n2693), .D(C91_DATA2_6), .Y(
        n2681) );
  oa21d1_hd U1214 ( .A(n2803), .B(n1284), .C(n2681), .Y(n421) );
  ao22d1_hd U1215 ( .A(z_e[5]), .B(n2690), .C(n2693), .D(C91_DATA2_5), .Y(
        n2682) );
  oa21d1_hd U1216 ( .A(n2823), .B(n1284), .C(n2682), .Y(n422) );
  ao22d1_hd U1217 ( .A(z_e[4]), .B(n2690), .C(n2693), .D(C91_DATA2_4), .Y(
        n2683) );
  oa21d1_hd U1218 ( .A(n2802), .B(n1284), .C(n2683), .Y(n423) );
  ao22d1_hd U1219 ( .A(z_e[3]), .B(n2690), .C(n2693), .D(C91_DATA2_3), .Y(
        n2684) );
  oa21d1_hd U1220 ( .A(n2832), .B(n1284), .C(n2684), .Y(n424) );
  ao22d1_hd U1221 ( .A(z_e[2]), .B(n2690), .C(n2693), .D(C91_DATA2_2), .Y(
        n2685) );
  oa21d1_hd U1222 ( .A(n2847), .B(n1284), .C(n2685), .Y(n425) );
  ao22d1_hd U1223 ( .A(z_e[1]), .B(n2690), .C(n2693), .D(C91_DATA2_1), .Y(
        n2686) );
  oa21d1_hd U1224 ( .A(n2798), .B(n1284), .C(n2686), .Y(n426) );
  ao22d1_hd U1225 ( .A(a_e[0]), .B(n2268), .C(n2693), .D(n2689), .Y(n2687) );
  oa21d1_hd U1226 ( .A(n2689), .B(n2688), .C(n2687), .Y(n427) );
  ao22d1_hd U1227 ( .A(a_e[9]), .B(n2268), .C(z_e[9]), .D(n2690), .Y(n2696) );
  ao22d1_hd U1228 ( .A(n1291), .B(z_e[9]), .C(n2691), .D(n2934), .Y(n2694) );
  oa211d1_hd U1229 ( .A(DP_OP_154J4_137_6175_n2), .B(n2694), .C(n2693), .D(
        n2692), .Y(n2695) );
  ao22d1_hd U1230 ( .A(b_m[25]), .B(n2949), .C(n2277), .D(b[21]), .Y(n2697) );
  oa21d1_hd U1231 ( .A(n2698), .B(n2275), .C(n2697), .Y(n429) );
  ao22d1_hd U1232 ( .A(b_m[24]), .B(n2949), .C(n2278), .D(b[20]), .Y(n2699) );
  oa21d1_hd U1233 ( .A(n2700), .B(n2275), .C(n2699), .Y(n430) );
  ao22d1_hd U1234 ( .A(b_m[23]), .B(n2949), .C(n2279), .D(b[19]), .Y(n2701) );
  oa21d1_hd U1235 ( .A(n2702), .B(n2275), .C(n2701), .Y(n431) );
  ao22d1_hd U1236 ( .A(b_m[22]), .B(n2949), .C(n2278), .D(b[18]), .Y(n2703) );
  oa21d1_hd U1237 ( .A(n2704), .B(n2275), .C(n2703), .Y(n432) );
  ao22d1_hd U1238 ( .A(b_m[21]), .B(n2949), .C(n2279), .D(b[17]), .Y(n2705) );
  oa21d1_hd U1239 ( .A(n2706), .B(n2275), .C(n2705), .Y(n433) );
  ao22d1_hd U1240 ( .A(b_m[20]), .B(n2949), .C(n2278), .D(b[16]), .Y(n2707) );
  oa21d1_hd U1241 ( .A(n2708), .B(n2275), .C(n2707), .Y(n434) );
  ao22d1_hd U1242 ( .A(b_m[19]), .B(n2949), .C(n2279), .D(b[15]), .Y(n2709) );
  oa21d1_hd U1243 ( .A(n2710), .B(n2275), .C(n2709), .Y(n435) );
  ao22d1_hd U1244 ( .A(b_m[18]), .B(n2949), .C(n2279), .D(b[14]), .Y(n2711) );
  oa21d1_hd U1245 ( .A(n2712), .B(n2275), .C(n2711), .Y(n436) );
  ao22d1_hd U1246 ( .A(b_m[17]), .B(n2949), .C(n2278), .D(b[13]), .Y(n2713) );
  oa21d1_hd U1247 ( .A(n2714), .B(n2275), .C(n2713), .Y(n437) );
  ao22d1_hd U1248 ( .A(b_m[16]), .B(n2949), .C(n2279), .D(b[12]), .Y(n2715) );
  oa21d1_hd U1249 ( .A(n2716), .B(n2275), .C(n2715), .Y(n438) );
  ao22d1_hd U1250 ( .A(b_m[15]), .B(n2949), .C(n2278), .D(b[11]), .Y(n2717) );
  oa21d1_hd U1251 ( .A(n2718), .B(n2275), .C(n2717), .Y(n439) );
  ao22d1_hd U1252 ( .A(b_m[14]), .B(n2949), .C(n2279), .D(b[10]), .Y(n2719) );
  oa21d1_hd U1253 ( .A(n2720), .B(n2275), .C(n2719), .Y(n440) );
  ao22d1_hd U1254 ( .A(b_m[13]), .B(n2949), .C(n2278), .D(b[9]), .Y(n2721) );
  oa21d1_hd U1255 ( .A(n2722), .B(n2275), .C(n2721), .Y(n441) );
  ao22d1_hd U1256 ( .A(b_m[12]), .B(n2949), .C(n2278), .D(b[8]), .Y(n2723) );
  oa21d1_hd U1257 ( .A(n2724), .B(n2275), .C(n2723), .Y(n442) );
  ao22d1_hd U1258 ( .A(b_m[11]), .B(n2949), .C(n2278), .D(b[7]), .Y(n2725) );
  oa21d1_hd U1259 ( .A(n2726), .B(n2275), .C(n2725), .Y(n443) );
  ao22d1_hd U1260 ( .A(b_m[10]), .B(n2949), .C(n2278), .D(b[6]), .Y(n2727) );
  oa21d1_hd U1261 ( .A(n2728), .B(n2275), .C(n2727), .Y(n444) );
  ao22d1_hd U1262 ( .A(b_m[9]), .B(n2949), .C(n2278), .D(b[5]), .Y(n2729) );
  oa21d1_hd U1263 ( .A(n2730), .B(n2275), .C(n2729), .Y(n445) );
  ao22d1_hd U1264 ( .A(b_m[8]), .B(n2949), .C(n2278), .D(b[4]), .Y(n2731) );
  oa21d1_hd U1265 ( .A(n2732), .B(n2275), .C(n2731), .Y(n446) );
  ao22d1_hd U1266 ( .A(b_m[7]), .B(n2949), .C(n2278), .D(b[3]), .Y(n2733) );
  oa21d1_hd U1267 ( .A(n2734), .B(n2275), .C(n2733), .Y(n447) );
  ao22d1_hd U1268 ( .A(b_m[6]), .B(n2949), .C(n2278), .D(b[2]), .Y(n2735) );
  oa21d1_hd U1269 ( .A(n2736), .B(n2275), .C(n2735), .Y(n448) );
  ao22d1_hd U1270 ( .A(b_m[5]), .B(n2949), .C(n2278), .D(b[1]), .Y(n2737) );
  oa21d1_hd U1271 ( .A(n2738), .B(n2275), .C(n2737), .Y(n449) );
  ao22d1_hd U1272 ( .A(b_m[4]), .B(n2949), .C(n2278), .D(b[0]), .Y(n2739) );
  oa21d1_hd U1273 ( .A(n2740), .B(n2275), .C(n2739), .Y(n450) );
  oa22d1_hd U1274 ( .A(n2741), .B(n2275), .C(n2740), .D(n2742), .Y(n451) );
  oa22d1_hd U1275 ( .A(n2743), .B(n2275), .C(n2741), .D(n2742), .Y(n452) );
  oa22d1_hd U1276 ( .A(n2279), .B(n2744), .C(n2743), .D(n2742), .Y(n453) );
  ao22d1_hd U1277 ( .A(a_m[25]), .B(n2793), .C(n2278), .D(a[21]), .Y(n2745) );
  oa21d1_hd U1278 ( .A(n2746), .B(n2273), .C(n2745), .Y(n454) );
  ao22d1_hd U1279 ( .A(a_m[24]), .B(n2793), .C(n2278), .D(a[20]), .Y(n2747) );
  oa21d1_hd U1280 ( .A(n2748), .B(n2273), .C(n2747), .Y(n455) );
  ao22d1_hd U1281 ( .A(a_m[23]), .B(n2793), .C(n2278), .D(a[19]), .Y(n2749) );
  oa21d1_hd U1282 ( .A(n2750), .B(n2273), .C(n2749), .Y(n456) );
  ao22d1_hd U1283 ( .A(a_m[22]), .B(n2793), .C(n2278), .D(a[18]), .Y(n2751) );
  oa21d1_hd U1284 ( .A(n2752), .B(n2273), .C(n2751), .Y(n457) );
  ao22d1_hd U1285 ( .A(a_m[21]), .B(n2793), .C(n2278), .D(a[17]), .Y(n2753) );
  oa21d1_hd U1286 ( .A(n2754), .B(n2273), .C(n2753), .Y(n458) );
  ao22d1_hd U1287 ( .A(a_m[20]), .B(n2793), .C(n2278), .D(a[16]), .Y(n2755) );
  oa21d1_hd U1288 ( .A(n2756), .B(n2273), .C(n2755), .Y(n459) );
  ao22d1_hd U1289 ( .A(a_m[19]), .B(n2793), .C(n2278), .D(a[15]), .Y(n2757) );
  oa21d1_hd U1290 ( .A(n2758), .B(n2273), .C(n2757), .Y(n460) );
  ao22d1_hd U1291 ( .A(a_m[18]), .B(n2793), .C(n2278), .D(a[14]), .Y(n2759) );
  oa21d1_hd U1292 ( .A(n2760), .B(n2273), .C(n2759), .Y(n461) );
  ao22d1_hd U1293 ( .A(a_m[17]), .B(n2793), .C(n2278), .D(a[13]), .Y(n2761) );
  oa21d1_hd U1294 ( .A(n2762), .B(n2273), .C(n2761), .Y(n462) );
  ao22d1_hd U1295 ( .A(a_m[16]), .B(n2793), .C(n2278), .D(a[12]), .Y(n2763) );
  oa21d1_hd U1296 ( .A(n2764), .B(n2273), .C(n2763), .Y(n463) );
  ao22d1_hd U1297 ( .A(a_m[15]), .B(n2793), .C(n2278), .D(a[11]), .Y(n2765) );
  oa21d1_hd U1298 ( .A(n2766), .B(n2273), .C(n2765), .Y(n464) );
  ao22d1_hd U1299 ( .A(a_m[14]), .B(n2793), .C(n2277), .D(a[10]), .Y(n2767) );
  oa21d1_hd U1300 ( .A(n2768), .B(n2273), .C(n2767), .Y(n465) );
  ao22d1_hd U1301 ( .A(a_m[13]), .B(n2793), .C(n2277), .D(a[9]), .Y(n2769) );
  oa21d1_hd U1302 ( .A(n2770), .B(n2273), .C(n2769), .Y(n466) );
  ao22d1_hd U1303 ( .A(a_m[12]), .B(n2793), .C(n2277), .D(a[8]), .Y(n2771) );
  oa21d1_hd U1304 ( .A(n2772), .B(n2273), .C(n2771), .Y(n467) );
  ao22d1_hd U1305 ( .A(a_m[11]), .B(n2793), .C(n2277), .D(a[7]), .Y(n2773) );
  oa21d1_hd U1306 ( .A(n2774), .B(n2273), .C(n2773), .Y(n468) );
  ao22d1_hd U1307 ( .A(a_m[10]), .B(n2793), .C(n2277), .D(a[6]), .Y(n2775) );
  oa21d1_hd U1308 ( .A(n2776), .B(n2273), .C(n2775), .Y(n469) );
  ao22d1_hd U1309 ( .A(a_m[9]), .B(n2793), .C(n2277), .D(a[5]), .Y(n2777) );
  oa21d1_hd U1310 ( .A(n2778), .B(n2273), .C(n2777), .Y(n470) );
  ao22d1_hd U1311 ( .A(a_m[8]), .B(n2793), .C(n2277), .D(a[4]), .Y(n2779) );
  oa21d1_hd U1312 ( .A(n2780), .B(n2273), .C(n2779), .Y(n471) );
  ao22d1_hd U1313 ( .A(a_m[7]), .B(n2793), .C(n2277), .D(a[3]), .Y(n2781) );
  oa21d1_hd U1314 ( .A(n2782), .B(n2796), .C(n2781), .Y(n472) );
  ao22d1_hd U1315 ( .A(a_m[6]), .B(n2793), .C(n2278), .D(a[2]), .Y(n2783) );
  oa21d1_hd U1316 ( .A(n2784), .B(n2796), .C(n2783), .Y(n473) );
  ao22d1_hd U1317 ( .A(a_m[5]), .B(n2793), .C(n2277), .D(a[1]), .Y(n2785) );
  oa21d1_hd U1318 ( .A(n2786), .B(n2796), .C(n2785), .Y(n474) );
  ao22d1_hd U1319 ( .A(a_m[4]), .B(n2793), .C(n2277), .D(a[0]), .Y(n2787) );
  oa21d1_hd U1320 ( .A(n2788), .B(n2796), .C(n2787), .Y(n475) );
  oa22d1_hd U1321 ( .A(n2789), .B(n2273), .C(n2788), .D(n2790), .Y(n476) );
  oa22d1_hd U1322 ( .A(n2791), .B(n2273), .C(n2789), .D(n2790), .Y(n477) );
  oa22d1_hd U1323 ( .A(n2279), .B(n2792), .C(n2791), .D(n2790), .Y(n478) );
  ao22d1_hd U1324 ( .A(a_m[26]), .B(n2793), .C(n2277), .D(a[22]), .Y(n2794) );
  oa21d1_hd U1325 ( .A(n2795), .B(n2796), .C(n2794), .Y(n479) );
  nr2d1_hd U1326 ( .A(n2838), .B(n2798), .Y(n2841) );
  ao21d1_hd U1327 ( .A(n2801), .B(n2889), .C(n2855), .Y(n2825) );
  ivd1_hd U1328 ( .A(n2825), .Y(n2834) );
  ao21d1_hd U1329 ( .A(n2889), .B(n2799), .C(n2834), .Y(n2824) );
  oa21d1_hd U1330 ( .A(n2803), .B(n2823), .C(n2889), .Y(n2800) );
  ao21d1_hd U1331 ( .A(n2840), .B(n2807), .C(n2809), .Y(n2858) );
  ivd1_hd U1332 ( .A(a[25]), .Y(n2843) );
  nr2d1_hd U1333 ( .A(n2851), .B(n2843), .Y(n2842) );
  ivd1_hd U1334 ( .A(a[27]), .Y(n2827) );
  nr2d1_hd U1335 ( .A(n2835), .B(n2827), .Y(n2826) );
  ivd1_hd U1336 ( .A(a[29]), .Y(n2813) );
  nr2d1_hd U1337 ( .A(n2820), .B(n2813), .Y(n2806) );
  nr2d1_hd U1338 ( .A(n2806), .B(n2280), .Y(n2816) );
  nr2d1_hd U1339 ( .A(n2859), .B(n2801), .Y(n2833) );
  nr2d1_hd U1340 ( .A(n2802), .B(n2831), .Y(n2819) );
  nr2d1_hd U1341 ( .A(n2803), .B(n2818), .Y(n2808) );
  nd3d1_hd U1342 ( .A(a_e[7]), .B(n2808), .C(n2805), .Y(n2804) );
  oa211d1_hd U1343 ( .A(n2858), .B(n2805), .C(n2860), .D(n2804), .Y(n480) );
  ao22d1_hd U1344 ( .A(a_e[7]), .B(n2809), .C(n2808), .D(n2807), .Y(n2810) );
  oa211d1_hd U1345 ( .A(n2812), .B(n2811), .C(n2810), .D(n2860), .Y(n481) );
  oa21d1_hd U1346 ( .A(a_e[5]), .B(n2859), .C(n2824), .Y(n2814) );
  ao22d1_hd U1347 ( .A(n2816), .B(n2815), .C(a_e[6]), .D(n2814), .Y(n2817) );
  oa211d1_hd U1348 ( .A(a_e[6]), .B(n2818), .C(n2817), .D(n2853), .Y(n482) );
  ao21d1_hd U1349 ( .A(n2819), .B(n2823), .C(n2861), .Y(n2822) );
  oa211d1_hd U1350 ( .A(n2826), .B(a[28]), .C(n2279), .D(n2820), .Y(n2821) );
  oa211d1_hd U1351 ( .A(n2824), .B(n2823), .C(n2822), .D(n2821), .Y(n483) );
  oa21d1_hd U1352 ( .A(a_e[3]), .B(n2859), .C(n2825), .Y(n2829) );
  ao211d1_hd U1353 ( .A(n2835), .B(n2827), .C(n2826), .D(n2280), .Y(n2828) );
  ao211d1_hd U1354 ( .A(a_e[4]), .B(n2829), .C(n2861), .D(n2828), .Y(n2830) );
  oa21d1_hd U1355 ( .A(a_e[4]), .B(n2831), .C(n2830), .Y(n484) );
  ao22d1_hd U1356 ( .A(a_e[3]), .B(n2834), .C(n2833), .D(n2832), .Y(n2837) );
  oa211d1_hd U1357 ( .A(n2842), .B(a[26]), .C(n2279), .D(n2835), .Y(n2836) );
  nd3d1_hd U1358 ( .A(n2837), .B(n2853), .C(n2836), .Y(n485) );
  nr2d1_hd U1359 ( .A(a_e[1]), .B(n2859), .Y(n2850) );
  nr2d1_hd U1360 ( .A(n2850), .B(n2849), .Y(n2848) );
  ao211d1_hd U1361 ( .A(n2851), .B(n2843), .C(n2842), .D(n2280), .Y(n2844) );
  nr2d1_hd U1362 ( .A(n2845), .B(n2844), .Y(n2846) );
  oa211d1_hd U1363 ( .A(n2848), .B(n2847), .C(n2846), .D(n2853), .Y(n486) );
  ao22d1_hd U1364 ( .A(a_e[0]), .B(n2850), .C(a_e[1]), .D(n2849), .Y(n2854) );
  oa211d1_hd U1365 ( .A(a[23]), .B(a[24]), .C(n2279), .D(n2851), .Y(n2852) );
  nd3d1_hd U1366 ( .A(n2854), .B(n2853), .C(n2852), .Y(n487) );
  oa211d1_hd U1367 ( .A(a[23]), .B(n2280), .C(n2857), .D(n2856), .Y(n488) );
  oa21d1_hd U1368 ( .A(a_e[8]), .B(n2859), .C(n2858), .Y(n2862) );
  scg17d1_hd U1369 ( .A(a_e[9]), .B(n2862), .C(n2861), .D(n2860), .Y(n489) );
  nr2d1_hd U1370 ( .A(n2912), .B(n2911), .Y(n2908) );
  nr2d1_hd U1371 ( .A(n2898), .B(n2897), .Y(n2888) );
  ao21d1_hd U1372 ( .A(n2889), .B(n2864), .C(n2919), .Y(n2887) );
  scg14d1_hd U1373 ( .A(n2865), .B(n2889), .C(n2887), .Y(n2871) );
  ao21d1_hd U1374 ( .A(n2909), .B(n2869), .C(n2871), .Y(n2953) );
  ivd1_hd U1375 ( .A(b[25]), .Y(n2904) );
  nr2d1_hd U1376 ( .A(n2914), .B(n2904), .Y(n2903) );
  ivd1_hd U1377 ( .A(b[27]), .Y(n2891) );
  nr2d1_hd U1378 ( .A(n2900), .B(n2891), .Y(n2890) );
  ivd1_hd U1379 ( .A(b[29]), .Y(n2875) );
  nr2d1_hd U1380 ( .A(n2883), .B(n2875), .Y(n2868) );
  nr2d1_hd U1381 ( .A(n2868), .B(n2280), .Y(n2877) );
  nr2d1_hd U1382 ( .A(n2954), .B(n2864), .Y(n2882) );
  ivd1_hd U1383 ( .A(n2882), .Y(n2881) );
  nr2d1_hd U1384 ( .A(n2865), .B(n2881), .Y(n2870) );
  nd3d1_hd U1385 ( .A(b_e[7]), .B(n2870), .C(n2867), .Y(n2866) );
  oa211d1_hd U1386 ( .A(n2953), .B(n2867), .C(n2955), .D(n2866), .Y(n490) );
  ao22d1_hd U1387 ( .A(b_e[7]), .B(n2871), .C(n2870), .D(n2869), .Y(n2872) );
  oa211d1_hd U1388 ( .A(n2280), .B(n2873), .C(n2872), .D(n2955), .Y(n491) );
  oa21d1_hd U1389 ( .A(b_e[5]), .B(n2954), .C(n2887), .Y(n2878) );
  ao22d1_hd U1390 ( .A(b_e[6]), .B(n2878), .C(n2877), .D(n2876), .Y(n2879) );
  oa211d1_hd U1391 ( .A(n2881), .B(n2880), .C(n2879), .D(n2956), .Y(n492) );
  ao21d1_hd U1392 ( .A(n2882), .B(n2886), .C(n2916), .Y(n2885) );
  oa211d1_hd U1393 ( .A(n2890), .B(b[28]), .C(n2279), .D(n2883), .Y(n2884) );
  oa211d1_hd U1394 ( .A(n2887), .B(n2886), .C(n2885), .D(n2884), .Y(n493) );
  ao21d1_hd U1395 ( .A(n2889), .B(n2897), .C(n2919), .Y(n2899) );
  ao211d1_hd U1396 ( .A(n2900), .B(n2891), .C(n2890), .D(n2280), .Y(n2892) );
  ao21d1_hd U1397 ( .A(n2893), .B(b_e[4]), .C(n2892), .Y(n2894) );
  oa211d1_hd U1398 ( .A(b_e[4]), .B(n2895), .C(n2894), .D(n2956), .Y(n494) );
  oa22d1_hd U1399 ( .A(n2899), .B(n2898), .C(n2897), .D(n2896), .Y(n2902) );
  oa211d1_hd U1400 ( .A(n2903), .B(b[26]), .C(n2279), .D(n2900), .Y(n2901) );
  scg13d1_hd U1401 ( .A(n2902), .B(n2916), .C(n2901), .Y(n495) );
  nr2d1_hd U1402 ( .A(b_e[0]), .B(n2954), .Y(n2918) );
  nr2d1_hd U1403 ( .A(n2919), .B(n2918), .Y(n2913) );
  ao211d1_hd U1404 ( .A(n2914), .B(n2904), .C(n2903), .D(n2280), .Y(n2905) );
  ao211d1_hd U1405 ( .A(b_e[2]), .B(n2906), .C(n2916), .D(n2905), .Y(n2907) );
  scg22d1_hd U1406 ( .A(n2909), .B(n2908), .C(b_e[2]), .D(n2907), .Y(n496) );
  oa22d1_hd U1407 ( .A(n2913), .B(n2912), .C(n2911), .D(n2910), .Y(n2917) );
  oa211d1_hd U1408 ( .A(b[23]), .B(b[24]), .C(n2279), .D(n2914), .Y(n2915) );
  scg13d1_hd U1409 ( .A(n2917), .B(n2916), .C(n2915), .Y(n497) );
  ao21d1_hd U1410 ( .A(n2919), .B(b_e[0]), .C(n2918), .Y(n2920) );
  oa21d1_hd U1411 ( .A(b[23]), .B(n2280), .C(n2920), .Y(n498) );
  scg21d1_hd U1412 ( .A(n2921), .B(o_AB_ACK), .C(i_RST), .D(n27), .Y(n499) );
  oa211d1_hd U1413 ( .A(state[3]), .B(n2926), .C(n2925), .D(n2924), .Y(n2941)
         );
  nd3d1_hd U1414 ( .A(n2281), .B(o_Z_STB), .C(i_Z_ACK), .Y(n2965) );
  nd4d1_hd U1415 ( .A(N41), .B(n2958), .C(n2965), .D(n1284), .Y(n2932) );
  ivd1_hd U1416 ( .A(n2927), .Y(n2929) );
  oa22d1_hd U1417 ( .A(n2930), .B(n2960), .C(n2929), .D(n2928), .Y(n2931) );
  nr4d1_hd U1418 ( .A(n27), .B(n2941), .C(n2932), .D(n2931), .Y(n2933) );
  ivd1_hd U1419 ( .A(n2961), .Y(n2938) );
  nr2d1_hd U1420 ( .A(n2936), .B(n2944), .Y(n2937) );
  ao22d1_hd U1421 ( .A(state[2]), .B(n2938), .C(N41), .D(n2937), .Y(n2939) );
  oa21d1_hd U1422 ( .A(n2940), .B(n2963), .C(n2939), .Y(n500) );
  nr2d1_hd U1423 ( .A(n1291), .B(n2941), .Y(n2943) );
  oa22d1_hd U1424 ( .A(n2943), .B(n2963), .C(n2942), .D(n2961), .Y(n501) );
  ao21d1_hd U1425 ( .A(state[1]), .B(n2944), .C(state[0]), .Y(n2945) );
  nr2d1_hd U1426 ( .A(n2946), .B(n2945), .Y(n2948) );
  oa22d1_hd U1427 ( .A(n2948), .B(n2963), .C(n2947), .D(n2961), .Y(n502) );
  ao22d1_hd U1428 ( .A(b_m[26]), .B(n2949), .C(n2277), .D(b[22]), .Y(n2950) );
  oa21d1_hd U1429 ( .A(n2952), .B(n2275), .C(n2950), .Y(n503) );
  oa21d1_hd U1430 ( .A(b_e[8]), .B(n2954), .C(n2953), .Y(n2957) );
  scg15d1_hd U1431 ( .A(b_e[9]), .B(n2957), .C(n2956), .D(n2955), .Y(n504) );
  oa22d1_hd U1432 ( .A(n2964), .B(n2963), .C(n2962), .D(n2961), .Y(n505) );
  ivd1_hd U1433 ( .A(n2965), .Y(n2966) );
  scg21d1_hd U1434 ( .A(n2281), .B(o_Z_STB), .C(i_RST), .D(n2966), .Y(n506) );
endmodule


module float_adder_0 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3, C91_DATA2_4,
         C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8, n1, n2, n27, n266,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n509, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23, C2_Z_22,
         C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16, C2_Z_15,
         C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8, C2_Z_7,
         C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_43J4_124_6938_n58, DP_OP_43J4_124_6938_n57,
         DP_OP_43J4_124_6938_n56, DP_OP_43J4_124_6938_n55,
         DP_OP_43J4_124_6938_n54, DP_OP_43J4_124_6938_n53,
         DP_OP_43J4_124_6938_n52, DP_OP_43J4_124_6938_n51,
         DP_OP_43J4_124_6938_n50, DP_OP_43J4_124_6938_n49,
         DP_OP_43J4_124_6938_n48, DP_OP_43J4_124_6938_n47,
         DP_OP_43J4_124_6938_n46, DP_OP_43J4_124_6938_n45,
         DP_OP_43J4_124_6938_n44, DP_OP_43J4_124_6938_n43,
         DP_OP_43J4_124_6938_n42, DP_OP_43J4_124_6938_n41,
         DP_OP_43J4_124_6938_n40, DP_OP_43J4_124_6938_n39,
         DP_OP_43J4_124_6938_n38, DP_OP_43J4_124_6938_n37,
         DP_OP_43J4_124_6938_n36, DP_OP_43J4_124_6938_n35,
         DP_OP_43J4_124_6938_n34, DP_OP_43J4_124_6938_n33,
         DP_OP_43J4_124_6938_n32, DP_OP_43J4_124_6938_n27,
         DP_OP_43J4_124_6938_n26, DP_OP_43J4_124_6938_n25,
         DP_OP_43J4_124_6938_n24, DP_OP_43J4_124_6938_n23,
         DP_OP_43J4_124_6938_n22, DP_OP_43J4_124_6938_n21,
         DP_OP_43J4_124_6938_n20, DP_OP_43J4_124_6938_n19,
         DP_OP_43J4_124_6938_n18, DP_OP_43J4_124_6938_n17,
         DP_OP_43J4_124_6938_n16, DP_OP_43J4_124_6938_n15,
         DP_OP_43J4_124_6938_n14, DP_OP_43J4_124_6938_n13,
         DP_OP_43J4_124_6938_n12, DP_OP_43J4_124_6938_n11,
         DP_OP_43J4_124_6938_n10, DP_OP_43J4_124_6938_n9,
         DP_OP_43J4_124_6938_n8, DP_OP_43J4_124_6938_n7,
         DP_OP_43J4_124_6938_n6, DP_OP_43J4_124_6938_n5,
         DP_OP_43J4_124_6938_n4, DP_OP_43J4_124_6938_n3,
         DP_OP_43J4_124_6938_n2, DP_OP_43J4_124_6938_n1,
         DP_OP_154J4_137_6175_n9, DP_OP_154J4_137_6175_n8,
         DP_OP_154J4_137_6175_n7, DP_OP_154J4_137_6175_n6,
         DP_OP_154J4_137_6175_n5, DP_OP_154J4_137_6175_n4,
         DP_OP_154J4_137_6175_n3, DP_OP_154J4_137_6175_n2, n2270, n1222, n1284,
         n1285, n1291, n1891, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J4_137_6175_U10 ( .A(n1291), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J4_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J4_137_6175_U9 ( .A(n1291), .B(z_e[2]), .CI(
        DP_OP_154J4_137_6175_n9), .CO(DP_OP_154J4_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J4_137_6175_U8 ( .A(n1291), .B(z_e[3]), .CI(
        DP_OP_154J4_137_6175_n8), .CO(DP_OP_154J4_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J4_137_6175_U7 ( .A(n1291), .B(z_e[4]), .CI(
        DP_OP_154J4_137_6175_n7), .CO(DP_OP_154J4_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J4_137_6175_U6 ( .A(n1291), .B(z_e[5]), .CI(
        DP_OP_154J4_137_6175_n6), .CO(DP_OP_154J4_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J4_137_6175_U5 ( .A(n1291), .B(z_e[6]), .CI(
        DP_OP_154J4_137_6175_n5), .CO(DP_OP_154J4_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J4_137_6175_U4 ( .A(n1291), .B(z_e[7]), .CI(
        DP_OP_154J4_137_6175_n4), .CO(DP_OP_154J4_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J4_137_6175_U3 ( .A(n1291), .B(z_e[8]), .CI(
        DP_OP_154J4_137_6175_n3), .CO(DP_OP_154J4_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n2286), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n2286), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n509), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n2286), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n2286), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n2286), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n2286), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n2286), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n509), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n509), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n509), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n509), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n2286), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n2286), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n2286), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n2286), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n2286), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n2286), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n2286), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n2286), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n2286), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n509), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n2286), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n2286), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n2286), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n2286), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n2286), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n2286), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n2286), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n2286), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n2286), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n2287), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n2287), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n2287), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n2287), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n2273), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n2273), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n2287), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n2287), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n2287), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n2287), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n2287), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n27), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n2287), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n2287), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n2287), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n27), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n27), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n27), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n27), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n27), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n27), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n2287), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n27), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n2287), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n2287), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n27), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n27), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n2287), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n2287), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n2287), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n2287), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n2287), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n2287), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n2287), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n2287), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n2287), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n2287), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n2287), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n2287), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n2287), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n2287), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n2287), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n2287), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n2287), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n2287), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n2287), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n2287), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n2287), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n2287), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n2287), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n2287), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n2287), .CK(i_CLK), .Q(b[22]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n2273), .CK(i_CLK), .Q(sum[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n2273), .CK(i_CLK), .Q(sum[2]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n2273), .CK(i_CLK), .Q(sum[26]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n2273), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n2273), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n2273), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n2273), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n2273), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n2273), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n2273), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n2273), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n2273), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n2273), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n2273), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n2273), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n2273), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n2273), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n2273), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n2273), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n2273), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n2273), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n2273), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n2273), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n2273), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n2273), .CK(i_CLK), .Q(sum[25]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n2273), .CK(i_CLK), .Q(sum[1]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n2287), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n2287), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n2287), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n2287), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n2273), .CK(i_CLK), .Q(sum[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n2287), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n2287), .CK(i_CLK), .Q(b[28]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n2287), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n2287), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n2287), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n2287), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n2287), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n2287), .CK(i_CLK), .Q(b[26]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n2287), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n2287), .CK(i_CLK), .Q(b[23]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n1222), .CK(i_CLK), .Q(guard) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n2282), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n2282), .CK(i_CLK), .Q(a_s) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n2270), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n2270), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J4_124_6938_U28 ( .A(C2_Z_0), .B(n1891), .CI(
        DP_OP_43J4_124_6938_n58), .CO(DP_OP_43J4_124_6938_n27), .S(N310) );
  fad1_hd DP_OP_43J4_124_6938_U27 ( .A(DP_OP_43J4_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J4_124_6938_n27), .CO(DP_OP_43J4_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J4_124_6938_U26 ( .A(DP_OP_43J4_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J4_124_6938_n26), .CO(DP_OP_43J4_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J4_124_6938_U25 ( .A(DP_OP_43J4_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J4_124_6938_n25), .CO(DP_OP_43J4_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J4_124_6938_U2 ( .A(DP_OP_43J4_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J4_124_6938_n2), .CO(DP_OP_43J4_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J4_124_6938_U16 ( .A(DP_OP_43J4_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J4_124_6938_n16), .CO(DP_OP_43J4_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J4_124_6938_U17 ( .A(DP_OP_43J4_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J4_124_6938_n17), .CO(DP_OP_43J4_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J4_124_6938_U18 ( .A(DP_OP_43J4_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J4_124_6938_n18), .CO(DP_OP_43J4_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J4_124_6938_U19 ( .A(DP_OP_43J4_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J4_124_6938_n19), .CO(DP_OP_43J4_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J4_124_6938_U20 ( .A(DP_OP_43J4_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J4_124_6938_n20), .CO(DP_OP_43J4_124_6938_n19), .S(N318)
         );
  fad1_hd DP_OP_43J4_124_6938_U21 ( .A(DP_OP_43J4_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J4_124_6938_n21), .CO(DP_OP_43J4_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J4_124_6938_U22 ( .A(DP_OP_43J4_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J4_124_6938_n22), .CO(DP_OP_43J4_124_6938_n21), .S(N316)
         );
  fad1_hd DP_OP_43J4_124_6938_U23 ( .A(DP_OP_43J4_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J4_124_6938_n23), .CO(DP_OP_43J4_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J4_124_6938_U24 ( .A(DP_OP_43J4_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J4_124_6938_n24), .CO(DP_OP_43J4_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J4_124_6938_U15 ( .A(DP_OP_43J4_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J4_124_6938_n15), .CO(DP_OP_43J4_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J4_124_6938_U14 ( .A(DP_OP_43J4_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J4_124_6938_n14), .CO(DP_OP_43J4_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J4_124_6938_U13 ( .A(DP_OP_43J4_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J4_124_6938_n13), .CO(DP_OP_43J4_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J4_124_6938_U12 ( .A(DP_OP_43J4_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J4_124_6938_n12), .CO(DP_OP_43J4_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J4_124_6938_U5 ( .A(DP_OP_43J4_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J4_124_6938_n5), .CO(DP_OP_43J4_124_6938_n4), .S(N333) );
  fad1_hd DP_OP_43J4_124_6938_U4 ( .A(DP_OP_43J4_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J4_124_6938_n4), .CO(DP_OP_43J4_124_6938_n3), .S(N334) );
  fad1_hd DP_OP_43J4_124_6938_U3 ( .A(DP_OP_43J4_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J4_124_6938_n3), .CO(DP_OP_43J4_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J4_124_6938_U11 ( .A(DP_OP_43J4_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J4_124_6938_n11), .CO(DP_OP_43J4_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J4_124_6938_U10 ( .A(DP_OP_43J4_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J4_124_6938_n10), .CO(DP_OP_43J4_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J4_124_6938_U9 ( .A(DP_OP_43J4_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J4_124_6938_n9), .CO(DP_OP_43J4_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J4_124_6938_U8 ( .A(DP_OP_43J4_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J4_124_6938_n8), .CO(DP_OP_43J4_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J4_124_6938_U7 ( .A(DP_OP_43J4_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J4_124_6938_n7), .CO(DP_OP_43J4_124_6938_n6), .S(N331) );
  fad1_hd DP_OP_43J4_124_6938_U6 ( .A(DP_OP_43J4_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J4_124_6938_n6), .CO(DP_OP_43J4_124_6938_n5), .S(N332) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  clknd2d1_hd U523 ( .A(a_m[24]), .B(n2703), .Y(n2326) );
  clknd2d1_hd U524 ( .A(a_m[7]), .B(n2737), .Y(n2296) );
  clknd2d1_hd U525 ( .A(a_m[11]), .B(n2729), .Y(n2303) );
  clknd2d1_hd U526 ( .A(a_e[3]), .B(n2903), .Y(n2396) );
  clknd2d1_hd U527 ( .A(b_e[6]), .B(n2808), .Y(n2399) );
  clknd2d1_hd U528 ( .A(b_m[19]), .B(n2761), .Y(n2316) );
  clknd2d1_hd U529 ( .A(a_m[18]), .B(n2715), .Y(n2314) );
  clknd2d1_hd U530 ( .A(n2386), .B(n2399), .Y(n2392) );
  clknd2d1_hd U531 ( .A(z_e[7]), .B(z_e[8]), .Y(n2506) );
  clknd2d1_hd U532 ( .A(b_e[0]), .B(n2843), .Y(n2387) );
  clknd2d1_hd U533 ( .A(b_e[4]), .B(n2893), .Y(n2869) );
  clknd2d1_hd U534 ( .A(b_e[6]), .B(b_e[5]), .Y(n2870) );
  clknd2d1_hd U535 ( .A(n2894), .B(n2411), .Y(n2933) );
  ad2bd1_hd U536 ( .B(n2519), .AN(n1222), .Y(n2640) );
  clknd2d1_hd U537 ( .A(n2662), .B(n2517), .Y(n2518) );
  clknd2d1_hd U538 ( .A(n2420), .B(n2418), .Y(n2439) );
  clknd2d1_hd U539 ( .A(n2432), .B(n2477), .Y(n2507) );
  clknd2d1_hd U540 ( .A(n2868), .B(n2417), .Y(n2415) );
  clknd2d1_hd U541 ( .A(n2802), .B(n2419), .Y(n2455) );
  clknd2d1_hd U542 ( .A(n2952), .B(n2947), .Y(n2672) );
  clknd2d1_hd U543 ( .A(a_e[2]), .B(n2846), .Y(n2806) );
  clknd2d1_hd U544 ( .A(state[0]), .B(n2947), .Y(n2931) );
  clknd2d1_hd U545 ( .A(z_m[19]), .B(z_m[20]), .Y(n2674) );
  clknd2d1_hd U546 ( .A(n2280), .B(n2894), .Y(n2747) );
  clknd2d1_hd U547 ( .A(n2278), .B(n2894), .Y(n2795) );
  clknd2d1_hd U548 ( .A(n2410), .B(n2952), .Y(n2413) );
  clknd2d1_hd U549 ( .A(n2845), .B(n2843), .Y(n2862) );
  clknd2d1_hd U550 ( .A(b_e[2]), .B(n2913), .Y(n2902) );
  clknd2d1_hd U551 ( .A(n2914), .B(n2903), .Y(n2901) );
  clknd2d1_hd U552 ( .A(n2829), .B(n2805), .Y(n2814) );
  clknd2d1_hd U553 ( .A(n2821), .B(n2817), .Y(n2865) );
  clknd2d1_hd U554 ( .A(n2895), .B(b[28]), .Y(n2888) );
  clknd2d1_hd U555 ( .A(n2410), .B(n2941), .Y(n2945) );
  clknd2d1_hd U556 ( .A(state[2]), .B(n2967), .Y(n2949) );
  clknd2d1_hd U557 ( .A(N41), .B(n2966), .Y(n2968) );
  clknd2d1_hd U558 ( .A(n2665), .B(n2655), .Y(n2646) );
  clknd2d1_hd U559 ( .A(z_m[0]), .B(n2665), .Y(n2638) );
  clknd2d1_hd U560 ( .A(n2651), .B(n2646), .Y(n2641) );
  clknd2d1_hd U561 ( .A(n2614), .B(n2665), .Y(n2621) );
  clknd2d1_hd U562 ( .A(n2590), .B(n2665), .Y(n2597) );
  clknd2d1_hd U563 ( .A(z_m[21]), .B(n2675), .Y(n2667) );
  clknd2d1_hd U564 ( .A(n2681), .B(sum[27]), .Y(n2679) );
  clknd2d1_hd U565 ( .A(n2567), .B(n2665), .Y(n2573) );
  clknd2d1_hd U566 ( .A(n2539), .B(n2665), .Y(n2546) );
  clknd2d1_hd U567 ( .A(z_m[15]), .B(z_m[16]), .Y(n2553) );
  clknd2d1_hd U568 ( .A(n2520), .B(n2535), .Y(n2668) );
  clknd2d1_hd U569 ( .A(n2808), .B(n2879), .Y(n2448) );
  clknd2d1_hd U570 ( .A(a_e[0]), .B(b_e[0]), .Y(n2489) );
  clknd2d1_hd U571 ( .A(n2482), .B(n2477), .Y(n2476) );
  clknd2d1_hd U572 ( .A(n2468), .B(n2464), .Y(n2463) );
  clknd2d1_hd U573 ( .A(a_e[7]), .B(b_e[7]), .Y(n2443) );
  clknd2d1_hd U574 ( .A(n2454), .B(n2450), .Y(n2449) );
  clknd2d1_hd U575 ( .A(n2493), .B(n2440), .Y(n2492) );
  ivd1_hd U576 ( .A(b_m[1]), .Y(n2748) );
  clknd2d1_hd U577 ( .A(n2364), .B(n1891), .Y(n2356) );
  ivd1_hd U578 ( .A(b_m[2]), .Y(n2746) );
  clknd2d1_hd U579 ( .A(n2508), .B(n2433), .Y(n2440) );
  clknd2d1_hd U580 ( .A(n2431), .B(n2430), .Y(n2434) );
  nid1_hd U581 ( .A(n2503), .Y(n2275) );
  ivd2_hd U582 ( .A(n2356), .Y(n2361) );
  ivd2_hd U583 ( .A(n2362), .Y(n1891) );
  clknd2d1_hd U584 ( .A(n2329), .B(a_m[26]), .Y(n2330) );
  nr2d1_hd U585 ( .A(n2329), .B(a_m[26]), .Y(n2331) );
  ivd4_hd U586 ( .A(n2364), .Y(n2274) );
  clknd2d1_hd U587 ( .A(state[1]), .B(n2952), .Y(n2928) );
  clknd2d1_hd U588 ( .A(a[23]), .B(a[24]), .Y(n2856) );
  clknd2d1_hd U589 ( .A(n2844), .B(n2862), .Y(n2854) );
  clknd2d1_hd U590 ( .A(a_e[3]), .B(n2838), .Y(n2836) );
  clknd2d1_hd U591 ( .A(n2847), .B(a[26]), .Y(n2840) );
  clknd2d1_hd U592 ( .A(b[23]), .B(b[24]), .Y(n2919) );
  clknd2d1_hd U593 ( .A(n2914), .B(n2917), .Y(n2915) );
  clknd2d1_hd U594 ( .A(a_e[5]), .B(n2824), .Y(n2823) );
  clknd2d1_hd U595 ( .A(n2844), .B(n2894), .Y(n2864) );
  clknd2d1_hd U596 ( .A(a_e[4]), .B(a_e[3]), .Y(n2804) );
  clknd2d1_hd U597 ( .A(n2831), .B(a[28]), .Y(n2825) );
  clknd2d1_hd U598 ( .A(n2908), .B(b[26]), .Y(n2905) );
  clknd2d1_hd U599 ( .A(n2904), .B(n2901), .Y(n2898) );
  clknd2d1_hd U600 ( .A(n2510), .B(n2509), .Y(n393) );
  clknd2d1_hd U601 ( .A(b[30]), .B(n2873), .Y(n2878) );
  clknd2d1_hd U602 ( .A(a_e[0]), .B(n2860), .Y(n2861) );
  clknd2d1_hd U603 ( .A(n2284), .B(n2811), .Y(n2816) );
  clknd2d1_hd U604 ( .A(b_e[5]), .B(n2879), .Y(n2885) );
  clknd2d1_hd U605 ( .A(n2888), .B(n2880), .Y(n2881) );
  clknd2d1_hd U606 ( .A(n2666), .B(n2646), .Y(n2648) );
  clknd2d1_hd U607 ( .A(n2701), .B(n2700), .Y(n428) );
  clknd2d1_hd U608 ( .A(DP_OP_154J4_137_6175_n2), .B(n2699), .Y(n2697) );
  clknd2d1_hd U609 ( .A(n2658), .B(z_m[14]), .Y(n2562) );
  clknd2d1_hd U610 ( .A(n2680), .B(n2513), .Y(n1222) );
  clknd2d1_hd U611 ( .A(n2658), .B(z_m[15]), .Y(n2555) );
  clknd2d1_hd U612 ( .A(n2491), .B(n2446), .Y(n362) );
  clknd2d1_hd U613 ( .A(n2498), .B(n2497), .Y(n2499) );
  clknd2d1_hd U614 ( .A(n2918), .B(n2915), .Y(n2911) );
  clknd2d1_hd U615 ( .A(n2825), .B(n2818), .Y(n2820) );
  clknd2d1_hd U616 ( .A(n2914), .B(n2893), .Y(n2900) );
  oa22ad1_hd U617 ( .A(n2328), .B(b_m[25]), .C(n2327), .D(a_m[25]), .Y(n2329)
         );
  ivd1_hd U618 ( .A(b_m[23]), .Y(n2705) );
  ivd1_hd U619 ( .A(b_m[3]), .Y(n2745) );
  ivd1_hd U620 ( .A(a_m[24]), .Y(n2751) );
  ivd1_hd U621 ( .A(b_m[21]), .Y(n2709) );
  nr2d1_hd U622 ( .A(n2327), .B(a_m[25]), .Y(n2328) );
  ao22d1_hd U623 ( .A(b_m[24]), .B(n2751), .C(n2326), .D(n2325), .Y(n2327) );
  oa22d1_hd U624 ( .A(a_m[23]), .B(n2705), .C(n2324), .D(n2323), .Y(n2325) );
  nr2d1_hd U625 ( .A(n2322), .B(n2321), .Y(n2324) );
  ao21d1_hd U626 ( .A(n2709), .B(a_m[21]), .C(n2320), .Y(n2321) );
  ivd3_hd U627 ( .A(n1284), .Y(n2273) );
  oa22d2_hd U628 ( .A(n2437), .B(n2421), .C(b_s), .D(a_s), .Y(n2362) );
  xo2d1_hd U629 ( .A(n1891), .B(DP_OP_43J4_124_6938_n1), .Y(N337) );
  oa211d8_hd U630 ( .A(b_m[26]), .B(n2331), .C(n1891), .D(n2330), .Y(n2364) );
  nid4_hd U631 ( .A(n27), .Y(n2287) );
  ad3d1_hd U632 ( .A(n2852), .B(n2846), .C(n2845), .Y(n2850) );
  scg6d1_hd U633 ( .A(b_m[17]), .B(n2315), .C(n2765), .Y(n2313) );
  scg6d1_hd U634 ( .A(b_m[10]), .B(n2304), .C(n2779), .Y(n2302) );
  scg9d1_hd U635 ( .A(n2963), .B(n2520), .C(n2533), .Y(n2524) );
  scg9d1_hd U636 ( .A(n2945), .B(n2411), .C(n2285), .Y(n2956) );
  ad3d1_hd U637 ( .A(n2965), .B(n2281), .C(n2963), .Y(n2969) );
  scg6d1_hd U638 ( .A(b_m[6]), .B(n2297), .C(n2787), .Y(n2295) );
  scg10d1_hd U639 ( .A(n2420), .B(n2419), .C(n2418), .D(n2417), .Y(n2497) );
  ivd2_hd U640 ( .A(n2679), .Y(n2653) );
  ad2d1_hd U641 ( .A(n2935), .B(n2516), .Y(n2512) );
  ivd2_hd U642 ( .A(n1285), .Y(n2285) );
  or2d1_hd U643 ( .A(n2949), .B(n2672), .Y(n1284) );
  or2d1_hd U644 ( .A(state[2]), .B(n2967), .Y(n2927) );
  ivd1_hd U645 ( .A(b_m[0]), .Y(n2749) );
  nr2ad1_hd U646 ( .A(n2963), .B(n2640), .Y(n2665) );
  nr2d2_hd U647 ( .A(n2494), .B(n2929), .Y(n2504) );
  nr2ad1_hd U648 ( .A(n2683), .B(n2695), .Y(n2698) );
  nr2ad1_hd U649 ( .A(n2965), .B(n2640), .Y(n2647) );
  nr2ad1_hd U650 ( .A(n2928), .B(n2949), .Y(n1291) );
  oa22ad1_hd U651 ( .A(n2301), .B(a_m[9]), .C(n2300), .D(b_m[9]), .Y(n2304) );
  oa22ad1_hd U652 ( .A(n2294), .B(a_m[5]), .C(n2293), .D(b_m[5]), .Y(n2297) );
  ivd1_hd U653 ( .A(b_m[4]), .Y(n2743) );
  ivd1_hd U654 ( .A(a_m[4]), .Y(n2791) );
  ivd1_hd U655 ( .A(a_m[3]), .Y(n2793) );
  nid2_hd U656 ( .A(n2964), .Y(n2281) );
  ivd1_hd U657 ( .A(n2665), .Y(n2639) );
  ivd1_hd U658 ( .A(n2693), .Y(n2695) );
  ivd1_hd U659 ( .A(n2801), .Y(n2279) );
  ivd1_hd U660 ( .A(n2945), .Y(n2894) );
  ivd1_hd U661 ( .A(b_m[7]), .Y(n2737) );
  ivd1_hd U662 ( .A(b_m[8]), .Y(n2735) );
  nid2_hd U663 ( .A(n2505), .Y(n2276) );
  ivd1_hd U664 ( .A(n2658), .Y(n2666) );
  nr2d1_hd U665 ( .A(n2939), .B(n2640), .Y(n2658) );
  ivd1_hd U666 ( .A(n2682), .Y(n2963) );
  nid2_hd U667 ( .A(n2652), .Y(n2277) );
  ivd1_hd U668 ( .A(n2647), .Y(n2654) );
  ivd1_hd U669 ( .A(n2681), .Y(n2513) );
  ivd1_hd U670 ( .A(n2285), .Y(n2282) );
  ivd2_hd U671 ( .A(n2795), .Y(n2798) );
  nr2d1_hd U672 ( .A(n2927), .B(n2672), .Y(n2682) );
  ivd2_hd U673 ( .A(n2956), .Y(n2280) );
  ivd2_hd U674 ( .A(n2279), .Y(n2278) );
  oa21d1_hd U675 ( .A(n2932), .B(n2933), .C(n2285), .Y(n2801) );
  nr2d1_hd U676 ( .A(n2423), .B(n2930), .Y(n2951) );
  ivd1_hd U677 ( .A(n2270), .Y(n2930) );
  ivd1_hd U678 ( .A(n2285), .Y(n2284) );
  ivd1_hd U679 ( .A(b_m[15]), .Y(n2721) );
  ivd1_hd U680 ( .A(b_m[14]), .Y(n2723) );
  ivd1_hd U681 ( .A(b_m[13]), .Y(n2725) );
  ivd1_hd U682 ( .A(a_m[12]), .Y(n2775) );
  ivd1_hd U683 ( .A(b_m[16]), .Y(n2719) );
  ivd1_hd U684 ( .A(b_m[18]), .Y(n2715) );
  ivd1_hd U685 ( .A(b_m[24]), .Y(n2703) );
  nid2_hd U686 ( .A(n509), .Y(n2286) );
  ivd1_hd U687 ( .A(n2493), .Y(n2929) );
  ad3d1_hd U688 ( .A(n2926), .B(i_AB_STB), .C(o_AB_ACK), .Y(n27) );
  ivd2_hd U689 ( .A(n2747), .Y(n2954) );
  ivd1_hd U690 ( .A(n2500), .Y(n2484) );
  nr2d1_hd U691 ( .A(n2931), .B(n2927), .Y(n2493) );
  ivd1_hd U692 ( .A(n2516), .Y(n2965) );
  ivd2_hd U693 ( .A(n2285), .Y(n2283) );
  ivd1_hd U694 ( .A(n1291), .Y(n2939) );
  nr2d1_hd U695 ( .A(n2931), .B(n2949), .Y(n2681) );
  nr2bd1_hd U696 ( .AN(n2941), .B(n2949), .Y(n2516) );
  nr2bd1_hd U697 ( .AN(z_e[1]), .B(n2506), .Y(n2508) );
  ivd1_hd U698 ( .A(n2866), .Y(n2858) );
  ivd1_hd U699 ( .A(n2914), .Y(n2959) );
  nr2d1_hd U700 ( .A(n2924), .B(n2945), .Y(n2914) );
  ao21d1_hd U701 ( .A(n2868), .B(n2951), .C(n2280), .Y(n2924) );
  ivd1_hd U702 ( .A(n2860), .Y(n2844) );
  ao21d1_hd U703 ( .A(n2802), .B(n2951), .C(n2278), .Y(n2860) );
  ivd1_hd U704 ( .A(b_e[7]), .Y(n2874) );
  ivd1_hd U705 ( .A(a_e[6]), .Y(n2808) );
  ivd1_hd U706 ( .A(a_e[5]), .Y(n2828) );
  ivd1_hd U707 ( .A(b_e[1]), .Y(n2917) );
  nr2d1_hd U708 ( .A(n2947), .B(n2413), .Y(n2270) );
  ivd1_hd U709 ( .A(b_e[8]), .Y(n2872) );
  ivd1_hd U710 ( .A(n2455), .Y(n2416) );
  ivd1_hd U711 ( .A(n2496), .Y(n2420) );
  ivd1_hd U712 ( .A(a_e[4]), .Y(n2807) );
  ivd1_hd U713 ( .A(a_e[0]), .Y(n2843) );
  nr2d1_hd U714 ( .A(n2952), .B(n2947), .Y(n2941) );
  ivd1_hd U715 ( .A(state[0]), .Y(n2952) );
  nr2bd1_hd U716 ( .AN(n2410), .B(n2931), .Y(n1285) );
  ivd1_hd U717 ( .A(state[1]), .Y(n2947) );
  ivd1_hd U718 ( .A(a_m[23]), .Y(n2753) );
  ivd1_hd U719 ( .A(a_m[22]), .Y(n2755) );
  ivd1_hd U720 ( .A(b_m[19]), .Y(n2713) );
  ivd1_hd U721 ( .A(b_m[20]), .Y(n2711) );
  ivd1_hd U722 ( .A(a_m[20]), .Y(n2759) );
  ivd1_hd U723 ( .A(b_m[22]), .Y(n2707) );
  ivd1_hd U724 ( .A(n2951), .Y(n2412) );
  ivd1_hd U725 ( .A(z_m[1]), .Y(n2655) );
  ivd1_hd U726 ( .A(z_m[14]), .Y(n2572) );
  ivd1_hd U727 ( .A(n2640), .Y(n2661) );
  nr4d1_hd U728 ( .A(n2496), .B(n2416), .C(n2415), .D(n2930), .Y(n2503) );
  oa21d1_hd U729 ( .A(n2940), .B(n2939), .C(n2938), .Y(n2966) );
  nr2d1_hd U730 ( .A(n2928), .B(n2927), .Y(n509) );
  ivd1_hd U731 ( .A(z_m[19]), .Y(n2544) );
  nr2d1_hd U732 ( .A(n2281), .B(n2930), .Y(n2500) );
  ao22d1_hd U733 ( .A(n2494), .B(n2493), .C(n2270), .D(n2439), .Y(n2491) );
  scg20d1_hd U734 ( .A(z_e[7]), .B(z_e[8]), .C(z_e[9]), .Y(n2494) );
  ivd1_hd U735 ( .A(z_m[22]), .Y(n2664) );
  ivd1_hd U736 ( .A(round_bit), .Y(n2517) );
  ivd1_hd U737 ( .A(z_m[0]), .Y(n2662) );
  ivd1_hd U738 ( .A(n2921), .Y(n2961) );
  ivd1_hd U739 ( .A(z_m[12]), .Y(n2583) );
  ivd1_hd U740 ( .A(z_m[11]), .Y(n2595) );
  ivd1_hd U741 ( .A(z_m[7]), .Y(n2619) );
  ivd1_hd U742 ( .A(z_m[8]), .Y(n2607) );
  ivd1_hd U743 ( .A(z_m[3]), .Y(n2645) );
  ivd1_hd U744 ( .A(z_m[4]), .Y(n2631) );
  ivd1_hd U745 ( .A(z_m[23]), .Y(n2675) );
  ivd1_hd U746 ( .A(state[3]), .Y(n2967) );
  ivd1_hd U747 ( .A(z_e[2]), .Y(n2477) );
  ivd1_hd U748 ( .A(z_e[0]), .Y(n2694) );
  nr2d1_hd U749 ( .A(n2924), .B(n2930), .Y(n2921) );
  ivd1_hd U750 ( .A(n2864), .Y(n2845) );
  ivd1_hd U751 ( .A(a_e[7]), .Y(n2812) );
  ivd1_hd U752 ( .A(b_e[3]), .Y(n2903) );
  nr4d1_hd U753 ( .A(n2409), .B(n2391), .C(n2392), .D(n2390), .Y(n2932) );
  ivd1_hd U754 ( .A(a_e[2]), .Y(n2852) );
  nr2d1_hd U755 ( .A(b_e[9]), .B(n2385), .Y(n2409) );
  scg13d1_hd U756 ( .A(n2439), .B(n2416), .C(n2415), .Y(n2423) );
  ivd1_hd U757 ( .A(b_e[0]), .Y(n2916) );
  ivd1_hd U758 ( .A(b_e[5]), .Y(n2891) );
  ivd1_hd U759 ( .A(b_e[6]), .Y(n2879) );
  ivd1_hd U760 ( .A(a_e[3]), .Y(n2837) );
  ivd1_hd U761 ( .A(a_e[9]), .Y(n2385) );
  ivd1_hd U762 ( .A(a_e[8]), .Y(n2810) );
  ivd1_hd U763 ( .A(a_e[1]), .Y(n2803) );
  nr2d1_hd U764 ( .A(state[2]), .B(state[3]), .Y(n2410) );
  ivd1_hd U765 ( .A(a[30]), .Y(n2817) );
  ivd1_hd U766 ( .A(a_m[0]), .Y(n2797) );
  ivd1_hd U767 ( .A(a_m[1]), .Y(n2796) );
  ivd1_hd U768 ( .A(a_m[2]), .Y(n2794) );
  ivd1_hd U769 ( .A(b_m[5]), .Y(n2741) );
  ivd1_hd U770 ( .A(a_m[5]), .Y(n2789) );
  ivd1_hd U771 ( .A(b_m[6]), .Y(n2739) );
  ivd1_hd U772 ( .A(b_m[9]), .Y(n2733) );
  ivd1_hd U773 ( .A(a_m[9]), .Y(n2781) );
  ivd1_hd U774 ( .A(b_m[10]), .Y(n2731) );
  ivd1_hd U775 ( .A(b_m[12]), .Y(n2727) );
  ivd1_hd U776 ( .A(a_m[14]), .Y(n2771) );
  ivd1_hd U777 ( .A(b_m[17]), .Y(n2717) );
  ivd1_hd U778 ( .A(a_m[18]), .Y(n2763) );
  ivd1_hd U779 ( .A(a_m[21]), .Y(n2757) );
  ivd1_hd U780 ( .A(b_m[25]), .Y(n2957) );
  ivd1_hd U781 ( .A(a_m[19]), .Y(n2761) );
  ivd1_hd U782 ( .A(a_m[17]), .Y(n2765) );
  ivd1_hd U783 ( .A(a_m[13]), .Y(n2773) );
  ivd1_hd U784 ( .A(a_m[10]), .Y(n2779) );
  ivd1_hd U785 ( .A(b_m[11]), .Y(n2729) );
  ivd1_hd U786 ( .A(a_m[6]), .Y(n2787) );
  ivd1_hd U787 ( .A(a_m[8]), .Y(n2783) );
  ivd1_hd U788 ( .A(a_m[7]), .Y(n2785) );
  ivd1_hd U789 ( .A(a_m[11]), .Y(n2777) );
  ivd1_hd U790 ( .A(a_m[16]), .Y(n2767) );
  ivd1_hd U791 ( .A(a_m[15]), .Y(n2769) );
  ivd1_hd U792 ( .A(b_s), .Y(n2421) );
  ivd1_hd U793 ( .A(a_s), .Y(n2437) );
  nr2d1_hd U794 ( .A(state[1]), .B(n2413), .Y(n2926) );
  nr2d1_hd U795 ( .A(sum[27]), .B(n2513), .Y(n2652) );
  nd2bd1_hd U796 ( .AN(b[30]), .B(n2882), .Y(n2960) );
  nr2d1_hd U797 ( .A(n2930), .B(n2860), .Y(n2866) );
  nd2bd1_hd U798 ( .AN(n2409), .B(n2408), .Y(n2411) );
  ivd1_hd U799 ( .A(b_e[9]), .Y(n2405) );
  ivd1_hd U800 ( .A(a_m[25]), .Y(n2800) );
  oa22d1_hd U801 ( .A(a_m[21]), .B(n2709), .C(a_m[22]), .D(n2707), .Y(n2322)
         );
  ao22d1_hd U802 ( .A(a_m[20]), .B(n2711), .C(a_m[19]), .D(n2713), .Y(n2319)
         );
  ao22d1_hd U803 ( .A(b_m[15]), .B(n2769), .C(b_m[16]), .D(n2767), .Y(n2312)
         );
  ao22d1_hd U804 ( .A(b_m[11]), .B(n2777), .C(b_m[12]), .D(n2775), .Y(n2307)
         );
  ao22d1_hd U805 ( .A(b_m[7]), .B(n2785), .C(b_m[8]), .D(n2783), .Y(n2299) );
  ao22d1_hd U806 ( .A(b_m[3]), .B(n2793), .C(b_m[4]), .D(n2791), .Y(n2292) );
  ao211d1_hd U807 ( .A(a_m[1]), .B(n2748), .C(a_m[0]), .D(n2749), .Y(n2290) );
  oa22d1_hd U808 ( .A(a_m[1]), .B(n2748), .C(a_m[2]), .D(n2746), .Y(n2289) );
  ao22d1_hd U809 ( .A(a_m[3]), .B(n2745), .C(a_m[2]), .D(n2746), .Y(n2288) );
  oa21d1_hd U810 ( .A(n2290), .B(n2289), .C(n2288), .Y(n2291) );
  ao22d1_hd U811 ( .A(a_m[4]), .B(n2743), .C(n2292), .D(n2291), .Y(n2293) );
  nr2d1_hd U812 ( .A(n2293), .B(b_m[5]), .Y(n2294) );
  oa211d1_hd U813 ( .A(b_m[6]), .B(n2297), .C(n2296), .D(n2295), .Y(n2298) );
  ao22d1_hd U814 ( .A(a_m[8]), .B(n2735), .C(n2299), .D(n2298), .Y(n2300) );
  nr2d1_hd U815 ( .A(n2300), .B(b_m[9]), .Y(n2301) );
  oa211d1_hd U816 ( .A(b_m[10]), .B(n2304), .C(n2303), .D(n2302), .Y(n2306) );
  oa22d1_hd U817 ( .A(b_m[13]), .B(n2773), .C(b_m[12]), .D(n2775), .Y(n2305)
         );
  ao21d1_hd U818 ( .A(n2307), .B(n2306), .C(n2305), .Y(n2310) );
  oa22d1_hd U819 ( .A(a_m[13]), .B(n2725), .C(a_m[14]), .D(n2723), .Y(n2309)
         );
  ao22d1_hd U820 ( .A(a_m[15]), .B(n2721), .C(a_m[14]), .D(n2723), .Y(n2308)
         );
  oa21d1_hd U821 ( .A(n2310), .B(n2309), .C(n2308), .Y(n2311) );
  ao22d1_hd U822 ( .A(a_m[16]), .B(n2719), .C(n2312), .D(n2311), .Y(n2315) );
  oa211d1_hd U823 ( .A(b_m[17]), .B(n2315), .C(n2314), .D(n2313), .Y(n2317) );
  oa211d1_hd U824 ( .A(a_m[18]), .B(n2715), .C(n2317), .D(n2316), .Y(n2318) );
  ao22d1_hd U825 ( .A(b_m[20]), .B(n2759), .C(n2319), .D(n2318), .Y(n2320) );
  oa22d1_hd U826 ( .A(b_m[22]), .B(n2755), .C(b_m[23]), .D(n2753), .Y(n2323)
         );
  ao22d1_hd U827 ( .A(n2274), .B(n2749), .C(n2797), .D(n2364), .Y(C2_Z_0) );
  ao22d1_hd U828 ( .A(n2274), .B(n2748), .C(n2796), .D(n2364), .Y(C2_Z_1) );
  ao22d1_hd U829 ( .A(n2274), .B(n2731), .C(n2779), .D(n2364), .Y(C2_Z_10) );
  ao22d1_hd U830 ( .A(n2274), .B(n2729), .C(n2777), .D(n2364), .Y(C2_Z_11) );
  ao22d1_hd U831 ( .A(n2274), .B(n2727), .C(n2775), .D(n2364), .Y(C2_Z_12) );
  ao22d1_hd U832 ( .A(n2274), .B(n2725), .C(n2773), .D(n2364), .Y(C2_Z_13) );
  ao22d1_hd U833 ( .A(n2274), .B(n2723), .C(n2771), .D(n2364), .Y(C2_Z_14) );
  ao22d1_hd U834 ( .A(n2274), .B(n2721), .C(n2769), .D(n2364), .Y(C2_Z_15) );
  ao22d1_hd U835 ( .A(n2274), .B(n2719), .C(n2767), .D(n2364), .Y(C2_Z_16) );
  ao22d1_hd U836 ( .A(n2274), .B(n2717), .C(n2765), .D(n2364), .Y(C2_Z_17) );
  ao22d1_hd U837 ( .A(n2274), .B(n2715), .C(n2763), .D(n2364), .Y(C2_Z_18) );
  ao22d1_hd U838 ( .A(n2274), .B(n2713), .C(n2761), .D(n2364), .Y(C2_Z_19) );
  ao22d1_hd U839 ( .A(n2274), .B(n2746), .C(n2794), .D(n2364), .Y(C2_Z_2) );
  ao22d1_hd U840 ( .A(n2274), .B(n2711), .C(n2759), .D(n2364), .Y(C2_Z_20) );
  ao22d1_hd U841 ( .A(n2274), .B(n2709), .C(n2757), .D(n2364), .Y(C2_Z_21) );
  ao22d1_hd U842 ( .A(n2274), .B(n2707), .C(n2755), .D(n2364), .Y(C2_Z_22) );
  ao22d1_hd U843 ( .A(n2274), .B(n2705), .C(n2753), .D(n2364), .Y(C2_Z_23) );
  ao22d1_hd U844 ( .A(n2274), .B(n2703), .C(n2751), .D(n2364), .Y(C2_Z_24) );
  ao22d1_hd U845 ( .A(n2274), .B(n2957), .C(n2800), .D(n2364), .Y(C2_Z_25) );
  ivd1_hd U846 ( .A(b_m[26]), .Y(n2333) );
  ivd1_hd U847 ( .A(a_m[26]), .Y(n2332) );
  oa21d1_hd U848 ( .A(n2333), .B(n2362), .C(n2332), .Y(C2_Z_26) );
  ao22d1_hd U849 ( .A(n2274), .B(n2745), .C(n2793), .D(n2364), .Y(C2_Z_3) );
  ao22d1_hd U850 ( .A(n2274), .B(n2743), .C(n2791), .D(n2364), .Y(C2_Z_4) );
  ao22d1_hd U851 ( .A(n2274), .B(n2741), .C(n2789), .D(n2364), .Y(C2_Z_5) );
  ao22d1_hd U852 ( .A(n2274), .B(n2739), .C(n2787), .D(n2364), .Y(C2_Z_6) );
  ao22d1_hd U853 ( .A(n2274), .B(n2737), .C(n2785), .D(n2364), .Y(C2_Z_7) );
  ao22d1_hd U854 ( .A(n2274), .B(n2735), .C(n2783), .D(n2364), .Y(C2_Z_8) );
  ao22d1_hd U855 ( .A(n2274), .B(n2733), .C(n2781), .D(n2364), .Y(C2_Z_9) );
  nr2d1_hd U856 ( .A(n2333), .B(n2332), .Y(n2334) );
  ao22d1_hd U857 ( .A(n1891), .B(n2334), .C(n2333), .D(n2362), .Y(
        DP_OP_43J4_124_6938_n32) );
  ao22d1_hd U858 ( .A(b_m[25]), .B(n2362), .C(n2361), .D(n2957), .Y(n2335) );
  oa21d1_hd U859 ( .A(a_m[25]), .B(n2364), .C(n2335), .Y(
        DP_OP_43J4_124_6938_n33) );
  ao22d1_hd U860 ( .A(n2274), .B(n2751), .C(n2361), .D(n2703), .Y(n2336) );
  oa21d1_hd U861 ( .A(n1891), .B(n2703), .C(n2336), .Y(DP_OP_43J4_124_6938_n34) );
  ao22d1_hd U862 ( .A(n2274), .B(n2753), .C(n2361), .D(n2705), .Y(n2337) );
  oa21d1_hd U863 ( .A(n1891), .B(n2705), .C(n2337), .Y(DP_OP_43J4_124_6938_n35) );
  ao22d1_hd U864 ( .A(n2274), .B(n2755), .C(n2361), .D(n2707), .Y(n2338) );
  oa21d1_hd U865 ( .A(n1891), .B(n2707), .C(n2338), .Y(DP_OP_43J4_124_6938_n36) );
  ao22d1_hd U866 ( .A(b_m[21]), .B(n2362), .C(n2361), .D(n2709), .Y(n2339) );
  oa21d1_hd U867 ( .A(a_m[21]), .B(n2364), .C(n2339), .Y(
        DP_OP_43J4_124_6938_n37) );
  ao22d1_hd U868 ( .A(n2274), .B(n2759), .C(n2361), .D(n2711), .Y(n2340) );
  oa21d1_hd U869 ( .A(n1891), .B(n2711), .C(n2340), .Y(DP_OP_43J4_124_6938_n38) );
  ao22d1_hd U870 ( .A(n2274), .B(n2761), .C(n2361), .D(n2713), .Y(n2341) );
  oa21d1_hd U871 ( .A(n1891), .B(n2713), .C(n2341), .Y(DP_OP_43J4_124_6938_n39) );
  ao22d1_hd U872 ( .A(b_m[18]), .B(n2362), .C(n2361), .D(n2715), .Y(n2342) );
  oa21d1_hd U873 ( .A(a_m[18]), .B(n2364), .C(n2342), .Y(
        DP_OP_43J4_124_6938_n40) );
  ao22d1_hd U874 ( .A(b_m[17]), .B(n2362), .C(n2361), .D(n2717), .Y(n2343) );
  oa21d1_hd U875 ( .A(a_m[17]), .B(n2364), .C(n2343), .Y(
        DP_OP_43J4_124_6938_n41) );
  ao22d1_hd U876 ( .A(n2274), .B(n2767), .C(n2361), .D(n2719), .Y(n2344) );
  oa21d1_hd U877 ( .A(n1891), .B(n2719), .C(n2344), .Y(DP_OP_43J4_124_6938_n42) );
  ao22d1_hd U878 ( .A(n2274), .B(n2769), .C(n2361), .D(n2721), .Y(n2345) );
  oa21d1_hd U879 ( .A(n1891), .B(n2721), .C(n2345), .Y(DP_OP_43J4_124_6938_n43) );
  ao22d1_hd U880 ( .A(b_m[14]), .B(n2362), .C(n2361), .D(n2723), .Y(n2346) );
  oa21d1_hd U881 ( .A(a_m[14]), .B(n2364), .C(n2346), .Y(
        DP_OP_43J4_124_6938_n44) );
  ao22d1_hd U882 ( .A(n2274), .B(n2773), .C(n2361), .D(n2725), .Y(n2347) );
  oa21d1_hd U883 ( .A(n1891), .B(n2725), .C(n2347), .Y(DP_OP_43J4_124_6938_n45) );
  ao22d1_hd U884 ( .A(n2274), .B(n2775), .C(b_m[12]), .D(n2362), .Y(n2348) );
  oa21d1_hd U885 ( .A(b_m[12]), .B(n2356), .C(n2348), .Y(
        DP_OP_43J4_124_6938_n46) );
  ao22d1_hd U886 ( .A(n2274), .B(n2777), .C(n2361), .D(n2729), .Y(n2349) );
  oa21d1_hd U887 ( .A(n1891), .B(n2729), .C(n2349), .Y(DP_OP_43J4_124_6938_n47) );
  ao22d1_hd U888 ( .A(n2274), .B(n2779), .C(b_m[10]), .D(n2362), .Y(n2350) );
  oa21d1_hd U889 ( .A(b_m[10]), .B(n2356), .C(n2350), .Y(
        DP_OP_43J4_124_6938_n48) );
  ao22d1_hd U890 ( .A(n2274), .B(n2781), .C(b_m[9]), .D(n2362), .Y(n2351) );
  oa21d1_hd U891 ( .A(b_m[9]), .B(n2356), .C(n2351), .Y(
        DP_OP_43J4_124_6938_n49) );
  ao22d1_hd U892 ( .A(n2274), .B(n2783), .C(n2361), .D(n2735), .Y(n2352) );
  oa21d1_hd U893 ( .A(n1891), .B(n2735), .C(n2352), .Y(DP_OP_43J4_124_6938_n50) );
  ao22d1_hd U894 ( .A(n2274), .B(n2785), .C(n2361), .D(n2737), .Y(n2353) );
  oa21d1_hd U895 ( .A(n1891), .B(n2737), .C(n2353), .Y(DP_OP_43J4_124_6938_n51) );
  ao22d1_hd U896 ( .A(n2274), .B(n2787), .C(b_m[6]), .D(n2362), .Y(n2354) );
  oa21d1_hd U897 ( .A(b_m[6]), .B(n2356), .C(n2354), .Y(
        DP_OP_43J4_124_6938_n52) );
  ao22d1_hd U898 ( .A(n2274), .B(n2789), .C(b_m[5]), .D(n2362), .Y(n2355) );
  oa21d1_hd U899 ( .A(b_m[5]), .B(n2356), .C(n2355), .Y(
        DP_OP_43J4_124_6938_n53) );
  ao22d1_hd U900 ( .A(n2274), .B(n2791), .C(n2361), .D(n2743), .Y(n2357) );
  oa21d1_hd U901 ( .A(n1891), .B(n2743), .C(n2357), .Y(DP_OP_43J4_124_6938_n54) );
  ao22d1_hd U902 ( .A(n2274), .B(n2793), .C(n2361), .D(n2745), .Y(n2358) );
  oa21d1_hd U903 ( .A(n1891), .B(n2745), .C(n2358), .Y(DP_OP_43J4_124_6938_n55) );
  ao22d1_hd U904 ( .A(b_m[2]), .B(n2362), .C(n2361), .D(n2746), .Y(n2359) );
  oa21d1_hd U905 ( .A(a_m[2]), .B(n2364), .C(n2359), .Y(
        DP_OP_43J4_124_6938_n56) );
  ao22d1_hd U906 ( .A(b_m[1]), .B(n2362), .C(n2361), .D(n2748), .Y(n2360) );
  oa21d1_hd U907 ( .A(a_m[1]), .B(n2364), .C(n2360), .Y(
        DP_OP_43J4_124_6938_n57) );
  ao22d1_hd U908 ( .A(b_m[0]), .B(n2362), .C(n2361), .D(n2749), .Y(n2363) );
  oa21d1_hd U909 ( .A(a_m[0]), .B(n2364), .C(n2363), .Y(
        DP_OP_43J4_124_6938_n58) );
  ao22d1_hd U910 ( .A(n2274), .B(n2421), .C(n2437), .D(n2364), .Y(N338) );
  nr4d1_hd U911 ( .A(a_e[6]), .B(a_e[2]), .C(a_e[1]), .D(a_e[5]), .Y(n2365) );
  nd4d1_hd U912 ( .A(a_e[7]), .B(n2365), .C(n2807), .D(n2837), .Y(n2366) );
  nr4d1_hd U913 ( .A(n2810), .B(n2843), .C(n2385), .D(n2366), .Y(n2802) );
  nr4d1_hd U914 ( .A(a_e[8]), .B(a_e[0]), .C(a_e[9]), .D(n2366), .Y(n2496) );
  nr4d1_hd U915 ( .A(b_e[2]), .B(b_e[1]), .C(b_e[3]), .D(b_e[4]), .Y(n2367) );
  nd4d1_hd U916 ( .A(b_e[7]), .B(n2367), .C(n2879), .D(n2891), .Y(n2376) );
  nr4d1_hd U917 ( .A(b_e[9]), .B(b_e[8]), .C(b_e[0]), .D(n2376), .Y(n2495) );
  ivd1_hd U918 ( .A(n2495), .Y(n2418) );
  nd4d1_hd U919 ( .A(n2753), .B(n2779), .C(n2797), .D(n2794), .Y(n2375) );
  nr4d1_hd U920 ( .A(a_m[25]), .B(a_m[11]), .C(a_m[12]), .D(a_m[26]), .Y(n2368) );
  nd4d1_hd U921 ( .A(n2368), .B(n2751), .C(n2759), .D(n2755), .Y(n2374) );
  nr4d1_hd U922 ( .A(a_m[13]), .B(a_m[14]), .C(a_m[15]), .D(a_m[16]), .Y(n2372) );
  nr4d1_hd U923 ( .A(a_m[21]), .B(a_m[17]), .C(a_m[18]), .D(a_m[19]), .Y(n2371) );
  nr4d1_hd U924 ( .A(a_m[5]), .B(a_m[1]), .C(a_m[3]), .D(a_m[4]), .Y(n2370) );
  nr4d1_hd U925 ( .A(a_m[9]), .B(a_m[6]), .C(a_m[7]), .D(a_m[8]), .Y(n2369) );
  nd4d1_hd U926 ( .A(n2372), .B(n2371), .C(n2370), .D(n2369), .Y(n2373) );
  nr3d1_hd U927 ( .A(n2375), .B(n2374), .C(n2373), .Y(n2419) );
  nr4d1_hd U928 ( .A(n2376), .B(n2872), .C(n2405), .D(n2916), .Y(n2868) );
  nd4d1_hd U929 ( .A(n2703), .B(n2717), .C(n2727), .D(n2719), .Y(n2384) );
  nr4d1_hd U930 ( .A(b_m[0]), .B(b_m[7]), .C(b_m[14]), .D(b_m[26]), .Y(n2377)
         );
  nd4d1_hd U931 ( .A(n2377), .B(n2705), .C(n2748), .D(n2746), .Y(n2383) );
  nr4d1_hd U932 ( .A(b_m[21]), .B(b_m[13]), .C(b_m[19]), .D(b_m[20]), .Y(n2381) );
  nr4d1_hd U933 ( .A(b_m[25]), .B(b_m[10]), .C(b_m[18]), .D(b_m[22]), .Y(n2380) );
  nr4d1_hd U934 ( .A(b_m[3]), .B(b_m[4]), .C(b_m[11]), .D(b_m[15]), .Y(n2379)
         );
  nr4d1_hd U935 ( .A(b_m[9]), .B(b_m[6]), .C(b_m[5]), .D(b_m[8]), .Y(n2378) );
  nd4d1_hd U936 ( .A(n2381), .B(n2380), .C(n2379), .D(n2378), .Y(n2382) );
  nr3d1_hd U937 ( .A(n2384), .B(n2383), .C(n2382), .Y(n2417) );
  nr2d1_hd U938 ( .A(a_e[1]), .B(n2917), .Y(n2391) );
  ao22d1_hd U939 ( .A(b_e[4]), .B(n2807), .C(b_e[5]), .D(n2828), .Y(n2386) );
  ao22d1_hd U940 ( .A(b_e[2]), .B(n2852), .C(b_e[3]), .D(n2837), .Y(n2393) );
  nr2d1_hd U941 ( .A(n2872), .B(a_e[8]), .Y(n2406) );
  ivd1_hd U942 ( .A(n2406), .Y(n2389) );
  nr2d1_hd U943 ( .A(n2874), .B(a_e[7]), .Y(n2402) );
  ivd1_hd U944 ( .A(n2402), .Y(n2388) );
  nd4d1_hd U945 ( .A(n2393), .B(n2389), .C(n2388), .D(n2387), .Y(n2390) );
  ivd1_hd U946 ( .A(n2392), .Y(n2401) );
  ao211d1_hd U947 ( .A(b_e[1]), .B(n2803), .C(b_e[0]), .D(n2843), .Y(n2395) );
  oa22d1_hd U948 ( .A(b_e[2]), .B(n2852), .C(b_e[1]), .D(n2803), .Y(n2394) );
  oa21d1_hd U949 ( .A(n2395), .B(n2394), .C(n2393), .Y(n2397) );
  oa211d1_hd U950 ( .A(b_e[4]), .B(n2807), .C(n2397), .D(n2396), .Y(n2400) );
  oa22d1_hd U951 ( .A(b_e[6]), .B(n2808), .C(b_e[5]), .D(n2828), .Y(n2398) );
  ao22d1_hd U952 ( .A(n2401), .B(n2400), .C(n2399), .D(n2398), .Y(n2403) );
  oa22d1_hd U953 ( .A(b_e[8]), .B(n2810), .C(n2403), .D(n2402), .Y(n2404) );
  ao21d1_hd U954 ( .A(a_e[7]), .B(n2874), .C(n2404), .Y(n2407) );
  oa22d1_hd U955 ( .A(n2407), .B(n2406), .C(a_e[9]), .D(n2405), .Y(n2408) );
  oa21d1_hd U956 ( .A(n2802), .B(n2412), .C(n2279), .Y(n1) );
  oa21d1_hd U957 ( .A(n2868), .B(n2412), .C(n2956), .Y(n2) );
  scg4d1_hd U958 ( .A(n1291), .B(round_bit), .C(z_m[0]), .D(n2516), .E(n2653), 
        .F(sum[3]), .G(n2277), .H(sum[2]), .Y(n266) );
  oa22d1_hd U959 ( .A(n2495), .B(n2420), .C(n2421), .D(n2455), .Y(n2414) );
  ao21d1_hd U960 ( .A(n2270), .B(n2414), .C(n2275), .Y(n2438) );
  ao21d1_hd U961 ( .A(n2416), .B(n2415), .C(n2495), .Y(n2422) );
  oa21d1_hd U962 ( .A(n2422), .B(n2421), .C(n2497), .Y(n2424) );
  ao21d1_hd U963 ( .A(n2270), .B(n2423), .C(n2493), .Y(n2964) );
  ao22d1_hd U964 ( .A(n2270), .B(n2424), .C(n2281), .D(z[31]), .Y(n2436) );
  ivd1_hd U965 ( .A(z_m[15]), .Y(n2560) );
  ivd1_hd U966 ( .A(z_m[16]), .Y(n2551) );
  ivd1_hd U967 ( .A(z_m[2]), .Y(n2637) );
  nd4d1_hd U968 ( .A(n2560), .B(n2551), .C(n2637), .D(n2631), .Y(n2425) );
  nr4d1_hd U969 ( .A(z_m[0]), .B(z_m[22]), .C(z_m[1]), .D(n2425), .Y(n2431) );
  ivd1_hd U970 ( .A(z_m[9]), .Y(n2596) );
  ivd1_hd U971 ( .A(z_m[10]), .Y(n2589) );
  nd4d1_hd U972 ( .A(n2619), .B(n2596), .C(n2589), .D(n2595), .Y(n2429) );
  ivd1_hd U973 ( .A(z_m[5]), .Y(n2620) );
  ivd1_hd U974 ( .A(z_m[6]), .Y(n2613) );
  nd4d1_hd U975 ( .A(n2645), .B(n2620), .C(n2613), .D(n2607), .Y(n2428) );
  ivd1_hd U976 ( .A(z_m[21]), .Y(n2676) );
  ivd1_hd U977 ( .A(z_m[20]), .Y(n2532) );
  ivd1_hd U978 ( .A(z_m[18]), .Y(n2538) );
  nd4d1_hd U979 ( .A(n2676), .B(n2544), .C(n2532), .D(n2538), .Y(n2427) );
  ivd1_hd U980 ( .A(z_m[13]), .Y(n2566) );
  ivd1_hd U981 ( .A(z_m[17]), .Y(n2545) );
  nd4d1_hd U982 ( .A(n2583), .B(n2566), .C(n2572), .D(n2545), .Y(n2426) );
  nr4d1_hd U983 ( .A(n2429), .B(n2428), .C(n2427), .D(n2426), .Y(n2430) );
  ivd1_hd U984 ( .A(z_e[9]), .Y(n2696) );
  nr4d1_hd U985 ( .A(z_e[6]), .B(z_e[4]), .C(z_e[3]), .D(z_e[5]), .Y(n2432) );
  nr4d1_hd U986 ( .A(z_m[23]), .B(z_e[0]), .C(n2696), .D(n2507), .Y(n2433) );
  oa211d1_hd U987 ( .A(n2434), .B(n2440), .C(n2493), .D(z_s), .Y(n2435) );
  oa211d1_hd U988 ( .A(n2438), .B(n2437), .C(n2436), .D(n2435), .Y(n361) );
  nr2d1_hd U989 ( .A(z_e[1]), .B(z_e[0]), .Y(n2482) );
  nr2d1_hd U990 ( .A(z_e[3]), .B(n2476), .Y(n2468) );
  ivd1_hd U991 ( .A(z_e[4]), .Y(n2464) );
  nr2d1_hd U992 ( .A(z_e[5]), .B(n2463), .Y(n2454) );
  ivd1_hd U993 ( .A(z_e[6]), .Y(n2450) );
  nr2d1_hd U994 ( .A(z_e[7]), .B(n2449), .Y(n2441) );
  ao211d1_hd U995 ( .A(z_e[7]), .B(n2449), .C(n2492), .D(n2441), .Y(n2445) );
  nd3d1_hd U996 ( .A(n2803), .B(n2917), .C(n2489), .Y(n2483) );
  nd2bd1_hd U997 ( .AN(b_e[2]), .B(n2852), .Y(n2475) );
  nr2d1_hd U998 ( .A(n2483), .B(n2475), .Y(n2474) );
  nd3d1_hd U999 ( .A(n2474), .B(n2837), .C(n2903), .Y(n2469) );
  nd2bd1_hd U1000 ( .AN(b_e[4]), .B(n2807), .Y(n2462) );
  nr2d1_hd U1001 ( .A(n2469), .B(n2462), .Y(n2461) );
  nd3d1_hd U1002 ( .A(n2461), .B(n2828), .C(n2891), .Y(n2456) );
  nr2d1_hd U1003 ( .A(n2456), .B(n2448), .Y(n2447) );
  nr2d1_hd U1004 ( .A(n2447), .B(n2443), .Y(n2442) );
  ao211d1_hd U1005 ( .A(n2447), .B(n2443), .C(n2484), .D(n2442), .Y(n2444) );
  ao211d1_hd U1006 ( .A(n2281), .B(z[30]), .C(n2445), .D(n2444), .Y(n2446) );
  ao21d1_hd U1007 ( .A(n2456), .B(n2448), .C(n2447), .Y(n2453) );
  ivd1_hd U1008 ( .A(n2492), .Y(n2479) );
  oa21d1_hd U1009 ( .A(n2454), .B(n2450), .C(n2449), .Y(n2451) );
  ao22d1_hd U1010 ( .A(n2281), .B(z[29]), .C(n2479), .D(n2451), .Y(n2452) );
  oa211d1_hd U1011 ( .A(n2453), .B(n2484), .C(n2491), .D(n2452), .Y(n363) );
  ao21d1_hd U1012 ( .A(z_e[5]), .B(n2463), .C(n2454), .Y(n2460) );
  nr3d1_hd U1013 ( .A(n2495), .B(n2455), .C(n2930), .Y(n2505) );
  ao22d1_hd U1014 ( .A(a_e[5]), .B(n2500), .C(b_e[5]), .D(n2276), .Y(n2457) );
  oa22d1_hd U1015 ( .A(n2461), .B(n2457), .C(n2484), .D(n2456), .Y(n2458) );
  ao21d1_hd U1016 ( .A(n2281), .B(z[28]), .C(n2458), .Y(n2459) );
  oa211d1_hd U1017 ( .A(n2460), .B(n2492), .C(n2491), .D(n2459), .Y(n364) );
  ao21d1_hd U1018 ( .A(n2469), .B(n2462), .C(n2461), .Y(n2467) );
  oa21d1_hd U1019 ( .A(n2468), .B(n2464), .C(n2463), .Y(n2465) );
  ao22d1_hd U1020 ( .A(n2281), .B(z[27]), .C(n2479), .D(n2465), .Y(n2466) );
  oa211d1_hd U1021 ( .A(n2467), .B(n2484), .C(n2491), .D(n2466), .Y(n365) );
  ao21d1_hd U1022 ( .A(z_e[3]), .B(n2476), .C(n2468), .Y(n2473) );
  ao22d1_hd U1023 ( .A(a_e[3]), .B(n2500), .C(b_e[3]), .D(n2276), .Y(n2470) );
  oa22d1_hd U1024 ( .A(n2474), .B(n2470), .C(n2484), .D(n2469), .Y(n2471) );
  ao21d1_hd U1025 ( .A(n2281), .B(z[26]), .C(n2471), .Y(n2472) );
  oa211d1_hd U1026 ( .A(n2473), .B(n2492), .C(n2491), .D(n2472), .Y(n366) );
  ao21d1_hd U1027 ( .A(n2483), .B(n2475), .C(n2474), .Y(n2481) );
  oa21d1_hd U1028 ( .A(n2482), .B(n2477), .C(n2476), .Y(n2478) );
  ao22d1_hd U1029 ( .A(n2281), .B(z[25]), .C(n2479), .D(n2478), .Y(n2480) );
  oa211d1_hd U1030 ( .A(n2481), .B(n2484), .C(n2491), .D(n2480), .Y(n367) );
  ao21d1_hd U1031 ( .A(z_e[0]), .B(z_e[1]), .C(n2482), .Y(n2488) );
  ao22d1_hd U1032 ( .A(a_e[1]), .B(n2500), .C(b_e[1]), .D(n2276), .Y(n2485) );
  oa22d1_hd U1033 ( .A(n2485), .B(n2489), .C(n2484), .D(n2483), .Y(n2486) );
  ao21d1_hd U1034 ( .A(n2281), .B(z[24]), .C(n2486), .Y(n2487) );
  oa211d1_hd U1035 ( .A(n2488), .B(n2492), .C(n2491), .D(n2487), .Y(n368) );
  ao22d1_hd U1036 ( .A(n2281), .B(z[23]), .C(n2500), .D(n2489), .Y(n2490) );
  oa211d1_hd U1037 ( .A(z_e[0]), .B(n2492), .C(n2491), .D(n2490), .Y(n369) );
  ao22d1_hd U1038 ( .A(b_m[25]), .B(n2276), .C(z_m[22]), .D(n2504), .Y(n2502)
         );
  nd3d1_hd U1039 ( .A(n2496), .B(n2495), .C(n1891), .Y(n2498) );
  ao22d1_hd U1040 ( .A(n2281), .B(z[22]), .C(n2500), .D(n2499), .Y(n2501) );
  scg15d1_hd U1041 ( .A(a_m[25]), .B(n2275), .C(n2502), .D(n2501), .Y(n370) );
  scg4d1_hd U1042 ( .A(b_m[24]), .B(n2276), .C(z_m[21]), .D(n2504), .E(a_m[24]), .F(n2275), .G(n2281), .H(z[21]), .Y(n371) );
  scg4d1_hd U1043 ( .A(b_m[23]), .B(n2276), .C(z_m[20]), .D(n2504), .E(a_m[23]), .F(n2503), .G(n2281), .H(z[20]), .Y(n372) );
  scg4d1_hd U1044 ( .A(b_m[22]), .B(n2276), .C(z_m[19]), .D(n2504), .E(a_m[22]), .F(n2275), .G(n2281), .H(z[19]), .Y(n373) );
  scg4d1_hd U1045 ( .A(b_m[21]), .B(n2276), .C(z_m[18]), .D(n2504), .E(a_m[21]), .F(n2275), .G(n2281), .H(z[18]), .Y(n374) );
  scg4d1_hd U1046 ( .A(b_m[20]), .B(n2276), .C(z_m[17]), .D(n2504), .E(a_m[20]), .F(n2275), .G(n2281), .H(z[17]), .Y(n375) );
  scg4d1_hd U1047 ( .A(b_m[19]), .B(n2276), .C(z_m[16]), .D(n2504), .E(a_m[19]), .F(n2275), .G(n2281), .H(z[16]), .Y(n376) );
  scg4d1_hd U1048 ( .A(b_m[18]), .B(n2276), .C(z_m[15]), .D(n2504), .E(a_m[18]), .F(n2275), .G(n2281), .H(z[15]), .Y(n377) );
  scg4d1_hd U1049 ( .A(a_m[17]), .B(n2275), .C(z_m[14]), .D(n2504), .E(n2276), 
        .F(b_m[17]), .G(n2281), .H(z[14]), .Y(n378) );
  scg4d1_hd U1050 ( .A(b_m[16]), .B(n2276), .C(z_m[13]), .D(n2504), .E(a_m[16]), .F(n2275), .G(n2281), .H(z[13]), .Y(n379) );
  scg4d1_hd U1051 ( .A(b_m[15]), .B(n2276), .C(z_m[12]), .D(n2504), .E(a_m[15]), .F(n2503), .G(n2281), .H(z[12]), .Y(n380) );
  scg4d1_hd U1052 ( .A(b_m[14]), .B(n2276), .C(z_m[11]), .D(n2504), .E(a_m[14]), .F(n2503), .G(n2281), .H(z[11]), .Y(n381) );
  scg4d1_hd U1053 ( .A(b_m[13]), .B(n2276), .C(z_m[10]), .D(n2504), .E(a_m[13]), .F(n2503), .G(n2281), .H(z[10]), .Y(n382) );
  scg4d1_hd U1054 ( .A(b_m[12]), .B(n2276), .C(z_m[9]), .D(n2504), .E(a_m[12]), 
        .F(n2503), .G(n2281), .H(z[9]), .Y(n383) );
  scg4d1_hd U1055 ( .A(b_m[11]), .B(n2276), .C(z_m[8]), .D(n2504), .E(a_m[11]), 
        .F(n2275), .G(n2281), .H(z[8]), .Y(n384) );
  scg4d1_hd U1056 ( .A(b_m[10]), .B(n2276), .C(z_m[7]), .D(n2504), .E(a_m[10]), 
        .F(n2275), .G(n2281), .H(z[7]), .Y(n385) );
  scg4d1_hd U1057 ( .A(b_m[9]), .B(n2276), .C(z_m[6]), .D(n2504), .E(a_m[9]), 
        .F(n2275), .G(n2281), .H(z[6]), .Y(n386) );
  scg4d1_hd U1058 ( .A(b_m[8]), .B(n2276), .C(z_m[5]), .D(n2504), .E(a_m[8]), 
        .F(n2275), .G(n2281), .H(z[5]), .Y(n387) );
  scg4d1_hd U1059 ( .A(b_m[7]), .B(n2276), .C(z_m[4]), .D(n2504), .E(a_m[7]), 
        .F(n2275), .G(n2281), .H(z[4]), .Y(n388) );
  scg4d1_hd U1060 ( .A(b_m[6]), .B(n2276), .C(z_m[3]), .D(n2504), .E(a_m[6]), 
        .F(n2275), .G(n2281), .H(z[3]), .Y(n389) );
  scg4d1_hd U1061 ( .A(b_m[5]), .B(n2276), .C(z_m[2]), .D(n2504), .E(a_m[5]), 
        .F(n2275), .G(n2281), .H(z[2]), .Y(n390) );
  scg4d1_hd U1062 ( .A(b_m[4]), .B(n2276), .C(z_m[1]), .D(n2504), .E(a_m[4]), 
        .F(n2275), .G(n2281), .H(z[1]), .Y(n391) );
  scg4d1_hd U1063 ( .A(b_m[3]), .B(n2276), .C(z_m[0]), .D(n2504), .E(a_m[3]), 
        .F(n2503), .G(n2281), .H(z[0]), .Y(n392) );
  ao22d1_hd U1064 ( .A(n2681), .B(sum[0]), .C(sticky), .D(n2513), .Y(n2510) );
  scg16d1_hd U1065 ( .A(n2507), .B(n2506), .C(z_e[9]), .Y(n2511) );
  nr2d1_hd U1066 ( .A(n2508), .B(n2511), .Y(n2935) );
  ao22d1_hd U1067 ( .A(n2512), .B(round_bit), .C(n2653), .D(sum[1]), .Y(n2509)
         );
  scg21d1_hd U1068 ( .A(n2511), .B(z_e[0]), .C(z_m[23]), .D(n2935), .Y(n2940)
         );
  ao21d1_hd U1069 ( .A(n2940), .B(n1291), .C(n2512), .Y(n2680) );
  ao22d1_hd U1070 ( .A(n2653), .B(sum[2]), .C(n2277), .D(sum[1]), .Y(n2515) );
  nd3d1_hd U1071 ( .A(n2516), .B(guard), .C(n1222), .Y(n2514) );
  oa211d1_hd U1072 ( .A(n2517), .B(n1222), .C(n2515), .D(n2514), .Y(n394) );
  oa211d1_hd U1073 ( .A(sticky), .B(n2518), .C(guard), .D(n2682), .Y(n2519) );
  ao22d1_hd U1074 ( .A(n2653), .B(sum[26]), .C(n2277), .D(sum[25]), .Y(n2523)
         );
  ivd1_hd U1075 ( .A(n2674), .Y(n2520) );
  nd3d1_hd U1076 ( .A(z_m[0]), .B(z_m[1]), .C(z_m[2]), .Y(n2626) );
  nr3d1_hd U1077 ( .A(n2626), .B(n2631), .C(n2645), .Y(n2614) );
  nd3d1_hd U1078 ( .A(n2614), .B(z_m[5]), .C(z_m[6]), .Y(n2602) );
  nr3d1_hd U1079 ( .A(n2602), .B(n2607), .C(n2619), .Y(n2590) );
  nd3d1_hd U1080 ( .A(n2590), .B(z_m[9]), .C(z_m[10]), .Y(n2578) );
  nr3d1_hd U1081 ( .A(n2578), .B(n2595), .C(n2583), .Y(n2567) );
  nd3d1_hd U1082 ( .A(n2567), .B(z_m[13]), .C(z_m[14]), .Y(n2552) );
  nr2d1_hd U1083 ( .A(n2553), .B(n2552), .Y(n2539) );
  nd3d1_hd U1084 ( .A(n2539), .B(z_m[17]), .C(z_m[18]), .Y(n2673) );
  nr2d1_hd U1085 ( .A(n2673), .B(n2639), .Y(n2535) );
  oa21d1_hd U1086 ( .A(z_m[22]), .B(n2668), .C(n2666), .Y(n2521) );
  ao21d1_hd U1087 ( .A(n2673), .B(n2682), .C(n2640), .Y(n2533) );
  oa21d1_hd U1088 ( .A(z_m[21]), .B(n2639), .C(n2524), .Y(n2663) );
  ao22d1_hd U1089 ( .A(z_m[21]), .B(n2521), .C(z_m[22]), .D(n2663), .Y(n2522)
         );
  oa211d1_hd U1090 ( .A(n2675), .B(n2654), .C(n2523), .D(n2522), .Y(n395) );
  ao22d1_hd U1091 ( .A(n2653), .B(sum[25]), .C(n2277), .D(sum[24]), .Y(n2527)
         );
  ao22d1_hd U1092 ( .A(z_m[21]), .B(n2524), .C(n2668), .D(n2676), .Y(n2525) );
  ao21d1_hd U1093 ( .A(n2658), .B(z_m[20]), .C(n2525), .Y(n2526) );
  oa211d1_hd U1094 ( .A(n2664), .B(n2654), .C(n2527), .D(n2526), .Y(n396) );
  ao21d1_hd U1095 ( .A(n2535), .B(n2532), .C(n2658), .Y(n2531) );
  ao22d1_hd U1096 ( .A(n2653), .B(sum[24]), .C(n2277), .D(sum[23]), .Y(n2530)
         );
  oa21d1_hd U1097 ( .A(z_m[19]), .B(n2639), .C(n2533), .Y(n2528) );
  ao22d1_hd U1098 ( .A(z_m[21]), .B(n2647), .C(z_m[20]), .D(n2528), .Y(n2529)
         );
  oa211d1_hd U1099 ( .A(n2531), .B(n2544), .C(n2530), .D(n2529), .Y(n397) );
  ao22d1_hd U1100 ( .A(n2653), .B(sum[23]), .C(n2277), .D(sum[22]), .Y(n2537)
         );
  oa22d1_hd U1101 ( .A(n2533), .B(n2544), .C(n2532), .D(n2654), .Y(n2534) );
  ao21d1_hd U1102 ( .A(n2535), .B(n2544), .C(n2534), .Y(n2536) );
  oa211d1_hd U1103 ( .A(n2666), .B(n2538), .C(n2537), .D(n2536), .Y(n398) );
  ao22d1_hd U1104 ( .A(n2653), .B(sum[22]), .C(n2277), .D(sum[21]), .Y(n2543)
         );
  oa21d1_hd U1105 ( .A(z_m[18]), .B(n2546), .C(n2666), .Y(n2541) );
  scg20d1_hd U1106 ( .A(n2963), .B(n2539), .C(n2640), .Y(n2547) );
  oa21d1_hd U1107 ( .A(z_m[17]), .B(n2639), .C(n2547), .Y(n2540) );
  ao22d1_hd U1108 ( .A(z_m[17]), .B(n2541), .C(z_m[18]), .D(n2540), .Y(n2542)
         );
  oa211d1_hd U1109 ( .A(n2544), .B(n2654), .C(n2543), .D(n2542), .Y(n399) );
  ao22d1_hd U1110 ( .A(n2653), .B(sum[21]), .C(n2277), .D(sum[20]), .Y(n2550)
         );
  ao22d1_hd U1111 ( .A(z_m[17]), .B(n2547), .C(n2546), .D(n2545), .Y(n2548) );
  ao21d1_hd U1112 ( .A(z_m[18]), .B(n2647), .C(n2548), .Y(n2549) );
  oa211d1_hd U1113 ( .A(n2666), .B(n2551), .C(n2550), .D(n2549), .Y(n400) );
  ao22d1_hd U1114 ( .A(n2653), .B(sum[20]), .C(n2277), .D(sum[19]), .Y(n2558)
         );
  ivd1_hd U1115 ( .A(n2552), .Y(n2561) );
  oa21d1_hd U1116 ( .A(n2561), .B(n2963), .C(n2661), .Y(n2559) );
  ao22d1_hd U1117 ( .A(z_m[16]), .B(n2559), .C(z_m[17]), .D(n2647), .Y(n2557)
         );
  nr2d1_hd U1118 ( .A(n2560), .B(n2552), .Y(n2554) );
  oa211d1_hd U1119 ( .A(z_m[16]), .B(n2554), .C(n2665), .D(n2553), .Y(n2556)
         );
  nd4d1_hd U1120 ( .A(n2558), .B(n2557), .C(n2556), .D(n2555), .Y(n401) );
  ao22d1_hd U1121 ( .A(n2653), .B(sum[19]), .C(n2277), .D(sum[18]), .Y(n2565)
         );
  ao22d1_hd U1122 ( .A(z_m[15]), .B(n2559), .C(z_m[16]), .D(n2647), .Y(n2564)
         );
  nd3d1_hd U1123 ( .A(n2561), .B(n2665), .C(n2560), .Y(n2563) );
  nd4d1_hd U1124 ( .A(n2565), .B(n2564), .C(n2563), .D(n2562), .Y(n402) );
  oa21d1_hd U1125 ( .A(n2567), .B(n2963), .C(n2661), .Y(n2575) );
  ao21d1_hd U1126 ( .A(n2665), .B(n2566), .C(n2575), .Y(n2571) );
  ao22d1_hd U1127 ( .A(n2653), .B(sum[18]), .C(n2277), .D(sum[17]), .Y(n2570)
         );
  oa21d1_hd U1128 ( .A(z_m[14]), .B(n2573), .C(n2666), .Y(n2568) );
  ao22d1_hd U1129 ( .A(z_m[15]), .B(n2647), .C(z_m[13]), .D(n2568), .Y(n2569)
         );
  oa211d1_hd U1130 ( .A(n2571), .B(n2572), .C(n2570), .D(n2569), .Y(n403) );
  ao22d1_hd U1131 ( .A(n2653), .B(sum[17]), .C(n2277), .D(sum[16]), .Y(n2577)
         );
  oa22d1_hd U1132 ( .A(z_m[13]), .B(n2573), .C(n2654), .D(n2572), .Y(n2574) );
  ao21d1_hd U1133 ( .A(z_m[13]), .B(n2575), .C(n2574), .Y(n2576) );
  oa211d1_hd U1134 ( .A(n2666), .B(n2583), .C(n2577), .D(n2576), .Y(n404) );
  nr2d1_hd U1135 ( .A(n2578), .B(n2639), .Y(n2586) );
  ao21d1_hd U1136 ( .A(n2586), .B(n2583), .C(n2658), .Y(n2582) );
  ao22d1_hd U1137 ( .A(n2653), .B(sum[16]), .C(n2277), .D(sum[15]), .Y(n2581)
         );
  ao21d1_hd U1138 ( .A(n2682), .B(n2578), .C(n2640), .Y(n2584) );
  oa21d1_hd U1139 ( .A(z_m[11]), .B(n2639), .C(n2584), .Y(n2579) );
  ao22d1_hd U1140 ( .A(z_m[12]), .B(n2579), .C(z_m[13]), .D(n2647), .Y(n2580)
         );
  oa211d1_hd U1141 ( .A(n2582), .B(n2595), .C(n2581), .D(n2580), .Y(n405) );
  ao22d1_hd U1142 ( .A(n2653), .B(sum[15]), .C(n2277), .D(sum[14]), .Y(n2588)
         );
  oa22d1_hd U1143 ( .A(n2584), .B(n2595), .C(n2583), .D(n2654), .Y(n2585) );
  ao21d1_hd U1144 ( .A(n2586), .B(n2595), .C(n2585), .Y(n2587) );
  oa211d1_hd U1145 ( .A(n2666), .B(n2589), .C(n2588), .D(n2587), .Y(n406) );
  ao22d1_hd U1146 ( .A(n2653), .B(sum[14]), .C(n2277), .D(sum[13]), .Y(n2594)
         );
  oa21d1_hd U1147 ( .A(z_m[10]), .B(n2597), .C(n2666), .Y(n2592) );
  scg20d1_hd U1148 ( .A(n2963), .B(n2590), .C(n2640), .Y(n2598) );
  oa21d1_hd U1149 ( .A(z_m[9]), .B(n2639), .C(n2598), .Y(n2591) );
  ao22d1_hd U1150 ( .A(z_m[9]), .B(n2592), .C(z_m[10]), .D(n2591), .Y(n2593)
         );
  oa211d1_hd U1151 ( .A(n2595), .B(n2654), .C(n2594), .D(n2593), .Y(n407) );
  ao22d1_hd U1152 ( .A(n2653), .B(sum[13]), .C(n2277), .D(sum[12]), .Y(n2601)
         );
  ao22d1_hd U1153 ( .A(z_m[9]), .B(n2598), .C(n2597), .D(n2596), .Y(n2599) );
  ao21d1_hd U1154 ( .A(z_m[10]), .B(n2647), .C(n2599), .Y(n2600) );
  oa211d1_hd U1155 ( .A(n2666), .B(n2607), .C(n2601), .D(n2600), .Y(n408) );
  nr2d1_hd U1156 ( .A(n2602), .B(n2639), .Y(n2610) );
  ao21d1_hd U1157 ( .A(n2610), .B(n2607), .C(n2658), .Y(n2606) );
  ao22d1_hd U1158 ( .A(n2653), .B(sum[12]), .C(n2277), .D(sum[11]), .Y(n2605)
         );
  ao21d1_hd U1159 ( .A(n2682), .B(n2602), .C(n2640), .Y(n2608) );
  oa21d1_hd U1160 ( .A(z_m[7]), .B(n2639), .C(n2608), .Y(n2603) );
  ao22d1_hd U1161 ( .A(z_m[8]), .B(n2603), .C(z_m[9]), .D(n2647), .Y(n2604) );
  oa211d1_hd U1162 ( .A(n2606), .B(n2619), .C(n2605), .D(n2604), .Y(n409) );
  ao22d1_hd U1163 ( .A(n2653), .B(sum[11]), .C(n2277), .D(sum[10]), .Y(n2612)
         );
  oa22d1_hd U1164 ( .A(n2608), .B(n2619), .C(n2607), .D(n2654), .Y(n2609) );
  ao21d1_hd U1165 ( .A(n2610), .B(n2619), .C(n2609), .Y(n2611) );
  oa211d1_hd U1166 ( .A(n2666), .B(n2613), .C(n2612), .D(n2611), .Y(n410) );
  ao22d1_hd U1167 ( .A(n2653), .B(sum[10]), .C(n2277), .D(sum[9]), .Y(n2618)
         );
  oa21d1_hd U1168 ( .A(z_m[6]), .B(n2621), .C(n2666), .Y(n2616) );
  scg20d1_hd U1169 ( .A(n2963), .B(n2614), .C(n2640), .Y(n2622) );
  oa21d1_hd U1170 ( .A(z_m[5]), .B(n2639), .C(n2622), .Y(n2615) );
  ao22d1_hd U1171 ( .A(z_m[5]), .B(n2616), .C(z_m[6]), .D(n2615), .Y(n2617) );
  oa211d1_hd U1172 ( .A(n2619), .B(n2654), .C(n2618), .D(n2617), .Y(n411) );
  ao22d1_hd U1173 ( .A(n2653), .B(sum[9]), .C(n2277), .D(sum[8]), .Y(n2625) );
  ao22d1_hd U1174 ( .A(z_m[5]), .B(n2622), .C(n2621), .D(n2620), .Y(n2623) );
  ao21d1_hd U1175 ( .A(z_m[6]), .B(n2647), .C(n2623), .Y(n2624) );
  oa211d1_hd U1176 ( .A(n2666), .B(n2631), .C(n2625), .D(n2624), .Y(n412) );
  nr2d1_hd U1177 ( .A(n2626), .B(n2639), .Y(n2634) );
  ao21d1_hd U1178 ( .A(n2634), .B(n2631), .C(n2658), .Y(n2630) );
  ao22d1_hd U1179 ( .A(n2653), .B(sum[8]), .C(n2277), .D(sum[7]), .Y(n2629) );
  ao21d1_hd U1180 ( .A(n2682), .B(n2626), .C(n2640), .Y(n2632) );
  oa21d1_hd U1181 ( .A(z_m[3]), .B(n2639), .C(n2632), .Y(n2627) );
  ao22d1_hd U1182 ( .A(z_m[4]), .B(n2627), .C(z_m[5]), .D(n2647), .Y(n2628) );
  oa211d1_hd U1183 ( .A(n2630), .B(n2645), .C(n2629), .D(n2628), .Y(n413) );
  ao22d1_hd U1184 ( .A(n2653), .B(sum[7]), .C(n2277), .D(sum[6]), .Y(n2636) );
  oa22d1_hd U1185 ( .A(n2632), .B(n2645), .C(n2631), .D(n2654), .Y(n2633) );
  ao21d1_hd U1186 ( .A(n2634), .B(n2645), .C(n2633), .Y(n2635) );
  oa211d1_hd U1187 ( .A(n2666), .B(n2637), .C(n2636), .D(n2635), .Y(n414) );
  ao22d1_hd U1188 ( .A(n2653), .B(sum[6]), .C(n2277), .D(sum[5]), .Y(n2644) );
  oa21d1_hd U1189 ( .A(z_m[2]), .B(n2638), .C(n2666), .Y(n2642) );
  nr2d1_hd U1190 ( .A(z_m[0]), .B(n2639), .Y(n2657) );
  nr2d1_hd U1191 ( .A(n2640), .B(n2657), .Y(n2651) );
  ao22d1_hd U1192 ( .A(z_m[1]), .B(n2642), .C(z_m[2]), .D(n2641), .Y(n2643) );
  oa211d1_hd U1193 ( .A(n2645), .B(n2654), .C(n2644), .D(n2643), .Y(n415) );
  ao22d1_hd U1194 ( .A(n2653), .B(sum[5]), .C(n2277), .D(sum[4]), .Y(n2650) );
  ao22d1_hd U1195 ( .A(z_m[0]), .B(n2648), .C(z_m[2]), .D(n2647), .Y(n2649) );
  oa211d1_hd U1196 ( .A(n2651), .B(n2655), .C(n2650), .D(n2649), .Y(n416) );
  ao22d1_hd U1197 ( .A(n2653), .B(sum[4]), .C(n2277), .D(sum[3]), .Y(n2660) );
  nr2d1_hd U1198 ( .A(n2655), .B(n2654), .Y(n2656) );
  ao211d1_hd U1199 ( .A(n2658), .B(guard), .C(n2657), .D(n2656), .Y(n2659) );
  oa211d1_hd U1200 ( .A(n2662), .B(n2661), .C(n2660), .D(n2659), .Y(n417) );
  ao21d1_hd U1201 ( .A(n2665), .B(n2664), .C(n2663), .Y(n2671) );
  oa21d1_hd U1202 ( .A(n2668), .B(n2667), .C(n2666), .Y(n2669) );
  ao22d1_hd U1203 ( .A(n2681), .B(sum[26]), .C(z_m[22]), .D(n2669), .Y(n2670)
         );
  oa211d1_hd U1204 ( .A(n2671), .B(n2675), .C(n2670), .D(n2679), .Y(n418) );
  nr4d1_hd U1205 ( .A(n2676), .B(n2675), .C(n2674), .D(n2673), .Y(n2677) );
  nd4d1_hd U1206 ( .A(n2682), .B(guard), .C(z_m[22]), .D(n2677), .Y(n2678) );
  nd4d1_hd U1207 ( .A(n2680), .B(n1284), .C(n2679), .D(n2678), .Y(n2693) );
  nr3d1_hd U1208 ( .A(n2682), .B(state[1]), .C(n2681), .Y(n2683) );
  ao22d1_hd U1209 ( .A(a_e[8]), .B(n2273), .C(n2698), .D(C91_DATA2_8), .Y(
        n2684) );
  scg14d1_hd U1210 ( .A(z_e[8]), .B(n2695), .C(n2684), .Y(n419) );
  ao22d1_hd U1211 ( .A(z_e[7]), .B(n2695), .C(n2698), .D(C91_DATA2_7), .Y(
        n2685) );
  oa21d1_hd U1212 ( .A(n2812), .B(n1284), .C(n2685), .Y(n420) );
  ao22d1_hd U1213 ( .A(z_e[6]), .B(n2695), .C(n2698), .D(C91_DATA2_6), .Y(
        n2686) );
  oa21d1_hd U1214 ( .A(n2808), .B(n1284), .C(n2686), .Y(n421) );
  ao22d1_hd U1215 ( .A(z_e[5]), .B(n2695), .C(n2698), .D(C91_DATA2_5), .Y(
        n2687) );
  oa21d1_hd U1216 ( .A(n2828), .B(n1284), .C(n2687), .Y(n422) );
  ao22d1_hd U1217 ( .A(z_e[4]), .B(n2695), .C(n2698), .D(C91_DATA2_4), .Y(
        n2688) );
  oa21d1_hd U1218 ( .A(n2807), .B(n1284), .C(n2688), .Y(n423) );
  ao22d1_hd U1219 ( .A(z_e[3]), .B(n2695), .C(n2698), .D(C91_DATA2_3), .Y(
        n2689) );
  oa21d1_hd U1220 ( .A(n2837), .B(n1284), .C(n2689), .Y(n424) );
  ao22d1_hd U1221 ( .A(z_e[2]), .B(n2695), .C(n2698), .D(C91_DATA2_2), .Y(
        n2690) );
  oa21d1_hd U1222 ( .A(n2852), .B(n1284), .C(n2690), .Y(n425) );
  ao22d1_hd U1223 ( .A(z_e[1]), .B(n2695), .C(n2698), .D(C91_DATA2_1), .Y(
        n2691) );
  oa21d1_hd U1224 ( .A(n2803), .B(n1284), .C(n2691), .Y(n426) );
  ao22d1_hd U1225 ( .A(a_e[0]), .B(n2273), .C(n2698), .D(n2694), .Y(n2692) );
  oa21d1_hd U1226 ( .A(n2694), .B(n2693), .C(n2692), .Y(n427) );
  ao22d1_hd U1227 ( .A(a_e[9]), .B(n2273), .C(z_e[9]), .D(n2695), .Y(n2701) );
  ao22d1_hd U1228 ( .A(n1291), .B(z_e[9]), .C(n2696), .D(n2939), .Y(n2699) );
  oa211d1_hd U1229 ( .A(DP_OP_154J4_137_6175_n2), .B(n2699), .C(n2698), .D(
        n2697), .Y(n2700) );
  ao22d1_hd U1230 ( .A(b_m[25]), .B(n2954), .C(n2282), .D(b[21]), .Y(n2702) );
  oa21d1_hd U1231 ( .A(n2703), .B(n2280), .C(n2702), .Y(n429) );
  ao22d1_hd U1232 ( .A(b_m[24]), .B(n2954), .C(n2283), .D(b[20]), .Y(n2704) );
  oa21d1_hd U1233 ( .A(n2705), .B(n2280), .C(n2704), .Y(n430) );
  ao22d1_hd U1234 ( .A(b_m[23]), .B(n2954), .C(n2284), .D(b[19]), .Y(n2706) );
  oa21d1_hd U1235 ( .A(n2707), .B(n2280), .C(n2706), .Y(n431) );
  ao22d1_hd U1236 ( .A(b_m[22]), .B(n2954), .C(n2283), .D(b[18]), .Y(n2708) );
  oa21d1_hd U1237 ( .A(n2709), .B(n2280), .C(n2708), .Y(n432) );
  ao22d1_hd U1238 ( .A(b_m[21]), .B(n2954), .C(n2284), .D(b[17]), .Y(n2710) );
  oa21d1_hd U1239 ( .A(n2711), .B(n2280), .C(n2710), .Y(n433) );
  ao22d1_hd U1240 ( .A(b_m[20]), .B(n2954), .C(n2283), .D(b[16]), .Y(n2712) );
  oa21d1_hd U1241 ( .A(n2713), .B(n2280), .C(n2712), .Y(n434) );
  ao22d1_hd U1242 ( .A(b_m[19]), .B(n2954), .C(n2284), .D(b[15]), .Y(n2714) );
  oa21d1_hd U1243 ( .A(n2715), .B(n2280), .C(n2714), .Y(n435) );
  ao22d1_hd U1244 ( .A(b_m[18]), .B(n2954), .C(n2284), .D(b[14]), .Y(n2716) );
  oa21d1_hd U1245 ( .A(n2717), .B(n2280), .C(n2716), .Y(n436) );
  ao22d1_hd U1246 ( .A(b_m[17]), .B(n2954), .C(n2283), .D(b[13]), .Y(n2718) );
  oa21d1_hd U1247 ( .A(n2719), .B(n2280), .C(n2718), .Y(n437) );
  ao22d1_hd U1248 ( .A(b_m[16]), .B(n2954), .C(n2284), .D(b[12]), .Y(n2720) );
  oa21d1_hd U1249 ( .A(n2721), .B(n2280), .C(n2720), .Y(n438) );
  ao22d1_hd U1250 ( .A(b_m[15]), .B(n2954), .C(n2283), .D(b[11]), .Y(n2722) );
  oa21d1_hd U1251 ( .A(n2723), .B(n2280), .C(n2722), .Y(n439) );
  ao22d1_hd U1252 ( .A(b_m[14]), .B(n2954), .C(n2284), .D(b[10]), .Y(n2724) );
  oa21d1_hd U1253 ( .A(n2725), .B(n2280), .C(n2724), .Y(n440) );
  ao22d1_hd U1254 ( .A(b_m[13]), .B(n2954), .C(n2283), .D(b[9]), .Y(n2726) );
  oa21d1_hd U1255 ( .A(n2727), .B(n2280), .C(n2726), .Y(n441) );
  ao22d1_hd U1256 ( .A(b_m[12]), .B(n2954), .C(n2283), .D(b[8]), .Y(n2728) );
  oa21d1_hd U1257 ( .A(n2729), .B(n2280), .C(n2728), .Y(n442) );
  ao22d1_hd U1258 ( .A(b_m[11]), .B(n2954), .C(n2283), .D(b[7]), .Y(n2730) );
  oa21d1_hd U1259 ( .A(n2731), .B(n2280), .C(n2730), .Y(n443) );
  ao22d1_hd U1260 ( .A(b_m[10]), .B(n2954), .C(n2283), .D(b[6]), .Y(n2732) );
  oa21d1_hd U1261 ( .A(n2733), .B(n2280), .C(n2732), .Y(n444) );
  ao22d1_hd U1262 ( .A(b_m[9]), .B(n2954), .C(n2283), .D(b[5]), .Y(n2734) );
  oa21d1_hd U1263 ( .A(n2735), .B(n2280), .C(n2734), .Y(n445) );
  ao22d1_hd U1264 ( .A(b_m[8]), .B(n2954), .C(n2283), .D(b[4]), .Y(n2736) );
  oa21d1_hd U1265 ( .A(n2737), .B(n2280), .C(n2736), .Y(n446) );
  ao22d1_hd U1266 ( .A(b_m[7]), .B(n2954), .C(n2283), .D(b[3]), .Y(n2738) );
  oa21d1_hd U1267 ( .A(n2739), .B(n2280), .C(n2738), .Y(n447) );
  ao22d1_hd U1268 ( .A(b_m[6]), .B(n2954), .C(n2283), .D(b[2]), .Y(n2740) );
  oa21d1_hd U1269 ( .A(n2741), .B(n2280), .C(n2740), .Y(n448) );
  ao22d1_hd U1270 ( .A(b_m[5]), .B(n2954), .C(n2283), .D(b[1]), .Y(n2742) );
  oa21d1_hd U1271 ( .A(n2743), .B(n2280), .C(n2742), .Y(n449) );
  ao22d1_hd U1272 ( .A(b_m[4]), .B(n2954), .C(n2283), .D(b[0]), .Y(n2744) );
  oa21d1_hd U1273 ( .A(n2745), .B(n2280), .C(n2744), .Y(n450) );
  oa22d1_hd U1274 ( .A(n2746), .B(n2280), .C(n2745), .D(n2747), .Y(n451) );
  oa22d1_hd U1275 ( .A(n2748), .B(n2280), .C(n2746), .D(n2747), .Y(n452) );
  oa22d1_hd U1276 ( .A(n2284), .B(n2749), .C(n2748), .D(n2747), .Y(n453) );
  ao22d1_hd U1277 ( .A(a_m[25]), .B(n2798), .C(n2283), .D(a[21]), .Y(n2750) );
  oa21d1_hd U1278 ( .A(n2751), .B(n2278), .C(n2750), .Y(n454) );
  ao22d1_hd U1279 ( .A(a_m[24]), .B(n2798), .C(n2283), .D(a[20]), .Y(n2752) );
  oa21d1_hd U1280 ( .A(n2753), .B(n2278), .C(n2752), .Y(n455) );
  ao22d1_hd U1281 ( .A(a_m[23]), .B(n2798), .C(n2283), .D(a[19]), .Y(n2754) );
  oa21d1_hd U1282 ( .A(n2755), .B(n2278), .C(n2754), .Y(n456) );
  ao22d1_hd U1283 ( .A(a_m[22]), .B(n2798), .C(n2283), .D(a[18]), .Y(n2756) );
  oa21d1_hd U1284 ( .A(n2757), .B(n2278), .C(n2756), .Y(n457) );
  ao22d1_hd U1285 ( .A(a_m[21]), .B(n2798), .C(n2283), .D(a[17]), .Y(n2758) );
  oa21d1_hd U1286 ( .A(n2759), .B(n2278), .C(n2758), .Y(n458) );
  ao22d1_hd U1287 ( .A(a_m[20]), .B(n2798), .C(n2283), .D(a[16]), .Y(n2760) );
  oa21d1_hd U1288 ( .A(n2761), .B(n2278), .C(n2760), .Y(n459) );
  ao22d1_hd U1289 ( .A(a_m[19]), .B(n2798), .C(n2283), .D(a[15]), .Y(n2762) );
  oa21d1_hd U1290 ( .A(n2763), .B(n2278), .C(n2762), .Y(n460) );
  ao22d1_hd U1291 ( .A(a_m[18]), .B(n2798), .C(n2283), .D(a[14]), .Y(n2764) );
  oa21d1_hd U1292 ( .A(n2765), .B(n2278), .C(n2764), .Y(n461) );
  ao22d1_hd U1293 ( .A(a_m[17]), .B(n2798), .C(n2283), .D(a[13]), .Y(n2766) );
  oa21d1_hd U1294 ( .A(n2767), .B(n2278), .C(n2766), .Y(n462) );
  ao22d1_hd U1295 ( .A(a_m[16]), .B(n2798), .C(n2283), .D(a[12]), .Y(n2768) );
  oa21d1_hd U1296 ( .A(n2769), .B(n2278), .C(n2768), .Y(n463) );
  ao22d1_hd U1297 ( .A(a_m[15]), .B(n2798), .C(n2283), .D(a[11]), .Y(n2770) );
  oa21d1_hd U1298 ( .A(n2771), .B(n2278), .C(n2770), .Y(n464) );
  ao22d1_hd U1299 ( .A(a_m[14]), .B(n2798), .C(n2282), .D(a[10]), .Y(n2772) );
  oa21d1_hd U1300 ( .A(n2773), .B(n2278), .C(n2772), .Y(n465) );
  ao22d1_hd U1301 ( .A(a_m[13]), .B(n2798), .C(n2282), .D(a[9]), .Y(n2774) );
  oa21d1_hd U1302 ( .A(n2775), .B(n2278), .C(n2774), .Y(n466) );
  ao22d1_hd U1303 ( .A(a_m[12]), .B(n2798), .C(n2282), .D(a[8]), .Y(n2776) );
  oa21d1_hd U1304 ( .A(n2777), .B(n2278), .C(n2776), .Y(n467) );
  ao22d1_hd U1305 ( .A(a_m[11]), .B(n2798), .C(n2282), .D(a[7]), .Y(n2778) );
  oa21d1_hd U1306 ( .A(n2779), .B(n2278), .C(n2778), .Y(n468) );
  ao22d1_hd U1307 ( .A(a_m[10]), .B(n2798), .C(n2282), .D(a[6]), .Y(n2780) );
  oa21d1_hd U1308 ( .A(n2781), .B(n2278), .C(n2780), .Y(n469) );
  ao22d1_hd U1309 ( .A(a_m[9]), .B(n2798), .C(n2282), .D(a[5]), .Y(n2782) );
  oa21d1_hd U1310 ( .A(n2783), .B(n2278), .C(n2782), .Y(n470) );
  ao22d1_hd U1311 ( .A(a_m[8]), .B(n2798), .C(n2282), .D(a[4]), .Y(n2784) );
  oa21d1_hd U1312 ( .A(n2785), .B(n2278), .C(n2784), .Y(n471) );
  ao22d1_hd U1313 ( .A(a_m[7]), .B(n2798), .C(n2282), .D(a[3]), .Y(n2786) );
  oa21d1_hd U1314 ( .A(n2787), .B(n2801), .C(n2786), .Y(n472) );
  ao22d1_hd U1315 ( .A(a_m[6]), .B(n2798), .C(n2283), .D(a[2]), .Y(n2788) );
  oa21d1_hd U1316 ( .A(n2789), .B(n2801), .C(n2788), .Y(n473) );
  ao22d1_hd U1317 ( .A(a_m[5]), .B(n2798), .C(n2282), .D(a[1]), .Y(n2790) );
  oa21d1_hd U1318 ( .A(n2791), .B(n2801), .C(n2790), .Y(n474) );
  ao22d1_hd U1319 ( .A(a_m[4]), .B(n2798), .C(n2282), .D(a[0]), .Y(n2792) );
  oa21d1_hd U1320 ( .A(n2793), .B(n2801), .C(n2792), .Y(n475) );
  oa22d1_hd U1321 ( .A(n2794), .B(n2278), .C(n2793), .D(n2795), .Y(n476) );
  oa22d1_hd U1322 ( .A(n2796), .B(n2278), .C(n2794), .D(n2795), .Y(n477) );
  oa22d1_hd U1323 ( .A(n2284), .B(n2797), .C(n2796), .D(n2795), .Y(n478) );
  ao22d1_hd U1324 ( .A(a_m[26]), .B(n2798), .C(n2282), .D(a[22]), .Y(n2799) );
  oa21d1_hd U1325 ( .A(n2800), .B(n2801), .C(n2799), .Y(n479) );
  nr2d1_hd U1326 ( .A(n2843), .B(n2803), .Y(n2846) );
  ao21d1_hd U1327 ( .A(n2806), .B(n2894), .C(n2860), .Y(n2830) );
  ivd1_hd U1328 ( .A(n2830), .Y(n2839) );
  ao21d1_hd U1329 ( .A(n2894), .B(n2804), .C(n2839), .Y(n2829) );
  oa21d1_hd U1330 ( .A(n2808), .B(n2828), .C(n2894), .Y(n2805) );
  ao21d1_hd U1331 ( .A(n2845), .B(n2812), .C(n2814), .Y(n2863) );
  ivd1_hd U1332 ( .A(a[25]), .Y(n2848) );
  nr2d1_hd U1333 ( .A(n2856), .B(n2848), .Y(n2847) );
  ivd1_hd U1334 ( .A(a[27]), .Y(n2832) );
  nr2d1_hd U1335 ( .A(n2840), .B(n2832), .Y(n2831) );
  ivd1_hd U1336 ( .A(a[29]), .Y(n2818) );
  nr2d1_hd U1337 ( .A(n2825), .B(n2818), .Y(n2811) );
  nr2d1_hd U1338 ( .A(n2811), .B(n2285), .Y(n2821) );
  nr2d1_hd U1339 ( .A(n2864), .B(n2806), .Y(n2838) );
  nr2d1_hd U1340 ( .A(n2807), .B(n2836), .Y(n2824) );
  nr2d1_hd U1341 ( .A(n2808), .B(n2823), .Y(n2813) );
  nd3d1_hd U1342 ( .A(a_e[7]), .B(n2813), .C(n2810), .Y(n2809) );
  oa211d1_hd U1343 ( .A(n2863), .B(n2810), .C(n2865), .D(n2809), .Y(n480) );
  ao22d1_hd U1344 ( .A(a_e[7]), .B(n2814), .C(n2813), .D(n2812), .Y(n2815) );
  oa211d1_hd U1345 ( .A(n2817), .B(n2816), .C(n2815), .D(n2865), .Y(n481) );
  oa21d1_hd U1346 ( .A(a_e[5]), .B(n2864), .C(n2829), .Y(n2819) );
  ao22d1_hd U1347 ( .A(n2821), .B(n2820), .C(a_e[6]), .D(n2819), .Y(n2822) );
  oa211d1_hd U1348 ( .A(a_e[6]), .B(n2823), .C(n2822), .D(n2858), .Y(n482) );
  ao21d1_hd U1349 ( .A(n2824), .B(n2828), .C(n2866), .Y(n2827) );
  oa211d1_hd U1350 ( .A(n2831), .B(a[28]), .C(n2284), .D(n2825), .Y(n2826) );
  oa211d1_hd U1351 ( .A(n2829), .B(n2828), .C(n2827), .D(n2826), .Y(n483) );
  oa21d1_hd U1352 ( .A(a_e[3]), .B(n2864), .C(n2830), .Y(n2834) );
  ao211d1_hd U1353 ( .A(n2840), .B(n2832), .C(n2831), .D(n2285), .Y(n2833) );
  ao211d1_hd U1354 ( .A(a_e[4]), .B(n2834), .C(n2866), .D(n2833), .Y(n2835) );
  oa21d1_hd U1355 ( .A(a_e[4]), .B(n2836), .C(n2835), .Y(n484) );
  ao22d1_hd U1356 ( .A(a_e[3]), .B(n2839), .C(n2838), .D(n2837), .Y(n2842) );
  oa211d1_hd U1357 ( .A(n2847), .B(a[26]), .C(n2284), .D(n2840), .Y(n2841) );
  nd3d1_hd U1358 ( .A(n2842), .B(n2858), .C(n2841), .Y(n485) );
  nr2d1_hd U1359 ( .A(a_e[1]), .B(n2864), .Y(n2855) );
  nr2d1_hd U1360 ( .A(n2855), .B(n2854), .Y(n2853) );
  ao211d1_hd U1361 ( .A(n2856), .B(n2848), .C(n2847), .D(n2285), .Y(n2849) );
  nr2d1_hd U1362 ( .A(n2850), .B(n2849), .Y(n2851) );
  oa211d1_hd U1363 ( .A(n2853), .B(n2852), .C(n2851), .D(n2858), .Y(n486) );
  ao22d1_hd U1364 ( .A(a_e[0]), .B(n2855), .C(a_e[1]), .D(n2854), .Y(n2859) );
  oa211d1_hd U1365 ( .A(a[23]), .B(a[24]), .C(n2284), .D(n2856), .Y(n2857) );
  nd3d1_hd U1366 ( .A(n2859), .B(n2858), .C(n2857), .Y(n487) );
  oa211d1_hd U1367 ( .A(a[23]), .B(n2285), .C(n2862), .D(n2861), .Y(n488) );
  oa21d1_hd U1368 ( .A(a_e[8]), .B(n2864), .C(n2863), .Y(n2867) );
  scg17d1_hd U1369 ( .A(a_e[9]), .B(n2867), .C(n2866), .D(n2865), .Y(n489) );
  nr2d1_hd U1370 ( .A(n2917), .B(n2916), .Y(n2913) );
  nr2d1_hd U1371 ( .A(n2903), .B(n2902), .Y(n2893) );
  ao21d1_hd U1372 ( .A(n2894), .B(n2869), .C(n2924), .Y(n2892) );
  scg14d1_hd U1373 ( .A(n2870), .B(n2894), .C(n2892), .Y(n2876) );
  ao21d1_hd U1374 ( .A(n2914), .B(n2874), .C(n2876), .Y(n2958) );
  ivd1_hd U1375 ( .A(b[25]), .Y(n2909) );
  nr2d1_hd U1376 ( .A(n2919), .B(n2909), .Y(n2908) );
  ivd1_hd U1377 ( .A(b[27]), .Y(n2896) );
  nr2d1_hd U1378 ( .A(n2905), .B(n2896), .Y(n2895) );
  ivd1_hd U1379 ( .A(b[29]), .Y(n2880) );
  nr2d1_hd U1380 ( .A(n2888), .B(n2880), .Y(n2873) );
  nr2d1_hd U1381 ( .A(n2873), .B(n2285), .Y(n2882) );
  nr2d1_hd U1382 ( .A(n2959), .B(n2869), .Y(n2887) );
  ivd1_hd U1383 ( .A(n2887), .Y(n2886) );
  nr2d1_hd U1384 ( .A(n2870), .B(n2886), .Y(n2875) );
  nd3d1_hd U1385 ( .A(b_e[7]), .B(n2875), .C(n2872), .Y(n2871) );
  oa211d1_hd U1386 ( .A(n2958), .B(n2872), .C(n2960), .D(n2871), .Y(n490) );
  ao22d1_hd U1387 ( .A(b_e[7]), .B(n2876), .C(n2875), .D(n2874), .Y(n2877) );
  oa211d1_hd U1388 ( .A(n2285), .B(n2878), .C(n2877), .D(n2960), .Y(n491) );
  oa21d1_hd U1389 ( .A(b_e[5]), .B(n2959), .C(n2892), .Y(n2883) );
  ao22d1_hd U1390 ( .A(b_e[6]), .B(n2883), .C(n2882), .D(n2881), .Y(n2884) );
  oa211d1_hd U1391 ( .A(n2886), .B(n2885), .C(n2884), .D(n2961), .Y(n492) );
  ao21d1_hd U1392 ( .A(n2887), .B(n2891), .C(n2921), .Y(n2890) );
  oa211d1_hd U1393 ( .A(n2895), .B(b[28]), .C(n2284), .D(n2888), .Y(n2889) );
  oa211d1_hd U1394 ( .A(n2892), .B(n2891), .C(n2890), .D(n2889), .Y(n493) );
  ao21d1_hd U1395 ( .A(n2894), .B(n2902), .C(n2924), .Y(n2904) );
  ao211d1_hd U1396 ( .A(n2905), .B(n2896), .C(n2895), .D(n2285), .Y(n2897) );
  ao21d1_hd U1397 ( .A(n2898), .B(b_e[4]), .C(n2897), .Y(n2899) );
  oa211d1_hd U1398 ( .A(b_e[4]), .B(n2900), .C(n2899), .D(n2961), .Y(n494) );
  oa22d1_hd U1399 ( .A(n2904), .B(n2903), .C(n2902), .D(n2901), .Y(n2907) );
  oa211d1_hd U1400 ( .A(n2908), .B(b[26]), .C(n2284), .D(n2905), .Y(n2906) );
  scg13d1_hd U1401 ( .A(n2907), .B(n2921), .C(n2906), .Y(n495) );
  nr2d1_hd U1402 ( .A(b_e[0]), .B(n2959), .Y(n2923) );
  nr2d1_hd U1403 ( .A(n2924), .B(n2923), .Y(n2918) );
  ao211d1_hd U1404 ( .A(n2919), .B(n2909), .C(n2908), .D(n2285), .Y(n2910) );
  ao211d1_hd U1405 ( .A(b_e[2]), .B(n2911), .C(n2921), .D(n2910), .Y(n2912) );
  scg22d1_hd U1406 ( .A(n2914), .B(n2913), .C(b_e[2]), .D(n2912), .Y(n496) );
  oa22d1_hd U1407 ( .A(n2918), .B(n2917), .C(n2916), .D(n2915), .Y(n2922) );
  oa211d1_hd U1408 ( .A(b[23]), .B(b[24]), .C(n2284), .D(n2919), .Y(n2920) );
  scg13d1_hd U1409 ( .A(n2922), .B(n2921), .C(n2920), .Y(n497) );
  ao21d1_hd U1410 ( .A(n2924), .B(b_e[0]), .C(n2923), .Y(n2925) );
  oa21d1_hd U1411 ( .A(b[23]), .B(n2285), .C(n2925), .Y(n498) );
  scg21d1_hd U1412 ( .A(n2926), .B(o_AB_ACK), .C(i_RST), .D(n27), .Y(n499) );
  oa211d1_hd U1413 ( .A(state[3]), .B(n2931), .C(n2930), .D(n2929), .Y(n2946)
         );
  nd3d1_hd U1414 ( .A(n2286), .B(o_Z_STB), .C(i_Z_ACK), .Y(n2970) );
  nd4d1_hd U1415 ( .A(N41), .B(n2963), .C(n2970), .D(n1284), .Y(n2937) );
  ivd1_hd U1416 ( .A(n2932), .Y(n2934) );
  oa22d1_hd U1417 ( .A(n2935), .B(n2965), .C(n2934), .D(n2933), .Y(n2936) );
  nr4d1_hd U1418 ( .A(n27), .B(n2946), .C(n2937), .D(n2936), .Y(n2938) );
  ivd1_hd U1419 ( .A(n2966), .Y(n2943) );
  nr2d1_hd U1420 ( .A(n2941), .B(n2949), .Y(n2942) );
  ao22d1_hd U1421 ( .A(state[2]), .B(n2943), .C(N41), .D(n2942), .Y(n2944) );
  oa21d1_hd U1422 ( .A(n2945), .B(n2968), .C(n2944), .Y(n500) );
  nr2d1_hd U1423 ( .A(n1291), .B(n2946), .Y(n2948) );
  oa22d1_hd U1424 ( .A(n2948), .B(n2968), .C(n2947), .D(n2966), .Y(n501) );
  ao21d1_hd U1425 ( .A(state[1]), .B(n2949), .C(state[0]), .Y(n2950) );
  nr2d1_hd U1426 ( .A(n2951), .B(n2950), .Y(n2953) );
  oa22d1_hd U1427 ( .A(n2953), .B(n2968), .C(n2952), .D(n2966), .Y(n502) );
  ao22d1_hd U1428 ( .A(b_m[26]), .B(n2954), .C(n2282), .D(b[22]), .Y(n2955) );
  oa21d1_hd U1429 ( .A(n2957), .B(n2280), .C(n2955), .Y(n503) );
  oa21d1_hd U1430 ( .A(b_e[8]), .B(n2959), .C(n2958), .Y(n2962) );
  scg15d1_hd U1431 ( .A(b_e[9]), .B(n2962), .C(n2961), .D(n2960), .Y(n504) );
  oa22d1_hd U1432 ( .A(n2969), .B(n2968), .C(n2967), .D(n2966), .Y(n505) );
  ivd1_hd U1433 ( .A(n2970), .Y(n2971) );
  scg21d1_hd U1434 ( .A(n2286), .B(o_Z_STB), .C(i_RST), .D(n2971), .Y(n506) );
endmodule


module iir_notch ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   w_add_1_AB_ACK, w_add_2_AB_ACK, w_add_1_Z_STB, w_add_2_Z_STB,
         r_add_1_AB_STB, r_add_1_Z_ACK, r_add_2_AB_STB, r_add_2_Z_ACK,
         w_mult_1_Z_STB, w_mult_2_Z_STB, w_mult_3_Z_STB, w_mult_1_AB_ACK,
         w_mult_2_AB_ACK, w_mult_3_AB_ACK, r_mult_1_AB_STB, r_mult_1_Z_ACK,
         n_2_net_, r_mult_2_AB_STB, r_mult_2_Z_ACK, n_3_net_, r_mult_3_AB_STB,
         r_mult_3_Z_ACK, n_4_net_, N23, r_pstate_0_, r_counter_1_, N1343,
         N1383, N1402, N1403, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n548, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n791, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n908, n1083, n1086, n1260, n1261, n1262,
         n1266, n1267, n1268, n1269, n1274, n1275, n1281, n1285, n1287, n1289,
         n1291, n1293, n1295, n1297, n1299, n1301, n1303, n1305, n1307, n1309,
         n1311, n1313, n1315, n1317, n1319, n1321, n1323, n1325, n1327, n1329,
         n1331, n1333, n1335, n1337, n1339, n1340, n1341, n1343, n1345, n1347,
         n1351, n1352, n1353, n1358, n1359, n1360, n1361, n1362, n1368, n1369,
         n1370, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1391, n1392, n1393,
         n1394, n1395, n1396, n1399, n1401, n1403, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1477, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n790, n792,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954;
  wire   [31:0] r_add_1_A;
  wire   [31:0] r_add_1_B;
  wire   [31:0] w_add_1_Z;
  wire   [31:0] r_add_2_A;
  wire   [31:0] r_add_2_B;
  wire   [31:0] w_add_2_Z;
  wire   [31:0] r_mult_1_A;
  wire   [31:0] r_mult_1_B;
  wire   [31:0] w_mult_1_Z;
  wire   [31:0] r_mult_2_A;
  wire   [31:0] r_mult_2_B;
  wire   [31:0] w_mult_2_Z;
  wire   [31:0] r_mult_3_A;
  wire   [31:0] r_mult_3_B;
  wire   [31:0] w_mult_3_Z;
  wire   [159:0] r_x_data;
  wire   [127:0] r_y_data;

  float_adder_1 add_1 ( .i_A(r_add_1_A), .i_B(r_add_1_B), .i_AB_STB(
        r_add_1_AB_STB), .o_AB_ACK(w_add_1_AB_ACK), .o_Z(w_add_1_Z), .o_Z_STB(
        w_add_1_Z_STB), .i_Z_ACK(r_add_1_Z_ACK), .i_CLK(i_CLK), .i_RST(N23) );
  float_adder_0 add_2 ( .i_A(r_add_2_A), .i_B(r_add_2_B), .i_AB_STB(
        r_add_2_AB_STB), .o_AB_ACK(w_add_2_AB_ACK), .o_Z(w_add_2_Z), .o_Z_STB(
        w_add_2_Z_STB), .i_Z_ACK(r_add_2_Z_ACK), .i_CLK(i_CLK), .i_RST(N23) );
  float_multiplier mult_1 ( .i_A(r_mult_1_A), .i_B(r_mult_1_B), .i_AB_STB(
        r_mult_1_AB_STB), .o_AB_ACK(w_mult_1_AB_ACK), .o_Z(w_mult_1_Z), 
        .o_Z_STB(w_mult_1_Z_STB), .i_Z_ACK(r_mult_1_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(n_2_net_) );
  float_multiplier mult_2 ( .i_A(r_mult_2_A), .i_B(r_mult_2_B), .i_AB_STB(
        r_mult_2_AB_STB), .o_AB_ACK(w_mult_2_AB_ACK), .o_Z(w_mult_2_Z), 
        .o_Z_STB(w_mult_2_Z_STB), .i_Z_ACK(r_mult_2_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(n_3_net_) );
  float_multiplier mult_3 ( .i_A(r_mult_3_A), .i_B(r_mult_3_B), .i_AB_STB(
        r_mult_3_AB_STB), .o_AB_ACK(w_mult_3_AB_ACK), .o_Z(w_mult_3_Z), 
        .o_Z_STB(w_mult_3_Z_STB), .i_Z_ACK(r_mult_3_Z_ACK), .i_CLK(i_CLK), 
        .i_RST(n_4_net_) );
  ivd1_hd I_10 ( .A(i_RSTN), .Y(n_4_net_) );
  ivd1_hd I_9 ( .A(i_RSTN), .Y(n_3_net_) );
  ivd1_hd I_8 ( .A(i_RSTN), .Y(n_2_net_) );
  ivd1_hd U833 ( .A(i_RSTN), .Y(N23) );
  fd2qd1_hd r_counter_reg_1_ ( .D(n791), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_counter_1_) );
  fd1eqd1_hd r_mult_3_AB_STB_reg ( .D(N1343), .E(N1403), .CK(i_CLK), .Q(
        r_mult_3_AB_STB) );
  fd2qd1_hd r_mult_3_Z_ACK_reg ( .D(n497), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_Z_ACK) );
  fd2qd1_hd r_mult_1_AB_STB_reg ( .D(n491), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_AB_STB) );
  fd2qd1_hd r_mult_2_AB_STB_reg ( .D(n490), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_AB_STB) );
  fd2qd1_hd r_mult_2_A_reg_2_ ( .D(n169), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[2]) );
  fd2qd1_hd r_mult_2_A_reg_11_ ( .D(n160), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[11]) );
  fd2qd1_hd r_mult_2_A_reg_16_ ( .D(n155), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[16]) );
  fd2qd1_hd r_mult_2_A_reg_23_ ( .D(n148), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[23]) );
  fd2qd1_hd r_mult_2_A_reg_30_ ( .D(n141), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[30]) );
  fd2qd1_hd r_mult_3_A_reg_30_ ( .D(n78), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[30]) );
  fd2qd1_hd r_mult_2_A_reg_1_ ( .D(n170), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[1]) );
  fd2qd1_hd r_mult_2_A_reg_4_ ( .D(n167), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[4]) );
  fd2qd1_hd r_mult_2_A_reg_7_ ( .D(n164), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[7]) );
  fd2qd1_hd r_mult_2_A_reg_9_ ( .D(n162), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[9]) );
  fd2qd1_hd r_mult_2_A_reg_13_ ( .D(n158), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[13]) );
  fd2qd1_hd r_mult_2_A_reg_14_ ( .D(n157), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[14]) );
  fd2qd1_hd r_mult_2_A_reg_19_ ( .D(n152), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[19]) );
  fd2qd1_hd r_mult_2_A_reg_20_ ( .D(n151), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[20]) );
  fd2qd1_hd r_mult_2_A_reg_21_ ( .D(n150), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[21]) );
  fd2qd1_hd r_mult_2_A_reg_31_ ( .D(n140), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[31]) );
  fd2qd1_hd r_mult_3_A_reg_2_ ( .D(n106), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[2]) );
  fd2qd1_hd r_mult_3_A_reg_10_ ( .D(n98), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[10]) );
  fd2qd1_hd r_mult_3_A_reg_11_ ( .D(n97), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[11]) );
  fd2qd1_hd r_mult_3_A_reg_15_ ( .D(n93), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[15]) );
  fd2qd1_hd r_mult_3_A_reg_18_ ( .D(n90), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[18]) );
  fd2qd1_hd r_mult_3_A_reg_21_ ( .D(n87), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[21]) );
  fd2qd1_hd r_mult_3_A_reg_22_ ( .D(n86), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[22]) );
  fd2qd1_hd r_mult_3_A_reg_23_ ( .D(n85), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[23]) );
  fd2qd1_hd r_mult_3_A_reg_24_ ( .D(n84), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[24]) );
  fd2qd1_hd r_mult_3_A_reg_31_ ( .D(n77), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[31]) );
  fd2qd1_hd r_mult_3_B_reg_31_ ( .D(n501), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[31]) );
  fd2qd1_hd r_mult_3_B_reg_0_ ( .D(n139), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[0]) );
  fd2qd1_hd r_mult_3_B_reg_1_ ( .D(n138), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[1]) );
  fd2qd1_hd r_mult_3_B_reg_2_ ( .D(n137), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[2]) );
  fd2qd1_hd r_mult_3_B_reg_3_ ( .D(n136), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[3]) );
  fd2qd1_hd r_mult_3_B_reg_4_ ( .D(n135), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[4]) );
  fd2qd1_hd r_mult_3_B_reg_5_ ( .D(n134), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[5]) );
  fd2qd1_hd r_mult_3_B_reg_6_ ( .D(n133), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[6]) );
  fd2qd1_hd r_mult_3_B_reg_7_ ( .D(n132), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[7]) );
  fd2qd1_hd r_mult_3_B_reg_8_ ( .D(n131), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[8]) );
  fd2qd1_hd r_mult_3_B_reg_9_ ( .D(n130), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[9]) );
  fd2qd1_hd r_mult_3_B_reg_10_ ( .D(n129), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[10]) );
  fd2qd1_hd r_mult_3_B_reg_11_ ( .D(n128), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[11]) );
  fd2qd1_hd r_mult_3_B_reg_12_ ( .D(n127), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[12]) );
  fd2qd1_hd r_mult_3_B_reg_13_ ( .D(n126), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[13]) );
  fd2qd1_hd r_mult_3_B_reg_14_ ( .D(n125), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[14]) );
  fd2qd1_hd r_mult_3_B_reg_15_ ( .D(n124), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[15]) );
  fd2qd1_hd r_mult_3_B_reg_16_ ( .D(n123), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[16]) );
  fd2qd1_hd r_mult_3_B_reg_17_ ( .D(n122), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[17]) );
  fd2qd1_hd r_mult_3_B_reg_18_ ( .D(n121), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[18]) );
  fd2qd1_hd r_mult_3_B_reg_19_ ( .D(n120), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[19]) );
  fd2qd1_hd r_mult_3_B_reg_20_ ( .D(n119), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[20]) );
  fd2qd1_hd r_mult_3_B_reg_21_ ( .D(n118), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[21]) );
  fd2qd1_hd r_mult_3_B_reg_22_ ( .D(n117), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[22]) );
  fd2qd1_hd r_mult_3_B_reg_23_ ( .D(n116), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[23]) );
  fd2qd1_hd r_mult_3_B_reg_24_ ( .D(n115), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[24]) );
  fd2qd1_hd r_mult_3_B_reg_25_ ( .D(n114), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[25]) );
  fd2qd1_hd r_mult_3_B_reg_26_ ( .D(n113), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[26]) );
  fd2qd1_hd r_mult_3_B_reg_27_ ( .D(n112), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[27]) );
  fd2qd1_hd r_mult_3_B_reg_28_ ( .D(n111), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[28]) );
  fd2qd1_hd r_mult_3_B_reg_29_ ( .D(n110), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[29]) );
  fd2qd1_hd r_mult_3_B_reg_30_ ( .D(n109), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_0_ ( .D(n76), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[0]) );
  fd2qd1_hd r_mult_1_B_reg_1_ ( .D(n75), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[1]) );
  fd2qd1_hd r_mult_1_B_reg_2_ ( .D(n74), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[2]) );
  fd2qd1_hd r_mult_1_B_reg_3_ ( .D(n73), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[3]) );
  fd2qd1_hd r_mult_1_B_reg_4_ ( .D(n72), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[4]) );
  fd2qd1_hd r_mult_1_B_reg_5_ ( .D(n71), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[5]) );
  fd2qd1_hd r_mult_1_B_reg_6_ ( .D(n70), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[6]) );
  fd2qd1_hd r_mult_1_B_reg_7_ ( .D(n69), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[7]) );
  fd2qd1_hd r_mult_1_B_reg_8_ ( .D(n68), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[8]) );
  fd2qd1_hd r_mult_1_B_reg_9_ ( .D(n67), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[9]) );
  fd2qd1_hd r_mult_1_B_reg_10_ ( .D(n66), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[10]) );
  fd2qd1_hd r_mult_1_B_reg_11_ ( .D(n65), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[11]) );
  fd2qd1_hd r_mult_1_B_reg_12_ ( .D(n64), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[12]) );
  fd2qd1_hd r_mult_1_B_reg_13_ ( .D(n63), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[13]) );
  fd2qd1_hd r_mult_1_B_reg_14_ ( .D(n62), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[14]) );
  fd2qd1_hd r_mult_1_B_reg_15_ ( .D(n61), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[15]) );
  fd2qd1_hd r_mult_1_B_reg_16_ ( .D(n60), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[16]) );
  fd2qd1_hd r_mult_1_B_reg_17_ ( .D(n59), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[17]) );
  fd2qd1_hd r_mult_1_B_reg_18_ ( .D(n58), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[18]) );
  fd2qd1_hd r_mult_1_B_reg_19_ ( .D(n57), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[19]) );
  fd2qd1_hd r_mult_1_B_reg_20_ ( .D(n56), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[20]) );
  fd2qd1_hd r_mult_1_B_reg_21_ ( .D(n55), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[21]) );
  fd2qd1_hd r_mult_1_B_reg_22_ ( .D(n54), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[22]) );
  fd2qd1_hd r_mult_1_B_reg_30_ ( .D(n46), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[30]) );
  fd2qd1_hd r_mult_1_B_reg_31_ ( .D(n45), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[31]) );
  fd2qd1_hd r_mult_2_B_reg_31_ ( .D(n499), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[31]) );
  fd2qd1_hd r_mult_1_Z_ACK_reg ( .D(n493), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_Z_ACK) );
  fd2qd1_hd r_mult_2_Z_ACK_reg ( .D(n492), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_Z_ACK) );
  fd2qd1_hd r_mult_2_B_reg_0_ ( .D(n202), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[0]) );
  fd2qd1_hd r_mult_2_B_reg_1_ ( .D(n201), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[1]) );
  fd2qd1_hd r_mult_2_B_reg_2_ ( .D(n200), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[2]) );
  fd2qd1_hd r_mult_2_B_reg_3_ ( .D(n199), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[3]) );
  fd2qd1_hd r_mult_2_B_reg_4_ ( .D(n198), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[4]) );
  fd2qd1_hd r_mult_2_B_reg_5_ ( .D(n197), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[5]) );
  fd2qd1_hd r_mult_2_B_reg_6_ ( .D(n196), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[6]) );
  fd2qd1_hd r_mult_2_B_reg_7_ ( .D(n195), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[7]) );
  fd2qd1_hd r_mult_2_B_reg_8_ ( .D(n194), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[8]) );
  fd2qd1_hd r_mult_2_B_reg_9_ ( .D(n193), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[9]) );
  fd2qd1_hd r_mult_2_B_reg_10_ ( .D(n192), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[10]) );
  fd2qd1_hd r_mult_2_B_reg_11_ ( .D(n191), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[11]) );
  fd2qd1_hd r_mult_2_B_reg_12_ ( .D(n190), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[12]) );
  fd2qd1_hd r_mult_2_B_reg_13_ ( .D(n189), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[13]) );
  fd2qd1_hd r_mult_2_B_reg_14_ ( .D(n188), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[14]) );
  fd2qd1_hd r_mult_2_B_reg_15_ ( .D(n187), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[15]) );
  fd2qd1_hd r_mult_2_B_reg_16_ ( .D(n186), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[16]) );
  fd2qd1_hd r_mult_2_B_reg_17_ ( .D(n185), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[17]) );
  fd2qd1_hd r_mult_2_B_reg_18_ ( .D(n184), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[18]) );
  fd2qd1_hd r_mult_2_B_reg_19_ ( .D(n183), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[19]) );
  fd2qd1_hd r_mult_2_B_reg_20_ ( .D(n182), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[20]) );
  fd2qd1_hd r_mult_2_B_reg_21_ ( .D(n181), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[21]) );
  fd2qd1_hd r_mult_2_B_reg_22_ ( .D(n180), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[22]) );
  fd2qd1_hd r_mult_2_B_reg_23_ ( .D(n179), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[23]) );
  fd2qd1_hd r_mult_2_B_reg_24_ ( .D(n178), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[24]) );
  fd2qd1_hd r_mult_2_B_reg_25_ ( .D(n177), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[25]) );
  fd2qd1_hd r_mult_2_B_reg_26_ ( .D(n176), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[26]) );
  fd2qd1_hd r_mult_2_B_reg_27_ ( .D(n175), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[27]) );
  fd2qd1_hd r_mult_2_B_reg_28_ ( .D(n174), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[28]) );
  fd2qd1_hd r_mult_2_B_reg_29_ ( .D(n173), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[29]) );
  fd2qd1_hd r_mult_2_B_reg_30_ ( .D(n172), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_B[30]) );
  fd2qd1_hd r_mult_2_A_reg_12_ ( .D(n159), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[12]) );
  fd2qd1_hd r_mult_2_A_reg_18_ ( .D(n153), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[18]) );
  fd2qd1_hd r_mult_1_B_reg_23_ ( .D(n53), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[23]) );
  fd2qd1_hd r_mult_1_B_reg_24_ ( .D(n52), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[24]) );
  fd2qd1_hd r_mult_1_B_reg_25_ ( .D(n51), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[25]) );
  fd2qd1_hd r_mult_1_B_reg_26_ ( .D(n50), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[26]) );
  fd2qd1_hd r_mult_1_B_reg_27_ ( .D(n49), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[27]) );
  fd2qd1_hd r_mult_1_B_reg_28_ ( .D(n48), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[28]) );
  fd2qd1_hd r_mult_1_B_reg_29_ ( .D(n47), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_B[29]) );
  fd2qd1_hd r_mult_2_A_reg_0_ ( .D(n171), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[0]) );
  fd2qd1_hd r_mult_2_A_reg_5_ ( .D(n166), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[5]) );
  fd2qd1_hd r_mult_2_A_reg_15_ ( .D(n156), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[15]) );
  fd2qd1_hd r_mult_2_A_reg_17_ ( .D(n154), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[17]) );
  fd2qd1_hd r_mult_2_A_reg_24_ ( .D(n147), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[24]) );
  fd2qd1_hd r_mult_3_A_reg_0_ ( .D(n108), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[0]) );
  fd2qd1_hd r_mult_3_A_reg_1_ ( .D(n107), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[1]) );
  fd2qd1_hd r_mult_3_A_reg_6_ ( .D(n102), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[6]) );
  fd2qd1_hd r_mult_3_A_reg_8_ ( .D(n100), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[8]) );
  fd2qd1_hd r_mult_3_A_reg_9_ ( .D(n99), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[9]) );
  fd2qd1_hd r_mult_3_A_reg_13_ ( .D(n95), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[13]) );
  fd2qd1_hd r_mult_3_A_reg_14_ ( .D(n94), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[14]) );
  fd2qd1_hd r_mult_3_A_reg_16_ ( .D(n92), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[16]) );
  fd2qd1_hd r_mult_3_A_reg_19_ ( .D(n89), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[19]) );
  fd2qd1_hd r_mult_3_A_reg_20_ ( .D(n88), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[20]) );
  fd2qd1_hd r_mult_2_A_reg_3_ ( .D(n168), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[3]) );
  fd2qd1_hd r_mult_2_A_reg_6_ ( .D(n165), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[6]) );
  fd2qd1_hd r_mult_2_A_reg_8_ ( .D(n163), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[8]) );
  fd2qd1_hd r_mult_2_A_reg_10_ ( .D(n161), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[10]) );
  fd2qd1_hd r_mult_2_A_reg_22_ ( .D(n149), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[22]) );
  fd2qd1_hd r_mult_2_A_reg_25_ ( .D(n146), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[25]) );
  fd2qd1_hd r_mult_2_A_reg_26_ ( .D(n145), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[26]) );
  fd2qd1_hd r_mult_2_A_reg_27_ ( .D(n144), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[27]) );
  fd2qd1_hd r_mult_2_A_reg_28_ ( .D(n143), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[28]) );
  fd2qd1_hd r_mult_2_A_reg_29_ ( .D(n142), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_2_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_0_ ( .D(n502), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[0]) );
  fd2qd1_hd r_mult_1_A_reg_2_ ( .D(n43), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[2]) );
  fd2qd1_hd r_mult_1_A_reg_3_ ( .D(n42), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[3]) );
  fd2qd1_hd r_mult_1_A_reg_4_ ( .D(n41), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[4]) );
  fd2qd1_hd r_mult_1_A_reg_5_ ( .D(n40), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[5]) );
  fd2qd1_hd r_mult_1_A_reg_7_ ( .D(n38), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[7]) );
  fd2qd1_hd r_mult_1_A_reg_10_ ( .D(n35), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[10]) );
  fd2qd1_hd r_mult_1_A_reg_11_ ( .D(n34), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[11]) );
  fd2qd1_hd r_mult_1_A_reg_13_ ( .D(n32), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[13]) );
  fd2qd1_hd r_mult_1_A_reg_14_ ( .D(n31), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[14]) );
  fd2qd1_hd r_mult_1_A_reg_15_ ( .D(n30), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[15]) );
  fd2qd1_hd r_mult_1_A_reg_17_ ( .D(n28), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[17]) );
  fd2qd1_hd r_mult_1_A_reg_18_ ( .D(n27), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[18]) );
  fd2qd1_hd r_mult_1_A_reg_19_ ( .D(n26), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[19]) );
  fd2qd1_hd r_mult_1_A_reg_21_ ( .D(n24), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[21]) );
  fd2qd1_hd r_mult_1_A_reg_22_ ( .D(n23), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[22]) );
  fd2qd1_hd r_mult_1_A_reg_23_ ( .D(n22), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[23]) );
  fd2qd1_hd r_mult_1_A_reg_24_ ( .D(n21), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[24]) );
  fd2qd1_hd r_mult_1_A_reg_25_ ( .D(n20), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[25]) );
  fd2qd1_hd r_mult_1_A_reg_26_ ( .D(n19), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[26]) );
  fd2qd1_hd r_mult_1_A_reg_27_ ( .D(n18), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[27]) );
  fd2qd1_hd r_mult_1_A_reg_28_ ( .D(n17), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[28]) );
  fd2qd1_hd r_mult_1_A_reg_29_ ( .D(n16), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[29]) );
  fd2qd1_hd r_mult_1_A_reg_1_ ( .D(n44), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[1]) );
  fd2qd1_hd r_mult_1_A_reg_6_ ( .D(n39), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[6]) );
  fd2qd1_hd r_mult_1_A_reg_8_ ( .D(n37), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[8]) );
  fd2qd1_hd r_mult_1_A_reg_9_ ( .D(n36), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[9]) );
  fd2qd1_hd r_mult_1_A_reg_12_ ( .D(n33), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[12]) );
  fd2qd1_hd r_mult_1_A_reg_16_ ( .D(n29), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[16]) );
  fd2qd1_hd r_mult_1_A_reg_20_ ( .D(n25), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[20]) );
  fd2qd1_hd r_mult_1_A_reg_30_ ( .D(n15), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[30]) );
  fd2qd1_hd r_mult_1_A_reg_31_ ( .D(n14), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_1_A[31]) );
  fd2qd1_hd r_add_2_B_reg_31_ ( .D(n794), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[31]) );
  fd2qd1_hd r_add_1_B_reg_19_ ( .D(n672), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[19]) );
  fd2qd1_hd r_add_2_B_reg_0_ ( .D(n755), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[0]) );
  fd2qd1_hd r_add_2_A_reg_0_ ( .D(n723), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[0]) );
  fd2qd1_hd r_add_2_B_reg_1_ ( .D(n754), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[1]) );
  fd2qd1_hd r_add_2_A_reg_1_ ( .D(n722), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[1]) );
  fd2qd1_hd r_add_2_B_reg_2_ ( .D(n753), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[2]) );
  fd2qd1_hd r_add_2_A_reg_2_ ( .D(n721), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[2]) );
  fd2qd1_hd r_add_2_B_reg_3_ ( .D(n752), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[3]) );
  fd2qd1_hd r_add_2_A_reg_3_ ( .D(n720), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[3]) );
  fd2qd1_hd r_add_2_B_reg_4_ ( .D(n751), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[4]) );
  fd2qd1_hd r_add_2_A_reg_4_ ( .D(n719), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[4]) );
  fd2qd1_hd r_add_2_B_reg_5_ ( .D(n750), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[5]) );
  fd2qd1_hd r_add_2_A_reg_5_ ( .D(n718), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[5]) );
  fd2qd1_hd r_add_2_B_reg_6_ ( .D(n749), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[6]) );
  fd2qd1_hd r_add_2_A_reg_6_ ( .D(n717), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[6]) );
  fd2qd1_hd r_add_2_B_reg_7_ ( .D(n748), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[7]) );
  fd2qd1_hd r_add_2_A_reg_7_ ( .D(n716), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[7]) );
  fd2qd1_hd r_add_2_B_reg_8_ ( .D(n747), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[8]) );
  fd2qd1_hd r_add_2_A_reg_8_ ( .D(n715), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[8]) );
  fd2qd1_hd r_add_2_B_reg_9_ ( .D(n746), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[9]) );
  fd2qd1_hd r_add_2_A_reg_9_ ( .D(n714), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[9]) );
  fd2qd1_hd r_add_2_B_reg_10_ ( .D(n745), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[10]) );
  fd2qd1_hd r_add_2_A_reg_10_ ( .D(n713), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[10]) );
  fd2qd1_hd r_add_2_B_reg_11_ ( .D(n744), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[11]) );
  fd2qd1_hd r_add_2_A_reg_11_ ( .D(n712), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[11]) );
  fd2qd1_hd r_add_2_B_reg_12_ ( .D(n743), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[12]) );
  fd2qd1_hd r_add_2_A_reg_12_ ( .D(n711), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[12]) );
  fd2qd1_hd r_add_2_B_reg_13_ ( .D(n742), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[13]) );
  fd2qd1_hd r_add_2_A_reg_13_ ( .D(n710), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[13]) );
  fd2qd1_hd r_add_2_B_reg_14_ ( .D(n741), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[14]) );
  fd2qd1_hd r_add_2_A_reg_14_ ( .D(n709), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[14]) );
  fd2qd1_hd r_add_2_B_reg_15_ ( .D(n740), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[15]) );
  fd2qd1_hd r_add_2_A_reg_15_ ( .D(n708), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[15]) );
  fd2qd1_hd r_add_2_B_reg_16_ ( .D(n739), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[16]) );
  fd2qd1_hd r_add_2_A_reg_16_ ( .D(n707), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[16]) );
  fd2qd1_hd r_add_2_B_reg_17_ ( .D(n738), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[17]) );
  fd2qd1_hd r_add_2_A_reg_17_ ( .D(n706), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[17]) );
  fd2qd1_hd r_add_2_B_reg_18_ ( .D(n737), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[18]) );
  fd2qd1_hd r_add_2_A_reg_18_ ( .D(n705), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[18]) );
  fd2qd1_hd r_add_2_B_reg_19_ ( .D(n736), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[19]) );
  fd2qd1_hd r_add_2_A_reg_19_ ( .D(n704), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[19]) );
  fd2qd1_hd r_add_2_B_reg_20_ ( .D(n735), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[20]) );
  fd2qd1_hd r_add_2_A_reg_20_ ( .D(n703), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[20]) );
  fd2qd1_hd r_add_2_B_reg_21_ ( .D(n734), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[21]) );
  fd2qd1_hd r_add_2_A_reg_21_ ( .D(n702), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[21]) );
  fd2qd1_hd r_add_2_B_reg_22_ ( .D(n733), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[22]) );
  fd2qd1_hd r_add_2_A_reg_22_ ( .D(n701), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[22]) );
  fd2qd1_hd r_add_2_B_reg_23_ ( .D(n732), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[23]) );
  fd2qd1_hd r_add_2_A_reg_23_ ( .D(n700), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[23]) );
  fd2qd1_hd r_add_2_B_reg_24_ ( .D(n731), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[24]) );
  fd2qd1_hd r_add_2_A_reg_24_ ( .D(n699), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[24]) );
  fd2qd1_hd r_add_2_B_reg_25_ ( .D(n730), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[25]) );
  fd2qd1_hd r_add_2_A_reg_25_ ( .D(n698), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[25]) );
  fd2qd1_hd r_add_2_B_reg_26_ ( .D(n729), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[26]) );
  fd2qd1_hd r_add_2_A_reg_26_ ( .D(n697), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[26]) );
  fd2qd1_hd r_add_2_B_reg_27_ ( .D(n728), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[27]) );
  fd2qd1_hd r_add_2_A_reg_27_ ( .D(n696), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[27]) );
  fd2qd1_hd r_add_2_B_reg_28_ ( .D(n727), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[28]) );
  fd2qd1_hd r_add_2_A_reg_28_ ( .D(n695), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[28]) );
  fd2qd1_hd r_add_2_B_reg_29_ ( .D(n726), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[29]) );
  fd2qd1_hd r_add_2_A_reg_29_ ( .D(n694), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[29]) );
  fd2qd1_hd r_add_2_B_reg_30_ ( .D(n725), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_B[30]) );
  fd2qd1_hd r_add_2_A_reg_30_ ( .D(n693), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[30]) );
  fd2qd1_hd r_add_2_A_reg_31_ ( .D(n692), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_A[31]) );
  fd2qd1_hd r_add_1_B_reg_31_ ( .D(n660), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[31]) );
  fd2qd1_hd r_add_1_B_reg_0_ ( .D(n691), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[0]) );
  fd2qd1_hd r_add_1_B_reg_1_ ( .D(n690), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[1]) );
  fd2qd1_hd r_add_1_B_reg_2_ ( .D(n689), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[2]) );
  fd2qd1_hd r_add_1_B_reg_3_ ( .D(n688), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[3]) );
  fd2qd1_hd r_add_1_B_reg_4_ ( .D(n687), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[4]) );
  fd2qd1_hd r_add_1_B_reg_5_ ( .D(n686), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[5]) );
  fd2qd1_hd r_add_1_B_reg_6_ ( .D(n685), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[6]) );
  fd2qd1_hd r_add_1_B_reg_7_ ( .D(n684), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[7]) );
  fd2qd1_hd r_add_1_B_reg_8_ ( .D(n683), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[8]) );
  fd2qd1_hd r_add_1_B_reg_9_ ( .D(n682), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[9]) );
  fd2qd1_hd r_add_1_B_reg_10_ ( .D(n681), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[10]) );
  fd2qd1_hd r_add_1_B_reg_11_ ( .D(n680), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[11]) );
  fd2qd1_hd r_add_1_B_reg_12_ ( .D(n679), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[12]) );
  fd2qd1_hd r_add_1_B_reg_13_ ( .D(n678), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[13]) );
  fd2qd1_hd r_add_1_B_reg_14_ ( .D(n677), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[14]) );
  fd2qd1_hd r_add_1_B_reg_15_ ( .D(n676), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[15]) );
  fd2qd1_hd r_add_1_B_reg_16_ ( .D(n675), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[16]) );
  fd2qd1_hd r_add_1_B_reg_17_ ( .D(n674), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[17]) );
  fd2qd1_hd r_add_1_B_reg_18_ ( .D(n673), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[18]) );
  fd2qd1_hd r_add_1_B_reg_20_ ( .D(n671), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[20]) );
  fd2qd1_hd r_add_1_B_reg_21_ ( .D(n670), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[21]) );
  fd2qd1_hd r_add_1_B_reg_22_ ( .D(n669), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[22]) );
  fd2qd1_hd r_add_1_B_reg_23_ ( .D(n668), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[23]) );
  fd2qd1_hd r_add_1_B_reg_24_ ( .D(n667), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[24]) );
  fd2qd1_hd r_add_1_B_reg_25_ ( .D(n666), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[25]) );
  fd2qd1_hd r_add_1_B_reg_26_ ( .D(n665), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[26]) );
  fd2qd1_hd r_add_1_B_reg_27_ ( .D(n664), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[27]) );
  fd2qd1_hd r_add_1_B_reg_28_ ( .D(n663), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[28]) );
  fd2qd1_hd r_add_1_B_reg_29_ ( .D(n662), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[29]) );
  fd2qd1_hd r_add_1_B_reg_30_ ( .D(n661), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_B[30]) );
  fd2qd1_hd r_x_data_reg_147_ ( .D(n342), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[147]) );
  fd2qd1_hd r_x_data_reg_128_ ( .D(n361), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[128]) );
  fd2qd1_hd r_x_data_reg_129_ ( .D(n360), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[129]) );
  fd2qd1_hd r_x_data_reg_130_ ( .D(n359), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[130]) );
  fd2qd1_hd r_x_data_reg_131_ ( .D(n358), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[131]) );
  fd2qd1_hd r_x_data_reg_132_ ( .D(n357), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[132]) );
  fd2qd1_hd r_x_data_reg_133_ ( .D(n356), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[133]) );
  fd2qd1_hd r_x_data_reg_134_ ( .D(n355), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[134]) );
  fd2qd1_hd r_x_data_reg_135_ ( .D(n354), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[135]) );
  fd2qd1_hd r_x_data_reg_136_ ( .D(n353), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[136]) );
  fd2qd1_hd r_x_data_reg_137_ ( .D(n352), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[137]) );
  fd2qd1_hd r_x_data_reg_138_ ( .D(n351), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[138]) );
  fd2qd1_hd r_x_data_reg_139_ ( .D(n350), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[139]) );
  fd2qd1_hd r_x_data_reg_140_ ( .D(n349), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[140]) );
  fd2qd1_hd r_x_data_reg_141_ ( .D(n348), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[141]) );
  fd2qd1_hd r_x_data_reg_142_ ( .D(n347), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[142]) );
  fd2qd1_hd r_x_data_reg_143_ ( .D(n346), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[143]) );
  fd2qd1_hd r_x_data_reg_144_ ( .D(n345), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[144]) );
  fd2qd1_hd r_x_data_reg_145_ ( .D(n344), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[145]) );
  fd2qd1_hd r_x_data_reg_146_ ( .D(n343), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[146]) );
  fd2qd1_hd r_x_data_reg_148_ ( .D(n341), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[148]) );
  fd2qd1_hd r_x_data_reg_149_ ( .D(n340), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[149]) );
  fd2qd1_hd r_x_data_reg_150_ ( .D(n339), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[150]) );
  fd2qd1_hd r_x_data_reg_151_ ( .D(n338), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[151]) );
  fd2qd1_hd r_x_data_reg_152_ ( .D(n337), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[152]) );
  fd2qd1_hd r_x_data_reg_153_ ( .D(n336), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[153]) );
  fd2qd1_hd r_x_data_reg_154_ ( .D(n335), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[154]) );
  fd2qd1_hd r_x_data_reg_155_ ( .D(n334), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[155]) );
  fd2qd1_hd r_x_data_reg_156_ ( .D(n333), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[156]) );
  fd2qd1_hd r_x_data_reg_157_ ( .D(n332), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[157]) );
  fd2qd1_hd r_x_data_reg_158_ ( .D(n331), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[158]) );
  fd2qd1_hd r_x_data_reg_159_ ( .D(n330), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[159]) );
  fd2qd1_hd r_y_data_reg_96_ ( .D(n234), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[96]) );
  fd2qd1_hd r_y_data_reg_97_ ( .D(n233), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[97]) );
  fd2qd1_hd r_y_data_reg_98_ ( .D(n232), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[98]) );
  fd2qd1_hd r_y_data_reg_99_ ( .D(n231), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[99]) );
  fd2qd1_hd r_y_data_reg_100_ ( .D(n230), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[100]) );
  fd2qd1_hd r_y_data_reg_101_ ( .D(n229), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[101]) );
  fd2qd1_hd r_y_data_reg_102_ ( .D(n228), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[102]) );
  fd2qd1_hd r_y_data_reg_103_ ( .D(n227), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[103]) );
  fd2qd1_hd r_y_data_reg_104_ ( .D(n226), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[104]) );
  fd2qd1_hd r_y_data_reg_105_ ( .D(n225), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[105]) );
  fd2qd1_hd r_y_data_reg_106_ ( .D(n224), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[106]) );
  fd2qd1_hd r_y_data_reg_107_ ( .D(n223), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[107]) );
  fd2qd1_hd r_y_data_reg_108_ ( .D(n222), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[108]) );
  fd2qd1_hd r_y_data_reg_109_ ( .D(n221), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[109]) );
  fd2qd1_hd r_y_data_reg_110_ ( .D(n220), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[110]) );
  fd2qd1_hd r_y_data_reg_111_ ( .D(n219), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[111]) );
  fd2qd1_hd r_y_data_reg_112_ ( .D(n218), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[112]) );
  fd2qd1_hd r_y_data_reg_113_ ( .D(n217), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[113]) );
  fd2qd1_hd r_y_data_reg_114_ ( .D(n216), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[114]) );
  fd2qd1_hd r_y_data_reg_115_ ( .D(n215), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[115]) );
  fd2qd1_hd r_y_data_reg_116_ ( .D(n214), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[116]) );
  fd2qd1_hd r_y_data_reg_117_ ( .D(n213), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[117]) );
  fd2qd1_hd r_y_data_reg_118_ ( .D(n212), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[118]) );
  fd2qd1_hd r_y_data_reg_119_ ( .D(n211), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[119]) );
  fd2qd1_hd r_y_data_reg_120_ ( .D(n210), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[120]) );
  fd2qd1_hd r_y_data_reg_121_ ( .D(n209), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[121]) );
  fd2qd1_hd r_y_data_reg_122_ ( .D(n208), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[122]) );
  fd2qd1_hd r_y_data_reg_123_ ( .D(n207), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[123]) );
  fd2qd1_hd r_y_data_reg_124_ ( .D(n206), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[124]) );
  fd2qd1_hd r_y_data_reg_125_ ( .D(n205), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[125]) );
  fd2qd1_hd r_y_data_reg_126_ ( .D(n204), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[126]) );
  fd2qd1_hd r_y_data_reg_127_ ( .D(n203), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[127]) );
  fd2qd1_hd r_add_1_A_reg_0_ ( .D(n787), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[0]) );
  fd2qd1_hd r_add_1_A_reg_1_ ( .D(n786), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[1]) );
  fd2qd1_hd r_add_1_A_reg_2_ ( .D(n785), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[2]) );
  fd2qd1_hd r_add_1_A_reg_3_ ( .D(n784), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[3]) );
  fd2qd1_hd r_add_1_A_reg_4_ ( .D(n783), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[4]) );
  fd2qd1_hd r_add_1_A_reg_5_ ( .D(n782), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[5]) );
  fd2qd1_hd r_add_1_A_reg_6_ ( .D(n781), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[6]) );
  fd2qd1_hd r_add_1_A_reg_7_ ( .D(n780), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[7]) );
  fd2qd1_hd r_add_1_A_reg_8_ ( .D(n779), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[8]) );
  fd2qd1_hd r_add_1_A_reg_9_ ( .D(n778), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[9]) );
  fd2qd1_hd r_add_1_A_reg_10_ ( .D(n777), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[10]) );
  fd2qd1_hd r_add_1_A_reg_11_ ( .D(n776), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[11]) );
  fd2qd1_hd r_add_1_A_reg_12_ ( .D(n775), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[12]) );
  fd2qd1_hd r_add_1_A_reg_13_ ( .D(n774), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[13]) );
  fd2qd1_hd r_add_1_A_reg_14_ ( .D(n773), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[14]) );
  fd2qd1_hd r_add_1_A_reg_15_ ( .D(n772), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[15]) );
  fd2qd1_hd r_add_1_A_reg_16_ ( .D(n771), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[16]) );
  fd2qd1_hd r_add_1_A_reg_17_ ( .D(n770), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[17]) );
  fd2qd1_hd r_add_1_A_reg_18_ ( .D(n769), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[18]) );
  fd2qd1_hd r_add_1_A_reg_19_ ( .D(n768), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[19]) );
  fd2qd1_hd r_add_1_A_reg_20_ ( .D(n767), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[20]) );
  fd2qd1_hd r_add_1_A_reg_21_ ( .D(n766), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[21]) );
  fd2qd1_hd r_add_1_A_reg_22_ ( .D(n765), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[22]) );
  fd2qd1_hd r_add_1_A_reg_23_ ( .D(n764), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[23]) );
  fd2qd1_hd r_add_1_A_reg_24_ ( .D(n763), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[24]) );
  fd2qd1_hd r_add_1_A_reg_25_ ( .D(n762), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[25]) );
  fd2qd1_hd r_add_1_A_reg_26_ ( .D(n761), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[26]) );
  fd2qd1_hd r_add_1_A_reg_27_ ( .D(n760), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[27]) );
  fd2qd1_hd r_add_1_A_reg_28_ ( .D(n759), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[28]) );
  fd2qd1_hd r_add_1_A_reg_29_ ( .D(n758), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[29]) );
  fd2qd1_hd r_add_1_A_reg_30_ ( .D(n757), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[30]) );
  fd2qd1_hd r_add_1_A_reg_31_ ( .D(n826), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_A[31]) );
  fd2qd1_hd r_mult_3_A_reg_3_ ( .D(n105), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[3]) );
  fd2qd1_hd r_mult_3_A_reg_4_ ( .D(n104), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[4]) );
  fd2qd1_hd r_mult_3_A_reg_5_ ( .D(n103), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[5]) );
  fd2qd1_hd r_mult_3_A_reg_7_ ( .D(n101), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[7]) );
  fd2qd1_hd r_mult_3_A_reg_12_ ( .D(n96), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[12]) );
  fd2qd1_hd r_mult_3_A_reg_17_ ( .D(n91), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[17]) );
  fd2qd1_hd r_mult_3_A_reg_25_ ( .D(n83), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[25]) );
  fd2qd1_hd r_mult_3_A_reg_26_ ( .D(n82), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[26]) );
  fd2qd1_hd r_mult_3_A_reg_27_ ( .D(n81), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[27]) );
  fd2qd1_hd r_mult_3_A_reg_28_ ( .D(n80), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[28]) );
  fd2qd1_hd r_mult_3_A_reg_29_ ( .D(n79), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_3_A[29]) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(n827), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[31]) );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(n795), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[0]) );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(n796), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[1]) );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(n797), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[2]) );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(n798), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[3]) );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(n799), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[4]) );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(n800), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[5]) );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(n801), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[6]) );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(n802), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[7]) );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(n803), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[8]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(n804), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[9]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(n805), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(n806), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(n807), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(n808), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(n809), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(n810), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(n811), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(n812), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(n813), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(n814), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(n815), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(n816), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(n817), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(n818), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(n819), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(n820), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(n821), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(n822), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(n823), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(n824), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(n825), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd r_x_data_reg_64_ ( .D(n425), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[64]) );
  fd2qd1_hd r_x_data_reg_65_ ( .D(n424), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[65]) );
  fd2qd1_hd r_x_data_reg_66_ ( .D(n423), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[66]) );
  fd2qd1_hd r_x_data_reg_67_ ( .D(n422), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[67]) );
  fd2qd1_hd r_x_data_reg_68_ ( .D(n421), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[68]) );
  fd2qd1_hd r_x_data_reg_69_ ( .D(n420), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[69]) );
  fd2qd1_hd r_x_data_reg_70_ ( .D(n419), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[70]) );
  fd2qd1_hd r_x_data_reg_71_ ( .D(n418), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[71]) );
  fd2qd1_hd r_x_data_reg_72_ ( .D(n417), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[72]) );
  fd2qd1_hd r_x_data_reg_73_ ( .D(n416), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[73]) );
  fd2qd1_hd r_x_data_reg_74_ ( .D(n415), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[74]) );
  fd2qd1_hd r_x_data_reg_75_ ( .D(n414), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[75]) );
  fd2qd1_hd r_x_data_reg_76_ ( .D(n413), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[76]) );
  fd2qd1_hd r_x_data_reg_77_ ( .D(n412), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[77]) );
  fd2qd1_hd r_x_data_reg_78_ ( .D(n411), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[78]) );
  fd2qd1_hd r_x_data_reg_79_ ( .D(n410), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[79]) );
  fd2qd1_hd r_x_data_reg_80_ ( .D(n409), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[80]) );
  fd2qd1_hd r_x_data_reg_81_ ( .D(n408), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[81]) );
  fd2qd1_hd r_x_data_reg_82_ ( .D(n407), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[82]) );
  fd2qd1_hd r_x_data_reg_83_ ( .D(n406), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[83]) );
  fd2qd1_hd r_x_data_reg_84_ ( .D(n405), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[84]) );
  fd2qd1_hd r_x_data_reg_85_ ( .D(n404), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[85]) );
  fd2qd1_hd r_x_data_reg_86_ ( .D(n403), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[86]) );
  fd2qd1_hd r_x_data_reg_94_ ( .D(n395), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[94]) );
  fd2qd1_hd r_x_data_reg_95_ ( .D(n394), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[95]) );
  fd2qd1_hd r_y_data_reg_64_ ( .D(n266), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[64]) );
  fd2qd1_hd r_y_data_reg_65_ ( .D(n265), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[65]) );
  fd2qd1_hd r_y_data_reg_66_ ( .D(n264), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[66]) );
  fd2qd1_hd r_y_data_reg_67_ ( .D(n263), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[67]) );
  fd2qd1_hd r_y_data_reg_68_ ( .D(n262), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[68]) );
  fd2qd1_hd r_y_data_reg_69_ ( .D(n261), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[69]) );
  fd2qd1_hd r_y_data_reg_70_ ( .D(n260), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[70]) );
  fd2qd1_hd r_y_data_reg_71_ ( .D(n259), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[71]) );
  fd2qd1_hd r_y_data_reg_72_ ( .D(n258), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[72]) );
  fd2qd1_hd r_y_data_reg_73_ ( .D(n257), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[73]) );
  fd2qd1_hd r_y_data_reg_74_ ( .D(n256), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[74]) );
  fd2qd1_hd r_y_data_reg_75_ ( .D(n255), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[75]) );
  fd2qd1_hd r_y_data_reg_76_ ( .D(n254), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[76]) );
  fd2qd1_hd r_y_data_reg_77_ ( .D(n253), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[77]) );
  fd2qd1_hd r_y_data_reg_78_ ( .D(n252), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[78]) );
  fd2qd1_hd r_y_data_reg_79_ ( .D(n251), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[79]) );
  fd2qd1_hd r_y_data_reg_80_ ( .D(n250), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[80]) );
  fd2qd1_hd r_y_data_reg_81_ ( .D(n249), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[81]) );
  fd2qd1_hd r_y_data_reg_82_ ( .D(n248), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[82]) );
  fd2qd1_hd r_y_data_reg_83_ ( .D(n247), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[83]) );
  fd2qd1_hd r_y_data_reg_84_ ( .D(n246), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[84]) );
  fd2qd1_hd r_y_data_reg_85_ ( .D(n245), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[85]) );
  fd2qd1_hd r_y_data_reg_86_ ( .D(n244), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[86]) );
  fd2qd1_hd r_y_data_reg_87_ ( .D(n243), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[87]) );
  fd2qd1_hd r_y_data_reg_88_ ( .D(n242), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[88]) );
  fd2qd1_hd r_y_data_reg_89_ ( .D(n241), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[89]) );
  fd2qd1_hd r_y_data_reg_90_ ( .D(n240), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[90]) );
  fd2qd1_hd r_y_data_reg_91_ ( .D(n239), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[91]) );
  fd2qd1_hd r_y_data_reg_92_ ( .D(n238), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[92]) );
  fd2qd1_hd r_y_data_reg_93_ ( .D(n237), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[93]) );
  fd2qd1_hd r_y_data_reg_94_ ( .D(n236), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[94]) );
  fd2qd1_hd r_y_data_reg_95_ ( .D(n235), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[95]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(n500), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_x_data_reg_32_ ( .D(n457), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[32]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(n456), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(n455), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[34]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(n454), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(n453), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(n452), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[37]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(n451), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(n450), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(n449), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(n448), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(n447), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(n446), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(n445), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(n444), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(n443), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(n442), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(n441), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(n440), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(n439), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(n438), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[51]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(n437), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(n436), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(n435), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(n434), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(n433), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(n432), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(n431), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[58]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(n430), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(n429), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(n428), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(n427), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_96_ ( .D(n393), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[96]) );
  fd2qd1_hd r_x_data_reg_97_ ( .D(n392), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[97]) );
  fd2qd1_hd r_x_data_reg_98_ ( .D(n391), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[98]) );
  fd2qd1_hd r_x_data_reg_99_ ( .D(n390), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[99]) );
  fd2qd1_hd r_x_data_reg_100_ ( .D(n389), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[100]) );
  fd2qd1_hd r_x_data_reg_101_ ( .D(n388), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[101]) );
  fd2qd1_hd r_x_data_reg_102_ ( .D(n387), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[102]) );
  fd2qd1_hd r_x_data_reg_103_ ( .D(n386), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[103]) );
  fd2qd1_hd r_x_data_reg_104_ ( .D(n385), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[104]) );
  fd2qd1_hd r_x_data_reg_105_ ( .D(n384), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[105]) );
  fd2qd1_hd r_x_data_reg_106_ ( .D(n383), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[106]) );
  fd2qd1_hd r_x_data_reg_107_ ( .D(n382), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[107]) );
  fd2qd1_hd r_x_data_reg_108_ ( .D(n381), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[108]) );
  fd2qd1_hd r_x_data_reg_109_ ( .D(n380), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[109]) );
  fd2qd1_hd r_x_data_reg_110_ ( .D(n379), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[110]) );
  fd2qd1_hd r_x_data_reg_111_ ( .D(n378), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[111]) );
  fd2qd1_hd r_x_data_reg_112_ ( .D(n377), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[112]) );
  fd2qd1_hd r_x_data_reg_113_ ( .D(n376), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[113]) );
  fd2qd1_hd r_x_data_reg_114_ ( .D(n375), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[114]) );
  fd2qd1_hd r_x_data_reg_115_ ( .D(n374), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[115]) );
  fd2qd1_hd r_x_data_reg_116_ ( .D(n373), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[116]) );
  fd2qd1_hd r_x_data_reg_117_ ( .D(n372), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[117]) );
  fd2qd1_hd r_x_data_reg_118_ ( .D(n371), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[118]) );
  fd2qd1_hd r_x_data_reg_119_ ( .D(n370), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[119]) );
  fd2qd1_hd r_x_data_reg_120_ ( .D(n369), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[120]) );
  fd2qd1_hd r_x_data_reg_121_ ( .D(n368), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[121]) );
  fd2qd1_hd r_x_data_reg_122_ ( .D(n367), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[122]) );
  fd2qd1_hd r_x_data_reg_123_ ( .D(n366), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[123]) );
  fd2qd1_hd r_x_data_reg_124_ ( .D(n365), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[124]) );
  fd2qd1_hd r_x_data_reg_125_ ( .D(n364), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[125]) );
  fd2qd1_hd r_x_data_reg_126_ ( .D(n363), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[126]) );
  fd2qd1_hd r_y_data_reg_0_ ( .D(n329), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[0]) );
  fd2qd1_hd r_y_data_reg_1_ ( .D(n328), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[1]) );
  fd2qd1_hd r_y_data_reg_2_ ( .D(n327), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[2]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(n326), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[3]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(n325), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(n324), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(n323), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(n322), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(n321), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(n320), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(n319), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(n318), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(n317), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(n316), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(n315), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(n314), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(n313), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(n312), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(n311), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(n310), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(n309), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(n308), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(n307), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(n306), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(n305), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(n304), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(n303), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(n302), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(n301), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(n300), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(n299), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_32_ ( .D(n298), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[32]) );
  fd2qd1_hd r_y_data_reg_33_ ( .D(n297), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[33]) );
  fd2qd1_hd r_y_data_reg_34_ ( .D(n296), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[34]) );
  fd2qd1_hd r_y_data_reg_35_ ( .D(n295), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[35]) );
  fd2qd1_hd r_y_data_reg_36_ ( .D(n294), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[36]) );
  fd2qd1_hd r_y_data_reg_37_ ( .D(n293), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[37]) );
  fd2qd1_hd r_y_data_reg_38_ ( .D(n292), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[38]) );
  fd2qd1_hd r_y_data_reg_39_ ( .D(n291), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[39]) );
  fd2qd1_hd r_y_data_reg_40_ ( .D(n290), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[40]) );
  fd2qd1_hd r_y_data_reg_41_ ( .D(n289), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[41]) );
  fd2qd1_hd r_y_data_reg_42_ ( .D(n288), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[42]) );
  fd2qd1_hd r_y_data_reg_43_ ( .D(n287), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[43]) );
  fd2qd1_hd r_y_data_reg_44_ ( .D(n286), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[44]) );
  fd2qd1_hd r_y_data_reg_45_ ( .D(n285), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[45]) );
  fd2qd1_hd r_y_data_reg_46_ ( .D(n284), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[46]) );
  fd2qd1_hd r_y_data_reg_47_ ( .D(n283), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[47]) );
  fd2qd1_hd r_y_data_reg_48_ ( .D(n282), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[48]) );
  fd2qd1_hd r_y_data_reg_49_ ( .D(n281), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[49]) );
  fd2qd1_hd r_y_data_reg_50_ ( .D(n280), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[50]) );
  fd2qd1_hd r_y_data_reg_51_ ( .D(n279), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[51]) );
  fd2qd1_hd r_y_data_reg_52_ ( .D(n278), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[52]) );
  fd2qd1_hd r_y_data_reg_53_ ( .D(n277), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[53]) );
  fd2qd1_hd r_y_data_reg_54_ ( .D(n276), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[54]) );
  fd2qd1_hd r_y_data_reg_55_ ( .D(n275), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[55]) );
  fd2qd1_hd r_y_data_reg_56_ ( .D(n274), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[56]) );
  fd2qd1_hd r_y_data_reg_57_ ( .D(n273), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[57]) );
  fd2qd1_hd r_y_data_reg_58_ ( .D(n272), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[58]) );
  fd2qd1_hd r_y_data_reg_59_ ( .D(n271), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[59]) );
  fd2qd1_hd r_y_data_reg_60_ ( .D(n270), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[60]) );
  fd2qd1_hd r_y_data_reg_61_ ( .D(n269), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[61]) );
  fd2qd1_hd r_y_data_reg_62_ ( .D(n268), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[62]) );
  fd2qd1_hd r_y_data_reg_63_ ( .D(n267), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[63]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(n426), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[63]) );
  fd2qd1_hd r_x_data_reg_127_ ( .D(n362), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[127]) );
  fd2qd1_hd r_x_data_reg_87_ ( .D(n402), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[87]) );
  fd2qd1_hd r_x_data_reg_88_ ( .D(n401), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[88]) );
  fd2qd1_hd r_x_data_reg_89_ ( .D(n400), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[89]) );
  fd2qd1_hd r_x_data_reg_90_ ( .D(n399), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[90]) );
  fd2qd1_hd r_x_data_reg_91_ ( .D(n398), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[91]) );
  fd2qd1_hd r_x_data_reg_92_ ( .D(n397), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[92]) );
  fd2qd1_hd r_x_data_reg_93_ ( .D(n396), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[93]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(n489), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(n488), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(n487), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(n486), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(n485), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(n484), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[5]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(n483), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(n482), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(n481), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(n480), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(n479), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(n478), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(n477), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(n476), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(n475), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(n474), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(n473), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(n472), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(n471), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(n470), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(n469), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(n468), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(n467), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(n466), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(n465), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(n464), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(n463), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(n462), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(n461), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(n460), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(n459), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(n458), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[31]) );
  fd2qd1_hd r_add_1_Z_ACK_reg ( .D(n793), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_Z_ACK) );
  fd2qd1_hd r_add_2_Z_ACK_reg ( .D(n756), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_Z_ACK) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n724), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_add_1_AB_STB_reg ( .D(n789), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_1_AB_STB) );
  fd2qd1_hd r_add_2_AB_STB_reg ( .D(n788), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_2_AB_STB) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n512), .E(N1402), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(N1383), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_pstate_0_) );
  fd3d1_hd r_pstate_reg_1_ ( .D(n498), .CK(i_CLK), .SN(i_RSTN), .Q(n11), .QN(
        n908) );
  fd3d1_hd r_counter_reg_0_ ( .D(n496), .CK(i_CLK), .SN(i_RSTN), .Q(n548), 
        .QN(n12) );
  fd3d1_hd r_counter_reg_2_ ( .D(n494), .CK(i_CLK), .SN(i_RSTN), .Q(n495), 
        .QN(n10) );
  scg14d1_hd U1024 ( .A(r_mult_3_A[9]), .B(n1260), .C(n1261), .Y(n99) );
  scg14d1_hd U1025 ( .A(r_mult_3_A[10]), .B(n1260), .C(n1269), .Y(n98) );
  scg14d1_hd U1026 ( .A(r_mult_3_A[11]), .B(n1260), .C(n1269), .Y(n97) );
  nd2bd1_hd U1027 ( .AN(r_mult_3_A[12]), .B(n1262), .Y(n96) );
  scg14d1_hd U1028 ( .A(r_mult_3_A[13]), .B(n1260), .C(n1261), .Y(n95) );
  scg14d1_hd U1029 ( .A(r_mult_3_A[14]), .B(n1260), .C(n1261), .Y(n94) );
  scg14d1_hd U1030 ( .A(r_mult_3_A[15]), .B(n1260), .C(n1269), .Y(n93) );
  scg14d1_hd U1031 ( .A(r_mult_3_A[16]), .B(n1260), .C(n1261), .Y(n92) );
  nd2bd1_hd U1032 ( .AN(r_mult_3_A[17]), .B(n1262), .Y(n91) );
  scg14d1_hd U1033 ( .A(r_mult_3_A[18]), .B(n1260), .C(n1269), .Y(n90) );
  scg14d1_hd U1034 ( .A(r_mult_3_A[19]), .B(n1260), .C(n1261), .Y(n89) );
  scg14d1_hd U1035 ( .A(r_mult_3_A[20]), .B(n1260), .C(n1261), .Y(n88) );
  scg14d1_hd U1036 ( .A(r_mult_3_A[21]), .B(n1260), .C(n1269), .Y(n87) );
  nd2bd1_hd U1037 ( .AN(r_mult_3_A[22]), .B(n1262), .Y(n86) );
  scg14d1_hd U1038 ( .A(r_mult_3_A[23]), .B(n1260), .C(n1269), .Y(n85) );
  scg14d1_hd U1039 ( .A(r_mult_3_A[24]), .B(n1260), .C(n1269), .Y(n84) );
  nd2bd1_hd U1040 ( .AN(r_mult_3_A[25]), .B(n1262), .Y(n83) );
  ao22d1_hd U1043 ( .A(n1267), .B(w_mult_2_Z[31]), .C(n1268), .D(
        w_mult_1_Z[31]), .Y(n1266) );
  nd2bd1_hd U1051 ( .AN(r_mult_3_A[26]), .B(n1262), .Y(n82) );
  nd2bd1_hd U1062 ( .AN(r_mult_3_A[27]), .B(n1262), .Y(n81) );
  nd2bd1_hd U1073 ( .AN(r_mult_3_A[28]), .B(n1262), .Y(n80) );
  scg4d1_hd U1081 ( .A(n1274), .B(r_add_2_B[31]), .C(w_mult_2_Z[31]), .D(n506), 
        .E(r_x_data[127]), .F(n509), .G(n511), .H(w_mult_3_Z[31]), .Y(n794) );
  nd2bd1_hd U1085 ( .AN(r_mult_3_A[29]), .B(n1262), .Y(n79) );
  ao22d1_hd U1089 ( .A(n1267), .B(w_mult_2_Z[0]), .C(n1268), .D(w_mult_1_Z[0]), 
        .Y(n1285) );
  ao22d1_hd U1092 ( .A(n1267), .B(w_mult_2_Z[1]), .C(n1268), .D(w_mult_1_Z[1]), 
        .Y(n1287) );
  ao22d1_hd U1095 ( .A(n1267), .B(w_mult_2_Z[2]), .C(n1268), .D(w_mult_1_Z[2]), 
        .Y(n1289) );
  ao22d1_hd U1098 ( .A(n1267), .B(w_mult_2_Z[3]), .C(n1268), .D(w_mult_1_Z[3]), 
        .Y(n1291) );
  ao22d1_hd U1101 ( .A(n1267), .B(w_mult_2_Z[4]), .C(n1268), .D(w_mult_1_Z[4]), 
        .Y(n1293) );
  ao22d1_hd U1104 ( .A(n1267), .B(w_mult_2_Z[5]), .C(n1268), .D(w_mult_1_Z[5]), 
        .Y(n1295) );
  ao22d1_hd U1107 ( .A(n1267), .B(w_mult_2_Z[6]), .C(n1268), .D(w_mult_1_Z[6]), 
        .Y(n1297) );
  ao22d1_hd U1110 ( .A(n1267), .B(w_mult_2_Z[7]), .C(n1268), .D(w_mult_1_Z[7]), 
        .Y(n1299) );
  ad2d1_hd U1112 ( .A(r_mult_3_A[30]), .B(n1260), .Y(n78) );
  ao22d1_hd U1114 ( .A(n1267), .B(w_mult_2_Z[8]), .C(n1268), .D(w_mult_1_Z[8]), 
        .Y(n1301) );
  ao22d1_hd U1117 ( .A(n1267), .B(w_mult_2_Z[9]), .C(n1268), .D(w_mult_1_Z[9]), 
        .Y(n1303) );
  ao22d1_hd U1120 ( .A(n1267), .B(w_mult_2_Z[10]), .C(n1268), .D(
        w_mult_1_Z[10]), .Y(n1305) );
  ao22d1_hd U1123 ( .A(n1267), .B(w_mult_2_Z[11]), .C(n1268), .D(
        w_mult_1_Z[11]), .Y(n1307) );
  ao22d1_hd U1126 ( .A(n1267), .B(w_mult_2_Z[12]), .C(n1268), .D(
        w_mult_1_Z[12]), .Y(n1309) );
  ao22d1_hd U1129 ( .A(n1267), .B(w_mult_2_Z[13]), .C(n1268), .D(
        w_mult_1_Z[13]), .Y(n1311) );
  ao22d1_hd U1132 ( .A(n1267), .B(w_mult_2_Z[14]), .C(n1268), .D(
        w_mult_1_Z[14]), .Y(n1313) );
  ao22d1_hd U1135 ( .A(n1267), .B(w_mult_2_Z[15]), .C(n1268), .D(
        w_mult_1_Z[15]), .Y(n1315) );
  ao22d1_hd U1138 ( .A(n1267), .B(w_mult_2_Z[16]), .C(n1268), .D(
        w_mult_1_Z[16]), .Y(n1317) );
  ao22d1_hd U1141 ( .A(n1267), .B(w_mult_2_Z[17]), .C(n1268), .D(
        w_mult_1_Z[17]), .Y(n1319) );
  scg14d1_hd U1143 ( .A(r_mult_3_A[31]), .B(n1260), .C(n1269), .Y(n77) );
  ao22d1_hd U1145 ( .A(n1267), .B(w_mult_2_Z[18]), .C(n1268), .D(
        w_mult_1_Z[18]), .Y(n1321) );
  ao22d1_hd U1148 ( .A(n1267), .B(w_mult_2_Z[19]), .C(n1268), .D(
        w_mult_1_Z[19]), .Y(n1323) );
  ao22d1_hd U1151 ( .A(n1267), .B(w_mult_2_Z[20]), .C(n1268), .D(
        w_mult_1_Z[20]), .Y(n1325) );
  ao22d1_hd U1154 ( .A(n1267), .B(w_mult_2_Z[21]), .C(n1268), .D(
        w_mult_1_Z[21]), .Y(n1327) );
  ao22d1_hd U1157 ( .A(n1267), .B(w_mult_2_Z[22]), .C(n1268), .D(
        w_mult_1_Z[22]), .Y(n1329) );
  ao22d1_hd U1160 ( .A(n1267), .B(w_mult_2_Z[23]), .C(n1268), .D(
        w_mult_1_Z[23]), .Y(n1331) );
  ao22d1_hd U1163 ( .A(n1267), .B(w_mult_2_Z[24]), .C(n1268), .D(
        w_mult_1_Z[24]), .Y(n1333) );
  ao22d1_hd U1166 ( .A(n1267), .B(w_mult_2_Z[25]), .C(n1268), .D(
        w_mult_1_Z[25]), .Y(n1335) );
  ao22d1_hd U1169 ( .A(n1267), .B(w_mult_2_Z[26]), .C(n1268), .D(
        w_mult_1_Z[26]), .Y(n1337) );
  ao22d1_hd U1172 ( .A(n1267), .B(w_mult_2_Z[27]), .C(n1268), .D(
        w_mult_1_Z[27]), .Y(n1339) );
  ao22d1_hd U1175 ( .A(n507), .B(r_x_data[64]), .C(r_mult_1_B[0]), .D(n9), .Y(
        n1340) );
  ao22d1_hd U1177 ( .A(n1267), .B(w_mult_2_Z[28]), .C(n1268), .D(
        w_mult_1_Z[28]), .Y(n1343) );
  ao22d1_hd U1180 ( .A(n1267), .B(w_mult_2_Z[29]), .C(n1268), .D(
        w_mult_1_Z[29]), .Y(n1345) );
  ao22d1_hd U1183 ( .A(n1267), .B(w_mult_2_Z[30]), .C(n1268), .D(
        w_mult_1_Z[30]), .Y(n1347) );
  scg4d1_hd U1187 ( .A(n1274), .B(r_add_2_B[0]), .C(w_mult_2_Z[0]), .D(n506), 
        .E(r_x_data[96]), .F(n507), .G(n511), .H(w_mult_3_Z[0]), .Y(n755) );
  scg4d1_hd U1188 ( .A(n1274), .B(r_add_2_B[1]), .C(w_mult_2_Z[1]), .D(n506), 
        .E(r_x_data[97]), .F(n508), .G(n511), .H(w_mult_3_Z[1]), .Y(n754) );
  scg4d1_hd U1189 ( .A(n1274), .B(r_add_2_B[2]), .C(w_mult_2_Z[2]), .D(n506), 
        .E(r_x_data[98]), .F(n509), .G(n511), .H(w_mult_3_Z[2]), .Y(n753) );
  scg4d1_hd U1190 ( .A(n1274), .B(r_add_2_B[3]), .C(w_mult_2_Z[3]), .D(n506), 
        .E(r_x_data[99]), .F(n508), .G(n511), .H(w_mult_3_Z[3]), .Y(n752) );
  scg4d1_hd U1191 ( .A(n1274), .B(r_add_2_B[4]), .C(w_mult_2_Z[4]), .D(n506), 
        .E(r_x_data[100]), .F(n2), .G(n511), .H(w_mult_3_Z[4]), .Y(n751) );
  scg4d1_hd U1192 ( .A(n1274), .B(r_add_2_B[5]), .C(w_mult_2_Z[5]), .D(n506), 
        .E(r_x_data[101]), .F(n509), .G(n511), .H(w_mult_3_Z[5]), .Y(n750) );
  ao22d1_hd U1194 ( .A(n507), .B(r_x_data[65]), .C(r_mult_1_B[1]), .D(n9), .Y(
        n1351) );
  scg4d1_hd U1195 ( .A(n1274), .B(r_add_2_B[6]), .C(w_mult_2_Z[6]), .D(n506), 
        .E(r_x_data[102]), .F(n508), .G(n511), .H(w_mult_3_Z[6]), .Y(n749) );
  scg4d1_hd U1196 ( .A(n1274), .B(r_add_2_B[7]), .C(w_mult_2_Z[7]), .D(n506), 
        .E(r_x_data[103]), .F(n507), .G(n511), .H(w_mult_3_Z[7]), .Y(n748) );
  scg4d1_hd U1197 ( .A(n1274), .B(r_add_2_B[8]), .C(w_mult_2_Z[8]), .D(n506), 
        .E(r_x_data[104]), .F(n507), .G(n511), .H(w_mult_3_Z[8]), .Y(n747) );
  scg4d1_hd U1198 ( .A(n1274), .B(r_add_2_B[9]), .C(w_mult_2_Z[9]), .D(n506), 
        .E(r_x_data[105]), .F(n507), .G(n511), .H(w_mult_3_Z[9]), .Y(n746) );
  scg4d1_hd U1199 ( .A(n1274), .B(r_add_2_B[10]), .C(w_mult_2_Z[10]), .D(n506), 
        .E(r_x_data[106]), .F(n508), .G(n511), .H(w_mult_3_Z[10]), .Y(n745) );
  scg4d1_hd U1200 ( .A(n1274), .B(r_add_2_B[11]), .C(w_mult_2_Z[11]), .D(n506), 
        .E(r_x_data[107]), .F(n2), .G(n511), .H(w_mult_3_Z[11]), .Y(n744) );
  scg4d1_hd U1201 ( .A(n1274), .B(r_add_2_B[12]), .C(w_mult_2_Z[12]), .D(n506), 
        .E(r_x_data[108]), .F(n507), .G(n511), .H(w_mult_3_Z[12]), .Y(n743) );
  scg4d1_hd U1202 ( .A(n1274), .B(r_add_2_B[13]), .C(w_mult_2_Z[13]), .D(n506), 
        .E(r_x_data[109]), .F(n509), .G(n511), .H(w_mult_3_Z[13]), .Y(n742) );
  scg4d1_hd U1203 ( .A(n1274), .B(r_add_2_B[14]), .C(w_mult_2_Z[14]), .D(n506), 
        .E(r_x_data[110]), .F(n507), .G(n511), .H(w_mult_3_Z[14]), .Y(n741) );
  scg4d1_hd U1204 ( .A(n1274), .B(r_add_2_B[15]), .C(w_mult_2_Z[15]), .D(n506), 
        .E(r_x_data[111]), .F(n507), .G(n511), .H(w_mult_3_Z[15]), .Y(n740) );
  ao22d1_hd U1206 ( .A(n2), .B(r_x_data[66]), .C(r_mult_1_B[2]), .D(n9), .Y(
        n1352) );
  scg4d1_hd U1207 ( .A(n1274), .B(r_add_2_B[16]), .C(w_mult_2_Z[16]), .D(n506), 
        .E(r_x_data[112]), .F(n508), .G(n511), .H(w_mult_3_Z[16]), .Y(n739) );
  scg4d1_hd U1208 ( .A(n1274), .B(r_add_2_B[17]), .C(w_mult_2_Z[17]), .D(n506), 
        .E(r_x_data[113]), .F(n508), .G(n511), .H(w_mult_3_Z[17]), .Y(n738) );
  scg4d1_hd U1209 ( .A(n1274), .B(r_add_2_B[18]), .C(w_mult_2_Z[18]), .D(n506), 
        .E(r_x_data[114]), .F(n509), .G(n511), .H(w_mult_3_Z[18]), .Y(n737) );
  scg4d1_hd U1210 ( .A(n1274), .B(r_add_2_B[19]), .C(w_mult_2_Z[19]), .D(n506), 
        .E(r_x_data[115]), .F(n510), .G(n511), .H(w_mult_3_Z[19]), .Y(n736) );
  scg4d1_hd U1211 ( .A(n1274), .B(r_add_2_B[20]), .C(w_mult_2_Z[20]), .D(n506), 
        .E(r_x_data[116]), .F(n2), .G(n511), .H(w_mult_3_Z[20]), .Y(n735) );
  scg4d1_hd U1212 ( .A(n1274), .B(r_add_2_B[21]), .C(w_mult_2_Z[21]), .D(n506), 
        .E(r_x_data[117]), .F(n507), .G(n511), .H(w_mult_3_Z[21]), .Y(n734) );
  scg4d1_hd U1213 ( .A(n1274), .B(r_add_2_B[22]), .C(w_mult_2_Z[22]), .D(n506), 
        .E(r_x_data[118]), .F(n510), .G(n511), .H(w_mult_3_Z[22]), .Y(n733) );
  scg4d1_hd U1214 ( .A(n1274), .B(r_add_2_B[23]), .C(w_mult_2_Z[23]), .D(n506), 
        .E(r_x_data[119]), .F(n510), .G(n511), .H(w_mult_3_Z[23]), .Y(n732) );
  scg4d1_hd U1215 ( .A(n1274), .B(r_add_2_B[24]), .C(w_mult_2_Z[24]), .D(n506), 
        .E(r_x_data[120]), .F(n510), .G(n511), .H(w_mult_3_Z[24]), .Y(n731) );
  scg4d1_hd U1216 ( .A(n1274), .B(r_add_2_B[25]), .C(w_mult_2_Z[25]), .D(n506), 
        .E(r_x_data[121]), .F(n510), .G(n511), .H(w_mult_3_Z[25]), .Y(n730) );
  ao22d1_hd U1218 ( .A(n507), .B(r_x_data[67]), .C(r_mult_1_B[3]), .D(n9), .Y(
        n1353) );
  scg4d1_hd U1219 ( .A(n1274), .B(r_add_2_B[26]), .C(w_mult_2_Z[26]), .D(n506), 
        .E(r_x_data[122]), .F(n510), .G(n511), .H(w_mult_3_Z[26]), .Y(n729) );
  scg4d1_hd U1220 ( .A(n1274), .B(r_add_2_B[27]), .C(w_mult_2_Z[27]), .D(n506), 
        .E(r_x_data[123]), .F(n510), .G(n511), .H(w_mult_3_Z[27]), .Y(n728) );
  scg4d1_hd U1221 ( .A(n1274), .B(r_add_2_B[28]), .C(w_mult_2_Z[28]), .D(n506), 
        .E(r_x_data[124]), .F(n510), .G(n511), .H(w_mult_3_Z[28]), .Y(n727) );
  scg4d1_hd U1222 ( .A(n1274), .B(r_add_2_B[29]), .C(w_mult_2_Z[29]), .D(n506), 
        .E(r_x_data[125]), .F(n510), .G(n511), .H(w_mult_3_Z[29]), .Y(n726) );
  scg4d1_hd U1223 ( .A(n1274), .B(r_add_2_B[30]), .C(w_mult_2_Z[30]), .D(n506), 
        .E(r_x_data[126]), .F(n510), .G(n511), .H(w_mult_3_Z[30]), .Y(n725) );
  scg4d1_hd U1226 ( .A(n1358), .B(w_add_2_Z[0]), .C(n1274), .D(r_add_2_A[0]), 
        .E(w_mult_2_Z[0]), .F(n1359), .G(n2), .H(r_x_data[32]), .Y(n723) );
  scg4d1_hd U1227 ( .A(n1358), .B(w_add_2_Z[1]), .C(n1274), .D(r_add_2_A[1]), 
        .E(w_mult_2_Z[1]), .F(n1359), .G(n2), .H(r_x_data[33]), .Y(n722) );
  scg4d1_hd U1228 ( .A(n1358), .B(w_add_2_Z[2]), .C(n1274), .D(r_add_2_A[2]), 
        .E(w_mult_2_Z[2]), .F(n1359), .G(n2), .H(r_x_data[34]), .Y(n721) );
  scg4d1_hd U1229 ( .A(n1358), .B(w_add_2_Z[3]), .C(n1274), .D(r_add_2_A[3]), 
        .E(w_mult_2_Z[3]), .F(n1359), .G(n2), .H(r_x_data[35]), .Y(n720) );
  ao22d1_hd U1231 ( .A(n510), .B(r_x_data[68]), .C(r_mult_1_B[4]), .D(n9), .Y(
        n1360) );
  scg4d1_hd U1232 ( .A(n1358), .B(w_add_2_Z[4]), .C(n1274), .D(r_add_2_A[4]), 
        .E(w_mult_2_Z[4]), .F(n1359), .G(n508), .H(r_x_data[36]), .Y(n719) );
  scg4d1_hd U1233 ( .A(n1358), .B(w_add_2_Z[5]), .C(n1274), .D(r_add_2_A[5]), 
        .E(w_mult_2_Z[5]), .F(n1359), .G(n2), .H(r_x_data[37]), .Y(n718) );
  scg4d1_hd U1234 ( .A(n1358), .B(w_add_2_Z[6]), .C(n1274), .D(r_add_2_A[6]), 
        .E(w_mult_2_Z[6]), .F(n1359), .G(n508), .H(r_x_data[38]), .Y(n717) );
  scg4d1_hd U1235 ( .A(n1358), .B(w_add_2_Z[7]), .C(n1274), .D(r_add_2_A[7]), 
        .E(w_mult_2_Z[7]), .F(n1359), .G(n2), .H(r_x_data[39]), .Y(n716) );
  scg4d1_hd U1236 ( .A(n1358), .B(w_add_2_Z[8]), .C(n1274), .D(r_add_2_A[8]), 
        .E(w_mult_2_Z[8]), .F(n1359), .G(n508), .H(r_x_data[40]), .Y(n715) );
  scg4d1_hd U1237 ( .A(n1358), .B(w_add_2_Z[9]), .C(n1274), .D(r_add_2_A[9]), 
        .E(w_mult_2_Z[9]), .F(n1359), .G(n508), .H(r_x_data[41]), .Y(n714) );
  scg4d1_hd U1238 ( .A(n1358), .B(w_add_2_Z[10]), .C(n1274), .D(r_add_2_A[10]), 
        .E(w_mult_2_Z[10]), .F(n1359), .G(n508), .H(r_x_data[42]), .Y(n713) );
  scg4d1_hd U1239 ( .A(n1358), .B(w_add_2_Z[11]), .C(n1274), .D(r_add_2_A[11]), 
        .E(w_mult_2_Z[11]), .F(n1359), .G(n2), .H(r_x_data[43]), .Y(n712) );
  scg4d1_hd U1240 ( .A(n1358), .B(w_add_2_Z[12]), .C(n1274), .D(r_add_2_A[12]), 
        .E(w_mult_2_Z[12]), .F(n1359), .G(n508), .H(r_x_data[44]), .Y(n711) );
  scg4d1_hd U1241 ( .A(n1358), .B(w_add_2_Z[13]), .C(n1274), .D(r_add_2_A[13]), 
        .E(w_mult_2_Z[13]), .F(n1359), .G(n2), .H(r_x_data[45]), .Y(n710) );
  ao22d1_hd U1243 ( .A(n507), .B(r_x_data[69]), .C(r_mult_1_B[5]), .D(n9), .Y(
        n1361) );
  scg4d1_hd U1244 ( .A(n1358), .B(w_add_2_Z[14]), .C(n1274), .D(r_add_2_A[14]), 
        .E(w_mult_2_Z[14]), .F(n1359), .G(n2), .H(r_x_data[46]), .Y(n709) );
  scg4d1_hd U1245 ( .A(n1358), .B(w_add_2_Z[15]), .C(n1274), .D(r_add_2_A[15]), 
        .E(w_mult_2_Z[15]), .F(n1359), .G(n508), .H(r_x_data[47]), .Y(n708) );
  scg4d1_hd U1246 ( .A(n1358), .B(w_add_2_Z[16]), .C(n1274), .D(r_add_2_A[16]), 
        .E(w_mult_2_Z[16]), .F(n1359), .G(n2), .H(r_x_data[48]), .Y(n707) );
  scg4d1_hd U1247 ( .A(n1358), .B(w_add_2_Z[17]), .C(n1274), .D(r_add_2_A[17]), 
        .E(w_mult_2_Z[17]), .F(n1359), .G(n508), .H(r_x_data[49]), .Y(n706) );
  scg4d1_hd U1248 ( .A(n1358), .B(w_add_2_Z[18]), .C(n1274), .D(r_add_2_A[18]), 
        .E(w_mult_2_Z[18]), .F(n1359), .G(n508), .H(r_x_data[50]), .Y(n705) );
  scg4d1_hd U1249 ( .A(n1358), .B(w_add_2_Z[19]), .C(n1274), .D(r_add_2_A[19]), 
        .E(w_mult_2_Z[19]), .F(n1359), .G(n508), .H(r_x_data[51]), .Y(n704) );
  scg4d1_hd U1250 ( .A(n1358), .B(w_add_2_Z[20]), .C(n1274), .D(r_add_2_A[20]), 
        .E(w_mult_2_Z[20]), .F(n1359), .G(n2), .H(r_x_data[52]), .Y(n703) );
  scg4d1_hd U1251 ( .A(n1358), .B(w_add_2_Z[21]), .C(n1274), .D(r_add_2_A[21]), 
        .E(w_mult_2_Z[21]), .F(n1359), .G(n508), .H(r_x_data[53]), .Y(n702) );
  scg4d1_hd U1252 ( .A(n1358), .B(w_add_2_Z[22]), .C(n1274), .D(r_add_2_A[22]), 
        .E(w_mult_2_Z[22]), .F(n1359), .G(n2), .H(r_x_data[54]), .Y(n701) );
  scg4d1_hd U1253 ( .A(n1358), .B(w_add_2_Z[23]), .C(n1274), .D(r_add_2_A[23]), 
        .E(w_mult_2_Z[23]), .F(n1359), .G(n508), .H(r_x_data[55]), .Y(n700) );
  ao22d1_hd U1255 ( .A(n507), .B(r_x_data[70]), .C(r_mult_1_B[6]), .D(n9), .Y(
        n1362) );
  scg4d1_hd U1256 ( .A(n1358), .B(w_add_2_Z[24]), .C(n1274), .D(r_add_2_A[24]), 
        .E(w_mult_2_Z[24]), .F(n1359), .G(n508), .H(r_x_data[56]), .Y(n699) );
  scg4d1_hd U1257 ( .A(n1358), .B(w_add_2_Z[25]), .C(n1274), .D(r_add_2_A[25]), 
        .E(w_mult_2_Z[25]), .F(n1359), .G(n509), .H(r_x_data[57]), .Y(n698) );
  scg4d1_hd U1258 ( .A(n1358), .B(w_add_2_Z[26]), .C(n1274), .D(r_add_2_A[26]), 
        .E(w_mult_2_Z[26]), .F(n1359), .G(n508), .H(r_x_data[58]), .Y(n697) );
  scg4d1_hd U1259 ( .A(n1358), .B(w_add_2_Z[27]), .C(n1274), .D(r_add_2_A[27]), 
        .E(w_mult_2_Z[27]), .F(n1359), .G(n509), .H(r_x_data[59]), .Y(n696) );
  scg4d1_hd U1260 ( .A(n1358), .B(w_add_2_Z[28]), .C(n1274), .D(r_add_2_A[28]), 
        .E(w_mult_2_Z[28]), .F(n1359), .G(n509), .H(r_x_data[60]), .Y(n695) );
  scg4d1_hd U1261 ( .A(n1358), .B(w_add_2_Z[29]), .C(n1274), .D(r_add_2_A[29]), 
        .E(w_mult_2_Z[29]), .F(n1359), .G(n509), .H(r_x_data[61]), .Y(n694) );
  scg4d1_hd U1262 ( .A(n1358), .B(w_add_2_Z[30]), .C(n1274), .D(r_add_2_A[30]), 
        .E(w_mult_2_Z[30]), .F(n1359), .G(n509), .H(r_x_data[62]), .Y(n693) );
  scg4d1_hd U1263 ( .A(n1358), .B(w_add_2_Z[31]), .C(n1274), .D(r_add_2_A[31]), 
        .E(w_mult_2_Z[31]), .F(n1359), .G(n509), .H(r_x_data[63]), .Y(n692) );
  ao22d1_hd U1272 ( .A(n507), .B(r_x_data[71]), .C(r_mult_1_B[7]), .D(n9), .Y(
        n1368) );
  ao22d1_hd U1284 ( .A(n2), .B(r_x_data[72]), .C(r_mult_1_B[8]), .D(n9), .Y(
        n1369) );
  ao22d1_hd U1296 ( .A(n507), .B(r_x_data[73]), .C(r_mult_1_B[9]), .D(n9), .Y(
        n1370) );
  ao22d1_hd U1315 ( .A(n2), .B(r_x_data[74]), .C(r_mult_1_B[10]), .D(n9), .Y(
        n1376) );
  ao22d1_hd U1317 ( .A(n507), .B(r_x_data[75]), .C(r_mult_1_B[11]), .D(n9), 
        .Y(n1377) );
  ao22d1_hd U1319 ( .A(n2), .B(r_x_data[76]), .C(r_mult_1_B[12]), .D(n9), .Y(
        n1378) );
  ao22d1_hd U1321 ( .A(n507), .B(r_x_data[77]), .C(r_mult_1_B[13]), .D(n9), 
        .Y(n1379) );
  ao22d1_hd U1323 ( .A(n510), .B(r_x_data[78]), .C(r_mult_1_B[14]), .D(n9), 
        .Y(n1380) );
  ao22d1_hd U1325 ( .A(n2), .B(r_x_data[79]), .C(r_mult_1_B[15]), .D(n9), .Y(
        n1381) );
  ao22d1_hd U1327 ( .A(n507), .B(r_x_data[80]), .C(r_mult_1_B[16]), .D(n9), 
        .Y(n1382) );
  ao22d1_hd U1329 ( .A(n510), .B(r_x_data[81]), .C(r_mult_1_B[17]), .D(n9), 
        .Y(n1383) );
  ao22d1_hd U1331 ( .A(n507), .B(r_x_data[82]), .C(r_mult_1_B[18]), .D(n9), 
        .Y(n1384) );
  ao22d1_hd U1333 ( .A(n2), .B(r_x_data[83]), .C(r_mult_1_B[19]), .D(n9), .Y(
        n1385) );
  ao22d1_hd U1335 ( .A(n507), .B(r_x_data[84]), .C(r_mult_1_B[20]), .D(n9), 
        .Y(n1386) );
  ao22d1_hd U1337 ( .A(n2), .B(r_x_data[85]), .C(r_mult_1_B[21]), .D(n9), .Y(
        n1387) );
  ao22d1_hd U1339 ( .A(n507), .B(r_x_data[86]), .C(r_mult_1_B[22]), .D(n9), 
        .Y(n1388) );
  ao22d1_hd U1341 ( .A(n507), .B(r_x_data[87]), .C(r_mult_1_B[23]), .D(n9), 
        .Y(n1389) );
  ao22d1_hd U1343 ( .A(n507), .B(r_x_data[88]), .C(r_mult_1_B[24]), .D(n9), 
        .Y(n1391) );
  ao22d1_hd U1345 ( .A(n507), .B(r_x_data[89]), .C(r_mult_1_B[25]), .D(n9), 
        .Y(n1392) );
  ao22d1_hd U1347 ( .A(w_mult_1_Z[0]), .B(n8), .C(r_mult_1_A[0]), .D(n9), .Y(
        n1393) );
  ao22d1_hd U1349 ( .A(n507), .B(r_y_data[63]), .C(r_mult_3_B[31]), .D(n1260), 
        .Y(n1394) );
  ao22d1_hd U1352 ( .A(n507), .B(r_x_data[90]), .C(r_mult_1_B[26]), .D(n9), 
        .Y(n1395) );
  scg4d1_hd U1353 ( .A(n9), .B(r_mult_2_B[31]), .C(n509), .D(r_y_data[31]), 
        .E(n1396), .F(w_add_2_Z[31]), .G(n8), .H(r_y_data[127]), .Y(n499) );
  scg14d1_hd U1357 ( .A(n1374), .B(r_mult_3_Z_ACK), .C(n1403), .Y(n497) );
  scg15d1_hd U1363 ( .A(n1374), .B(r_mult_1_Z_ACK), .C(n1375), .D(n1403), .Y(
        n493) );
  scg15d1_hd U1364 ( .A(n1374), .B(r_mult_2_Z_ACK), .C(n1375), .D(n1403), .Y(
        n492) );
  scg6d1_hd U1366 ( .A(n1281), .B(r_mult_1_AB_STB), .C(n1406), .Y(n491) );
  scg6d1_hd U1367 ( .A(n1281), .B(r_mult_2_AB_STB), .C(n1406), .Y(n490) );
  ao22d1_hd U1372 ( .A(n507), .B(r_x_data[91]), .C(r_mult_1_B[27]), .D(n9), 
        .Y(n1407) );
  ao22d1_hd U1384 ( .A(n507), .B(r_x_data[92]), .C(r_mult_1_B[28]), .D(n9), 
        .Y(n1408) );
  ao22d1_hd U1396 ( .A(n507), .B(r_x_data[93]), .C(r_mult_1_B[29]), .D(n9), 
        .Y(n1409) );
  ao22d1_hd U1408 ( .A(n507), .B(r_x_data[94]), .C(r_mult_1_B[30]), .D(n9), 
        .Y(n1410) );
  ao22d1_hd U1420 ( .A(n507), .B(r_x_data[95]), .C(r_mult_1_B[31]), .D(n9), 
        .Y(n1411) );
  ao22d1_hd U1443 ( .A(w_mult_1_Z[2]), .B(n8), .C(r_mult_1_A[2]), .D(n9), .Y(
        n1412) );
  ao22d1_hd U1455 ( .A(w_mult_1_Z[3]), .B(n8), .C(r_mult_1_A[3]), .D(n9), .Y(
        n1414) );
  ao22d1_hd U1467 ( .A(w_mult_1_Z[4]), .B(n8), .C(r_mult_1_A[4]), .D(n9), .Y(
        n1415) );
  ao22d1_hd U1479 ( .A(w_mult_1_Z[5]), .B(n8), .C(r_mult_1_A[5]), .D(n9), .Y(
        n1416) );
  ao22d1_hd U1502 ( .A(w_mult_1_Z[7]), .B(n8), .C(r_mult_1_A[7]), .D(n9), .Y(
        n1417) );
  ao22d1_hd U1536 ( .A(w_mult_1_Z[10]), .B(n8), .C(r_mult_1_A[10]), .D(n9), 
        .Y(n1418) );
  ao22d1_hd U1548 ( .A(w_mult_1_Z[11]), .B(n8), .C(r_mult_1_A[11]), .D(n9), 
        .Y(n1419) );
  ao22d1_hd U1571 ( .A(w_mult_1_Z[13]), .B(n8), .C(r_mult_1_A[13]), .D(n9), 
        .Y(n1420) );
  ao22d1_hd U1583 ( .A(w_mult_1_Z[14]), .B(n8), .C(r_mult_1_A[14]), .D(n9), 
        .Y(n1421) );
  ao22d1_hd U1595 ( .A(w_mult_1_Z[15]), .B(n8), .C(r_mult_1_A[15]), .D(n9), 
        .Y(n1422) );
  ao22d1_hd U1618 ( .A(w_mult_1_Z[17]), .B(n8), .C(r_mult_1_A[17]), .D(n9), 
        .Y(n1423) );
  ao22d1_hd U1630 ( .A(w_mult_1_Z[18]), .B(n8), .C(r_mult_1_A[18]), .D(n9), 
        .Y(n1424) );
  ao22d1_hd U1642 ( .A(w_mult_1_Z[19]), .B(n8), .C(r_mult_1_A[19]), .D(n9), 
        .Y(n1425) );
  ao22d1_hd U1665 ( .A(w_mult_1_Z[21]), .B(n8), .C(r_mult_1_A[21]), .D(n9), 
        .Y(n1426) );
  ao22d1_hd U1677 ( .A(w_mult_1_Z[22]), .B(n8), .C(r_mult_1_A[22]), .D(n9), 
        .Y(n1427) );
  ao22d1_hd U1689 ( .A(w_mult_1_Z[23]), .B(n8), .C(r_mult_1_A[23]), .D(n9), 
        .Y(n1428) );
  ao22d1_hd U1701 ( .A(w_mult_1_Z[24]), .B(n8), .C(r_mult_1_A[24]), .D(n9), 
        .Y(n1429) );
  scg4d1_hd U1709 ( .A(n9), .B(r_mult_2_B[0]), .C(w_add_2_Z[0]), .D(n1396), 
        .E(r_y_data[0]), .F(n509), .G(n8), .H(r_y_data[96]), .Y(n202) );
  scg4d1_hd U1710 ( .A(n9), .B(r_mult_2_B[1]), .C(w_add_2_Z[1]), .D(n1396), 
        .E(r_y_data[1]), .F(n509), .G(n8), .H(r_y_data[97]), .Y(n201) );
  scg4d1_hd U1711 ( .A(n1341), .B(r_mult_2_B[2]), .C(w_add_2_Z[2]), .D(n1396), 
        .E(r_y_data[2]), .F(n509), .G(n8), .H(r_y_data[98]), .Y(n200) );
  ao22d1_hd U1713 ( .A(w_mult_1_Z[25]), .B(n8), .C(r_mult_1_A[25]), .D(n9), 
        .Y(n1430) );
  scg4d1_hd U1714 ( .A(n1341), .B(r_mult_2_B[3]), .C(w_add_2_Z[3]), .D(n1396), 
        .E(r_y_data[3]), .F(n509), .G(n8), .H(r_y_data[99]), .Y(n199) );
  scg4d1_hd U1715 ( .A(n1341), .B(r_mult_2_B[4]), .C(w_add_2_Z[4]), .D(n1396), 
        .E(r_y_data[4]), .F(n509), .G(n8), .H(r_y_data[100]), .Y(n198) );
  scg4d1_hd U1716 ( .A(n1341), .B(r_mult_2_B[5]), .C(w_add_2_Z[5]), .D(n1396), 
        .E(r_y_data[5]), .F(n508), .G(n8), .H(r_y_data[101]), .Y(n197) );
  scg4d1_hd U1717 ( .A(n1341), .B(r_mult_2_B[6]), .C(w_add_2_Z[6]), .D(n1396), 
        .E(r_y_data[6]), .F(n509), .G(n8), .H(r_y_data[102]), .Y(n196) );
  scg4d1_hd U1718 ( .A(n1341), .B(r_mult_2_B[7]), .C(w_add_2_Z[7]), .D(n1396), 
        .E(r_y_data[7]), .F(n508), .G(n8), .H(r_y_data[103]), .Y(n195) );
  scg4d1_hd U1719 ( .A(n1341), .B(r_mult_2_B[8]), .C(w_add_2_Z[8]), .D(n1396), 
        .E(r_y_data[8]), .F(n509), .G(n8), .H(r_y_data[104]), .Y(n194) );
  scg4d1_hd U1720 ( .A(n1341), .B(r_mult_2_B[9]), .C(w_add_2_Z[9]), .D(n1396), 
        .E(r_y_data[9]), .F(n508), .G(n8), .H(r_y_data[105]), .Y(n193) );
  scg4d1_hd U1721 ( .A(n1341), .B(r_mult_2_B[10]), .C(w_add_2_Z[10]), .D(n1396), .E(r_y_data[10]), .F(n509), .G(n8), .H(r_y_data[106]), .Y(n192) );
  scg4d1_hd U1722 ( .A(n1341), .B(r_mult_2_B[11]), .C(w_add_2_Z[11]), .D(n1396), .E(r_y_data[11]), .F(n508), .G(n8), .H(r_y_data[107]), .Y(n191) );
  scg4d1_hd U1723 ( .A(n9), .B(r_mult_2_B[12]), .C(w_add_2_Z[12]), .D(n1396), 
        .E(r_y_data[12]), .F(n509), .G(n8), .H(r_y_data[108]), .Y(n190) );
  ao22d1_hd U1725 ( .A(w_mult_1_Z[26]), .B(n8), .C(r_mult_1_A[26]), .D(n9), 
        .Y(n1431) );
  scg4d1_hd U1726 ( .A(n9), .B(r_mult_2_B[13]), .C(w_add_2_Z[13]), .D(n1396), 
        .E(r_y_data[13]), .F(n508), .G(n8), .H(r_y_data[109]), .Y(n189) );
  scg4d1_hd U1727 ( .A(n9), .B(r_mult_2_B[14]), .C(w_add_2_Z[14]), .D(n1396), 
        .E(r_y_data[14]), .F(n509), .G(n8), .H(r_y_data[110]), .Y(n188) );
  scg4d1_hd U1728 ( .A(n9), .B(r_mult_2_B[15]), .C(w_add_2_Z[15]), .D(n1396), 
        .E(r_y_data[15]), .F(n509), .G(n8), .H(r_y_data[111]), .Y(n187) );
  scg4d1_hd U1729 ( .A(n9), .B(r_mult_2_B[16]), .C(w_add_2_Z[16]), .D(n1396), 
        .E(r_y_data[16]), .F(n508), .G(n8), .H(r_y_data[112]), .Y(n186) );
  scg4d1_hd U1730 ( .A(n9), .B(r_mult_2_B[17]), .C(w_add_2_Z[17]), .D(n1396), 
        .E(r_y_data[17]), .F(n508), .G(n8), .H(r_y_data[113]), .Y(n185) );
  scg4d1_hd U1731 ( .A(n9), .B(r_mult_2_B[18]), .C(w_add_2_Z[18]), .D(n1396), 
        .E(r_y_data[18]), .F(n508), .G(n8), .H(r_y_data[114]), .Y(n184) );
  scg4d1_hd U1732 ( .A(n9), .B(r_mult_2_B[19]), .C(w_add_2_Z[19]), .D(n1396), 
        .E(r_y_data[19]), .F(n509), .G(n8), .H(r_y_data[115]), .Y(n183) );
  scg4d1_hd U1733 ( .A(n9), .B(r_mult_2_B[20]), .C(w_add_2_Z[20]), .D(n1396), 
        .E(r_y_data[20]), .F(n510), .G(n8), .H(r_y_data[116]), .Y(n182) );
  scg4d1_hd U1734 ( .A(n9), .B(r_mult_2_B[21]), .C(w_add_2_Z[21]), .D(n1396), 
        .E(r_y_data[21]), .F(n510), .G(n8), .H(r_y_data[117]), .Y(n181) );
  scg4d1_hd U1735 ( .A(n9), .B(r_mult_2_B[22]), .C(w_add_2_Z[22]), .D(n1396), 
        .E(r_y_data[22]), .F(n510), .G(n8), .H(r_y_data[118]), .Y(n180) );
  ao22d1_hd U1737 ( .A(w_mult_1_Z[27]), .B(n8), .C(r_mult_1_A[27]), .D(n9), 
        .Y(n1432) );
  scg4d1_hd U1738 ( .A(n9), .B(r_mult_2_B[23]), .C(w_add_2_Z[23]), .D(n1396), 
        .E(r_y_data[23]), .F(n510), .G(n8), .H(r_y_data[119]), .Y(n179) );
  scg4d1_hd U1739 ( .A(n9), .B(r_mult_2_B[24]), .C(w_add_2_Z[24]), .D(n1396), 
        .E(r_y_data[24]), .F(n510), .G(n8), .H(r_y_data[120]), .Y(n178) );
  scg4d1_hd U1740 ( .A(n9), .B(r_mult_2_B[25]), .C(w_add_2_Z[25]), .D(n1396), 
        .E(r_y_data[25]), .F(n510), .G(n8), .H(r_y_data[121]), .Y(n177) );
  scg4d1_hd U1741 ( .A(n9), .B(r_mult_2_B[26]), .C(w_add_2_Z[26]), .D(n1396), 
        .E(r_y_data[26]), .F(n2), .G(n8), .H(r_y_data[122]), .Y(n176) );
  scg4d1_hd U1742 ( .A(n9), .B(r_mult_2_B[27]), .C(w_add_2_Z[27]), .D(n1396), 
        .E(r_y_data[27]), .F(n507), .G(n8), .H(r_y_data[123]), .Y(n175) );
  scg4d1_hd U1743 ( .A(n9), .B(r_mult_2_B[28]), .C(w_add_2_Z[28]), .D(n1396), 
        .E(r_y_data[28]), .F(n507), .G(n8), .H(r_y_data[124]), .Y(n174) );
  scg4d1_hd U1744 ( .A(n9), .B(r_mult_2_B[29]), .C(w_add_2_Z[29]), .D(n1396), 
        .E(r_y_data[29]), .F(n2), .G(n8), .H(r_y_data[125]), .Y(n173) );
  scg4d1_hd U1745 ( .A(n9), .B(r_mult_2_B[30]), .C(w_add_2_Z[30]), .D(n1396), 
        .E(r_y_data[30]), .F(n509), .G(r_y_data[126]), .H(n8), .Y(n172) );
  scg14d1_hd U1746 ( .A(r_mult_2_A[0]), .B(n9), .C(n1083), .Y(n171) );
  scg14d1_hd U1747 ( .A(r_mult_2_A[1]), .B(n9), .C(n1269), .Y(n170) );
  ao22d1_hd U1749 ( .A(w_mult_1_Z[28]), .B(n8), .C(r_mult_1_A[28]), .D(n9), 
        .Y(n1433) );
  ad2d1_hd U1750 ( .A(r_mult_2_A[2]), .B(n9), .Y(n169) );
  nd2bd1_hd U1751 ( .AN(r_mult_2_A[3]), .B(n1434), .Y(n168) );
  scg14d1_hd U1752 ( .A(r_mult_2_A[4]), .B(n9), .C(n1269), .Y(n167) );
  scg14d1_hd U1753 ( .A(r_mult_2_A[5]), .B(n9), .C(n5), .Y(n166) );
  nd2bd1_hd U1754 ( .AN(r_mult_2_A[6]), .B(n1434), .Y(n165) );
  scg14d1_hd U1755 ( .A(r_mult_2_A[7]), .B(n9), .C(n1403), .Y(n164) );
  nd2bd1_hd U1756 ( .AN(r_mult_2_A[8]), .B(n1434), .Y(n163) );
  scg14d1_hd U1757 ( .A(r_mult_2_A[9]), .B(n9), .C(n1413), .Y(n162) );
  nd2bd1_hd U1758 ( .AN(r_mult_2_A[10]), .B(n1434), .Y(n161) );
  ad2d1_hd U1759 ( .A(r_mult_2_A[11]), .B(n9), .Y(n160) );
  ao22d1_hd U1761 ( .A(w_mult_1_Z[29]), .B(n8), .C(r_mult_1_A[29]), .D(n9), 
        .Y(n1435) );
  scg15d1_hd U1762 ( .A(r_mult_2_A[12]), .B(n9), .C(n1269), .D(n1083), .Y(n159) );
  scg14d1_hd U1763 ( .A(r_mult_2_A[13]), .B(n9), .C(n1269), .Y(n158) );
  scg14d1_hd U1764 ( .A(r_mult_2_A[14]), .B(n9), .C(n1403), .Y(n157) );
  scg14d1_hd U1765 ( .A(r_mult_2_A[15]), .B(n9), .C(n1083), .Y(n156) );
  ad2d1_hd U1766 ( .A(r_mult_2_A[16]), .B(n9), .Y(n155) );
  scg14d1_hd U1767 ( .A(r_mult_2_A[17]), .B(n9), .C(n1083), .Y(n154) );
  scg15d1_hd U1768 ( .A(r_mult_2_A[18]), .B(n9), .C(n1269), .D(n1083), .Y(n153) );
  scg14d1_hd U1769 ( .A(r_mult_2_A[19]), .B(n9), .C(n1403), .Y(n152) );
  scg14d1_hd U1770 ( .A(r_mult_2_A[20]), .B(n9), .C(n1269), .Y(n151) );
  scg14d1_hd U1771 ( .A(r_mult_2_A[21]), .B(n9), .C(n1413), .Y(n150) );
  nd2bd1_hd U1775 ( .AN(r_mult_2_A[22]), .B(n1434), .Y(n149) );
  ad2d1_hd U1776 ( .A(r_mult_2_A[23]), .B(n9), .Y(n148) );
  scg14d1_hd U1777 ( .A(r_mult_2_A[24]), .B(n9), .C(n1083), .Y(n147) );
  nd2bd1_hd U1778 ( .AN(r_mult_2_A[25]), .B(n1434), .Y(n146) );
  nd2bd1_hd U1779 ( .AN(r_mult_2_A[26]), .B(n1434), .Y(n145) );
  nd2bd1_hd U1780 ( .AN(r_mult_2_A[27]), .B(n1434), .Y(n144) );
  nd2bd1_hd U1781 ( .AN(r_mult_2_A[28]), .B(n1434), .Y(n143) );
  nd2bd1_hd U1782 ( .AN(r_mult_2_A[29]), .B(n1434), .Y(n142) );
  ad2d1_hd U1784 ( .A(r_mult_2_A[30]), .B(n9), .Y(n141) );
  scg14d1_hd U1785 ( .A(r_mult_2_A[31]), .B(n9), .C(n1403), .Y(n140) );
  ao22d1_hd U1795 ( .A(n507), .B(r_y_data[32]), .C(r_mult_3_B[0]), .D(n1260), 
        .Y(n1439) );
  ao22d1_hd U1797 ( .A(n507), .B(r_y_data[33]), .C(r_mult_3_B[1]), .D(n1260), 
        .Y(n1440) );
  ao22d1_hd U1799 ( .A(n510), .B(r_y_data[34]), .C(r_mult_3_B[2]), .D(n1260), 
        .Y(n1441) );
  ao22d1_hd U1801 ( .A(n2), .B(r_y_data[35]), .C(r_mult_3_B[3]), .D(n1260), 
        .Y(n1442) );
  ao22d1_hd U1803 ( .A(n507), .B(r_y_data[36]), .C(r_mult_3_B[4]), .D(n1260), 
        .Y(n1443) );
  ao22d1_hd U1805 ( .A(n509), .B(r_y_data[37]), .C(r_mult_3_B[5]), .D(n1260), 
        .Y(n1444) );
  ao22d1_hd U1807 ( .A(n508), .B(r_y_data[38]), .C(r_mult_3_B[6]), .D(n1260), 
        .Y(n1445) );
  ao22d1_hd U1809 ( .A(n507), .B(r_y_data[39]), .C(r_mult_3_B[7]), .D(n1260), 
        .Y(n1446) );
  ao22d1_hd U1811 ( .A(n510), .B(r_y_data[40]), .C(r_mult_3_B[8]), .D(n1260), 
        .Y(n1447) );
  ao22d1_hd U1813 ( .A(n510), .B(r_y_data[41]), .C(r_mult_3_B[9]), .D(n1260), 
        .Y(n1448) );
  ao22d1_hd U1815 ( .A(n510), .B(r_y_data[42]), .C(r_mult_3_B[10]), .D(n1260), 
        .Y(n1449) );
  ao22d1_hd U1817 ( .A(n510), .B(r_y_data[43]), .C(r_mult_3_B[11]), .D(n1260), 
        .Y(n1450) );
  ao22d1_hd U1819 ( .A(n510), .B(r_y_data[44]), .C(r_mult_3_B[12]), .D(n1260), 
        .Y(n1451) );
  ao22d1_hd U1821 ( .A(n510), .B(r_y_data[45]), .C(r_mult_3_B[13]), .D(n1260), 
        .Y(n1452) );
  ao22d1_hd U1823 ( .A(n510), .B(r_y_data[46]), .C(r_mult_3_B[14]), .D(n1260), 
        .Y(n1453) );
  ao22d1_hd U1825 ( .A(n510), .B(r_y_data[47]), .C(r_mult_3_B[15]), .D(n1260), 
        .Y(n1454) );
  ao22d1_hd U1827 ( .A(n510), .B(r_y_data[48]), .C(r_mult_3_B[16]), .D(n1260), 
        .Y(n1455) );
  ao22d1_hd U1829 ( .A(n510), .B(r_y_data[49]), .C(r_mult_3_B[17]), .D(n1260), 
        .Y(n1456) );
  ao22d1_hd U1831 ( .A(n510), .B(r_y_data[50]), .C(r_mult_3_B[18]), .D(n1260), 
        .Y(n1457) );
  ao22d1_hd U1833 ( .A(n508), .B(r_y_data[51]), .C(r_mult_3_B[19]), .D(n1260), 
        .Y(n1458) );
  ao22d1_hd U1835 ( .A(n507), .B(r_y_data[52]), .C(r_mult_3_B[20]), .D(n1260), 
        .Y(n1459) );
  ao22d1_hd U1837 ( .A(n2), .B(r_y_data[53]), .C(r_mult_3_B[21]), .D(n1260), 
        .Y(n1460) );
  ao22d1_hd U1839 ( .A(n510), .B(r_y_data[54]), .C(r_mult_3_B[22]), .D(n1260), 
        .Y(n1461) );
  ao22d1_hd U1841 ( .A(n507), .B(r_y_data[55]), .C(r_mult_3_B[23]), .D(n1260), 
        .Y(n1462) );
  ao22d1_hd U1843 ( .A(n2), .B(r_y_data[56]), .C(r_mult_3_B[24]), .D(n1260), 
        .Y(n1463) );
  ao22d1_hd U1845 ( .A(n507), .B(r_y_data[57]), .C(r_mult_3_B[25]), .D(n1260), 
        .Y(n1464) );
  ao22d1_hd U1847 ( .A(n510), .B(r_y_data[58]), .C(r_mult_3_B[26]), .D(n1260), 
        .Y(n1465) );
  ao22d1_hd U1849 ( .A(n507), .B(r_y_data[59]), .C(r_mult_3_B[27]), .D(n1260), 
        .Y(n1466) );
  ao22d1_hd U1851 ( .A(n2), .B(r_y_data[60]), .C(r_mult_3_B[28]), .D(n1260), 
        .Y(n1467) );
  ao22d1_hd U1853 ( .A(n507), .B(r_y_data[61]), .C(r_mult_3_B[29]), .D(n1260), 
        .Y(n1468) );
  ao22d1_hd U1855 ( .A(n2), .B(r_y_data[62]), .C(r_mult_3_B[30]), .D(n1260), 
        .Y(n1469) );
  scg14d1_hd U1856 ( .A(r_mult_3_A[0]), .B(n1260), .C(n1261), .Y(n108) );
  scg14d1_hd U1857 ( .A(r_mult_3_A[1]), .B(n1260), .C(n1261), .Y(n107) );
  scg14d1_hd U1858 ( .A(r_mult_3_A[2]), .B(n1260), .C(n1269), .Y(n106) );
  nd2bd1_hd U1859 ( .AN(r_mult_3_A[3]), .B(n1262), .Y(n105) );
  nd2bd1_hd U1860 ( .AN(r_mult_3_A[4]), .B(n1262), .Y(n104) );
  nd2bd1_hd U1861 ( .AN(r_mult_3_A[5]), .B(n1262), .Y(n103) );
  scg14d1_hd U1862 ( .A(r_mult_3_A[6]), .B(n1260), .C(n1261), .Y(n102) );
  nd2bd1_hd U1864 ( .AN(r_mult_3_A[7]), .B(n1262), .Y(n101) );
  scg14d1_hd U1867 ( .A(r_mult_3_A[8]), .B(n1260), .C(n1269), .Y(n100) );
  nd4d1_hd U1893 ( .A(w_add_1_Z_STB), .B(w_add_2_Z_STB), .C(w_mult_2_Z_STB), 
        .D(w_mult_1_Z_STB), .Y(n1401) );
  nr2bd1_hd U1892 ( .AN(w_mult_3_Z_STB), .B(n1401), .Y(n1399) );
  ad4d1_hd U1895 ( .A(w_mult_2_AB_ACK), .B(w_mult_3_AB_ACK), .C(
        w_mult_1_AB_ACK), .D(w_add_1_AB_ACK), .Y(n1477) );
  clknd2d1_hd U844 ( .A(n884), .B(n1399), .Y(n517) );
  clknd2d1_hd U845 ( .A(n792), .B(n12), .Y(n882) );
  clknd2d1_hd U846 ( .A(n884), .B(n835), .Y(n832) );
  clknd2d1_hd U847 ( .A(n1375), .B(n1374), .Y(n835) );
  clknd2d1_hd U848 ( .A(n652), .B(n1269), .Y(n520) );
  clknd2d1_hd U849 ( .A(n548), .B(n792), .Y(n522) );
  clknd2d1_hd U850 ( .A(n880), .B(n519), .Y(n521) );
  clknd2d1_hd U851 ( .A(w_add_2_AB_ACK), .B(n1477), .Y(n516) );
  clknd2d1_hd U852 ( .A(n11), .B(n651), .Y(n514) );
  clknd2d1_hd U853 ( .A(n495), .B(n873), .Y(n872) );
  clknd2d1_hd U854 ( .A(n884), .B(n839), .Y(n840) );
  clknd2d4_hd U855 ( .A(n884), .B(n505), .Y(n953) );
  scg6d2_hd U856 ( .A(n12), .B(n511), .C(n1275), .Y(n1358) );
  ad2bd2_hd U857 ( .B(n511), .AN(n12), .Y(n1359) );
  clknd2d1_hd U858 ( .A(n839), .B(n834), .Y(n948) );
  clknd2d4_hd U859 ( .A(n884), .B(n518), .Y(n1261) );
  clknd2d1_hd U860 ( .A(r_counter_1_), .B(n12), .Y(n874) );
  clknd2d1_hd U861 ( .A(w_add_1_Z_STB), .B(w_add_2_Z_STB), .Y(n653) );
  clknd2d1_hd U862 ( .A(n4), .B(i_X_DATA[31]), .Y(n618) );
  clknd2d1_hd U863 ( .A(n4), .B(i_X_DATA[30]), .Y(n619) );
  clknd2d1_hd U864 ( .A(n4), .B(i_X_DATA[29]), .Y(n620) );
  clknd2d1_hd U865 ( .A(n4), .B(i_X_DATA[28]), .Y(n621) );
  clknd2d1_hd U866 ( .A(n4), .B(i_X_DATA[27]), .Y(n622) );
  clknd2d1_hd U867 ( .A(n4), .B(i_X_DATA[26]), .Y(n623) );
  clknd2d1_hd U868 ( .A(n4), .B(i_X_DATA[25]), .Y(n624) );
  clknd2d1_hd U869 ( .A(n4), .B(i_X_DATA[24]), .Y(n625) );
  clknd2d1_hd U870 ( .A(n4), .B(i_X_DATA[23]), .Y(n626) );
  clknd2d1_hd U871 ( .A(n4), .B(i_X_DATA[22]), .Y(n627) );
  clknd2d1_hd U872 ( .A(n4), .B(i_X_DATA[21]), .Y(n628) );
  clknd2d1_hd U873 ( .A(n4), .B(i_X_DATA[20]), .Y(n629) );
  clknd2d1_hd U874 ( .A(n4), .B(i_X_DATA[19]), .Y(n630) );
  clknd2d1_hd U875 ( .A(n4), .B(i_X_DATA[18]), .Y(n631) );
  clknd2d1_hd U876 ( .A(n4), .B(i_X_DATA[17]), .Y(n632) );
  clknd2d1_hd U877 ( .A(n4), .B(i_X_DATA[16]), .Y(n633) );
  clknd2d1_hd U878 ( .A(n4), .B(i_X_DATA[15]), .Y(n634) );
  clknd2d1_hd U879 ( .A(n4), .B(i_X_DATA[14]), .Y(n635) );
  clknd2d1_hd U880 ( .A(n4), .B(i_X_DATA[13]), .Y(n636) );
  clknd2d1_hd U881 ( .A(n4), .B(i_X_DATA[12]), .Y(n637) );
  clknd2d1_hd U882 ( .A(n4), .B(i_X_DATA[11]), .Y(n638) );
  clknd2d1_hd U883 ( .A(n4), .B(i_X_DATA[10]), .Y(n639) );
  clknd2d1_hd U884 ( .A(n4), .B(i_X_DATA[9]), .Y(n640) );
  clknd2d1_hd U885 ( .A(n4), .B(i_X_DATA[8]), .Y(n641) );
  clknd2d1_hd U886 ( .A(n4), .B(i_X_DATA[7]), .Y(n642) );
  clknd2d1_hd U887 ( .A(n4), .B(i_X_DATA[6]), .Y(n643) );
  clknd2d1_hd U888 ( .A(n3), .B(i_X_DATA[5]), .Y(n644) );
  clknd2d1_hd U889 ( .A(n4), .B(i_X_DATA[4]), .Y(n645) );
  clknd2d1_hd U890 ( .A(n3), .B(i_X_DATA[3]), .Y(n646) );
  clknd2d1_hd U891 ( .A(n4), .B(i_X_DATA[2]), .Y(n647) );
  clknd2d1_hd U892 ( .A(n4), .B(i_X_DATA[1]), .Y(n648) );
  clknd2d1_hd U893 ( .A(n3), .B(i_X_DATA[0]), .Y(n649) );
  clknd2d1_hd U894 ( .A(n1413), .B(n1435), .Y(n16) );
  clknd2d1_hd U895 ( .A(n1413), .B(n1433), .Y(n17) );
  clknd2d1_hd U896 ( .A(n1413), .B(n1432), .Y(n18) );
  clknd2d1_hd U897 ( .A(n1413), .B(n1431), .Y(n19) );
  clknd2d1_hd U898 ( .A(n1413), .B(n1430), .Y(n20) );
  clknd2d1_hd U899 ( .A(n1413), .B(n1429), .Y(n21) );
  clknd2d1_hd U900 ( .A(n1428), .B(n1269), .Y(n22) );
  clknd2d1_hd U901 ( .A(n1413), .B(n1427), .Y(n23) );
  clknd2d1_hd U902 ( .A(n1413), .B(n1426), .Y(n24) );
  clknd2d1_hd U903 ( .A(n1425), .B(n1269), .Y(n26) );
  clknd2d1_hd U904 ( .A(n1424), .B(n5), .Y(n27) );
  clknd2d1_hd U905 ( .A(n1423), .B(n5), .Y(n28) );
  clknd2d1_hd U906 ( .A(n1422), .B(n5), .Y(n30) );
  clknd2d1_hd U907 ( .A(n1421), .B(n1269), .Y(n31) );
  clknd2d1_hd U908 ( .A(n1420), .B(n1269), .Y(n32) );
  clknd2d1_hd U909 ( .A(n1419), .B(n5), .Y(n34) );
  clknd2d1_hd U910 ( .A(n1418), .B(n5), .Y(n35) );
  clknd2d1_hd U911 ( .A(n1413), .B(n1417), .Y(n38) );
  clknd2d1_hd U912 ( .A(n1416), .B(n1269), .Y(n40) );
  clknd2d1_hd U913 ( .A(n1415), .B(n5), .Y(n41) );
  clknd2d1_hd U914 ( .A(n1413), .B(n1414), .Y(n42) );
  clknd2d1_hd U915 ( .A(n1412), .B(n5), .Y(n43) );
  clknd2d1_hd U916 ( .A(n1393), .B(n1269), .Y(n502) );
  clknd2d1_hd U917 ( .A(n875), .B(n874), .Y(n877) );
  ivd3_hd U918 ( .A(n1269), .Y(n2) );
  nid6_hd U919 ( .A(n828), .Y(n1) );
  nid8_hd U920 ( .A(n828), .Y(n512) );
  clknd2d3_hd U921 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(n828) );
  ivd6_hd U922 ( .A(n828), .Y(n3) );
  ivd6_hd U923 ( .A(n828), .Y(n4) );
  nid6_hd U924 ( .A(n1341), .Y(n9) );
  ivd3_hd U925 ( .A(n1396), .Y(n5) );
  scg10d1_hd U926 ( .A(n1), .B(r_x_data[16]), .C(r_x_data[48]), .D(n3), .Y(
        n441) );
  scg10d1_hd U927 ( .A(n1), .B(r_x_data[19]), .C(r_x_data[51]), .D(n3), .Y(
        n438) );
  scg10d1_hd U928 ( .A(n1), .B(r_x_data[65]), .C(r_x_data[97]), .D(n3), .Y(
        n392) );
  scg10d1_hd U929 ( .A(n1), .B(r_x_data[18]), .C(r_x_data[50]), .D(n3), .Y(
        n439) );
  scg10d1_hd U930 ( .A(n1), .B(r_x_data[17]), .C(r_x_data[49]), .D(n3), .Y(
        n440) );
  scg10d1_hd U931 ( .A(n1), .B(r_x_data[40]), .C(r_x_data[72]), .D(n3), .Y(
        n417) );
  scg10d1_hd U932 ( .A(n1), .B(r_x_data[39]), .C(r_x_data[71]), .D(n3), .Y(
        n418) );
  scg10d1_hd U933 ( .A(n1), .B(r_x_data[57]), .C(r_x_data[89]), .D(n4), .Y(
        n400) );
  scg10d1_hd U934 ( .A(n1), .B(r_x_data[55]), .C(r_x_data[87]), .D(n3), .Y(
        n402) );
  scg10d1_hd U935 ( .A(n1), .B(r_x_data[9]), .C(r_x_data[41]), .D(n3), .Y(n448) );
  scg10d1_hd U936 ( .A(n1), .B(r_x_data[10]), .C(r_x_data[42]), .D(n3), .Y(
        n447) );
  scg10d1_hd U937 ( .A(n1), .B(r_x_data[37]), .C(r_x_data[69]), .D(n4), .Y(
        n420) );
  scg10d1_hd U938 ( .A(n1), .B(r_x_data[11]), .C(r_x_data[43]), .D(n3), .Y(
        n446) );
  scg10d1_hd U939 ( .A(n1), .B(r_x_data[58]), .C(r_x_data[90]), .D(n3), .Y(
        n399) );
  scg10d1_hd U940 ( .A(n1), .B(r_x_data[12]), .C(r_x_data[44]), .D(n3), .Y(
        n445) );
  scg10d1_hd U941 ( .A(n512), .B(r_x_data[59]), .C(r_x_data[91]), .D(n4), .Y(
        n398) );
  scg10d1_hd U942 ( .A(n1), .B(r_x_data[13]), .C(r_x_data[45]), .D(n3), .Y(
        n444) );
  scg10d1_hd U943 ( .A(n512), .B(r_x_data[60]), .C(r_x_data[92]), .D(n3), .Y(
        n397) );
  scg10d1_hd U944 ( .A(n1), .B(r_x_data[61]), .C(r_x_data[93]), .D(n4), .Y(
        n396) );
  scg10d1_hd U945 ( .A(n1), .B(r_x_data[14]), .C(r_x_data[46]), .D(n3), .Y(
        n443) );
  scg10d1_hd U946 ( .A(n828), .B(r_x_data[66]), .C(r_x_data[98]), .D(n3), .Y(
        n391) );
  scg10d1_hd U947 ( .A(n1), .B(r_x_data[15]), .C(r_x_data[47]), .D(n3), .Y(
        n442) );
  scg10d1_hd U948 ( .A(n1), .B(r_x_data[20]), .C(r_x_data[52]), .D(n3), .Y(
        n437) );
  scg10d1_hd U949 ( .A(n1), .B(r_x_data[21]), .C(r_x_data[53]), .D(n3), .Y(
        n436) );
  scg10d1_hd U950 ( .A(n828), .B(r_x_data[64]), .C(r_x_data[96]), .D(n4), .Y(
        n393) );
  scg10d1_hd U951 ( .A(n1), .B(r_x_data[56]), .C(r_x_data[88]), .D(n3), .Y(
        n401) );
  scg10d1_hd U952 ( .A(n828), .B(r_y_data[95]), .C(r_y_data[127]), .D(n4), .Y(
        n203) );
  scg10d1_hd U953 ( .A(n1), .B(r_x_data[6]), .C(r_x_data[38]), .D(n3), .Y(n451) );
  scg10d1_hd U954 ( .A(n512), .B(r_x_data[44]), .C(r_x_data[76]), .D(n3), .Y(
        n413) );
  scg10d1_hd U955 ( .A(n1), .B(r_x_data[53]), .C(r_x_data[85]), .D(n4), .Y(
        n404) );
  scg10d1_hd U956 ( .A(n1), .B(r_x_data[52]), .C(r_x_data[84]), .D(n3), .Y(
        n405) );
  scg10d1_hd U957 ( .A(n828), .B(r_x_data[46]), .C(r_x_data[78]), .D(n4), .Y(
        n411) );
  scg10d1_hd U958 ( .A(n1), .B(r_x_data[50]), .C(r_x_data[82]), .D(n3), .Y(
        n407) );
  scg10d1_hd U959 ( .A(n1), .B(r_x_data[4]), .C(r_x_data[36]), .D(n3), .Y(n453) );
  scg10d1_hd U960 ( .A(n1), .B(r_x_data[48]), .C(r_x_data[80]), .D(n4), .Y(
        n409) );
  scg10d1_hd U961 ( .A(n1), .B(r_x_data[2]), .C(r_x_data[34]), .D(n3), .Y(n455) );
  scg10d1_hd U962 ( .A(n1), .B(r_x_data[7]), .C(r_x_data[39]), .D(n3), .Y(n450) );
  scg10d1_hd U963 ( .A(n1), .B(r_x_data[42]), .C(r_x_data[74]), .D(n3), .Y(
        n415) );
  scg10d1_hd U964 ( .A(n828), .B(r_x_data[63]), .C(r_x_data[95]), .D(n4), .Y(
        n394) );
  scg10d1_hd U965 ( .A(n1), .B(r_x_data[8]), .C(r_x_data[40]), .D(n3), .Y(n449) );
  scg10d1_hd U966 ( .A(n1), .B(r_x_data[54]), .C(r_x_data[86]), .D(n3), .Y(
        n403) );
  ivd4_hd U967 ( .A(n828), .Y(n6) );
  ivd3_hd U968 ( .A(n504), .Y(n7) );
  nr2d4_hd U969 ( .A(n12), .B(n840), .Y(n1268) );
  nr2d4_hd U970 ( .A(n840), .B(n882), .Y(n1267) );
  ivd4_hd U971 ( .A(n1083), .Y(n8) );
  or2d4_hd U972 ( .A(n883), .B(n522), .Y(n1269) );
  scg10d1_hd U973 ( .A(n1), .B(r_x_data[23]), .C(r_x_data[55]), .D(n4), .Y(
        n434) );
  scg10d1_hd U974 ( .A(n1), .B(r_x_data[22]), .C(r_x_data[54]), .D(n4), .Y(
        n435) );
  scg10d1_hd U975 ( .A(n1), .B(r_x_data[5]), .C(r_x_data[37]), .D(n4), .Y(n452) );
  scg10d1_hd U976 ( .A(n1), .B(r_x_data[3]), .C(r_x_data[35]), .D(n4), .Y(n454) );
  ivd2_hd U977 ( .A(n950), .Y(n504) );
  nd2d4_hd U978 ( .A(n835), .B(n834), .Y(n1274) );
  or2d2_hd U979 ( .A(n1403), .B(n548), .Y(n1083) );
  nr2d4_hd U980 ( .A(n522), .B(n1403), .Y(n1396) );
  scg10d1_hd U981 ( .A(n1), .B(r_x_data[49]), .C(r_x_data[81]), .D(n4), .Y(
        n408) );
  scg10d1_hd U982 ( .A(n1), .B(r_x_data[32]), .C(r_x_data[64]), .D(n4), .Y(
        n425) );
  scg10d1_hd U983 ( .A(n1), .B(r_x_data[36]), .C(r_x_data[68]), .D(n4), .Y(
        n421) );
  nd2d4_hd U984 ( .A(n834), .B(n518), .Y(n1260) );
  scg10d1_hd U985 ( .A(n1), .B(r_x_data[35]), .C(r_x_data[67]), .D(n4), .Y(
        n422) );
  scg10d1_hd U986 ( .A(n1), .B(r_x_data[41]), .C(r_x_data[73]), .D(n4), .Y(
        n416) );
  scg10d1_hd U987 ( .A(n1), .B(r_x_data[33]), .C(r_x_data[65]), .D(n4), .Y(
        n424) );
  scg10d1_hd U988 ( .A(n1), .B(r_x_data[51]), .C(r_x_data[83]), .D(n4), .Y(
        n406) );
  scg10d1_hd U989 ( .A(n512), .B(r_x_data[0]), .C(r_x_data[32]), .D(n3), .Y(
        n457) );
  scg10d1_hd U990 ( .A(n1), .B(r_x_data[34]), .C(r_x_data[66]), .D(n4), .Y(
        n423) );
  scg10d1_hd U991 ( .A(n1), .B(r_x_data[45]), .C(r_x_data[77]), .D(n4), .Y(
        n412) );
  scg10d1_hd U992 ( .A(n1), .B(r_x_data[43]), .C(r_x_data[75]), .D(n4), .Y(
        n414) );
  scg10d1_hd U993 ( .A(n1), .B(r_x_data[38]), .C(r_x_data[70]), .D(n4), .Y(
        n419) );
  scg10d1_hd U994 ( .A(n512), .B(r_y_data[81]), .C(r_y_data[113]), .D(n3), .Y(
        n217) );
  scg10d1_hd U995 ( .A(n512), .B(r_x_data[122]), .C(r_x_data[154]), .D(n6), 
        .Y(n335) );
  scg10d1_hd U996 ( .A(n512), .B(r_y_data[82]), .C(r_y_data[114]), .D(n3), .Y(
        n216) );
  scg10d1_hd U997 ( .A(n512), .B(r_y_data[83]), .C(r_y_data[115]), .D(n3), .Y(
        n215) );
  scg10d1_hd U998 ( .A(n512), .B(r_x_data[121]), .C(r_x_data[153]), .D(n3), 
        .Y(n336) );
  scg10d1_hd U999 ( .A(n512), .B(r_y_data[84]), .C(r_y_data[116]), .D(n3), .Y(
        n214) );
  scg10d1_hd U1000 ( .A(n512), .B(r_y_data[85]), .C(r_y_data[117]), .D(n3), 
        .Y(n213) );
  scg10d1_hd U1001 ( .A(n512), .B(r_x_data[120]), .C(r_x_data[152]), .D(n6), 
        .Y(n337) );
  scg10d1_hd U1002 ( .A(n512), .B(r_y_data[86]), .C(r_y_data[118]), .D(n3), 
        .Y(n212) );
  scg10d1_hd U1003 ( .A(n512), .B(r_x_data[119]), .C(r_x_data[151]), .D(n3), 
        .Y(n338) );
  scg10d1_hd U1004 ( .A(n512), .B(r_x_data[118]), .C(r_x_data[150]), .D(n6), 
        .Y(n339) );
  scg10d1_hd U1005 ( .A(n1), .B(r_x_data[78]), .C(r_x_data[110]), .D(n4), .Y(
        n379) );
  scg10d1_hd U1006 ( .A(n512), .B(r_y_data[87]), .C(r_y_data[119]), .D(n3), 
        .Y(n211) );
  scg10d1_hd U1007 ( .A(n512), .B(r_y_data[88]), .C(r_y_data[120]), .D(n3), 
        .Y(n210) );
  scg10d1_hd U1008 ( .A(n512), .B(r_x_data[117]), .C(r_x_data[149]), .D(n3), 
        .Y(n340) );
  scg10d1_hd U1009 ( .A(n512), .B(r_x_data[116]), .C(r_x_data[148]), .D(n6), 
        .Y(n341) );
  scg10d1_hd U1010 ( .A(n512), .B(r_y_data[89]), .C(r_y_data[121]), .D(n3), 
        .Y(n209) );
  scg10d1_hd U1011 ( .A(n512), .B(r_x_data[114]), .C(r_x_data[146]), .D(n6), 
        .Y(n343) );
  scg10d1_hd U1012 ( .A(n512), .B(r_x_data[113]), .C(r_x_data[145]), .D(n3), 
        .Y(n344) );
  scg10d1_hd U1013 ( .A(n512), .B(r_y_data[90]), .C(r_y_data[122]), .D(n3), 
        .Y(n208) );
  scg10d1_hd U1014 ( .A(n512), .B(r_x_data[112]), .C(r_x_data[144]), .D(n6), 
        .Y(n345) );
  scg10d1_hd U1015 ( .A(n512), .B(r_x_data[111]), .C(r_x_data[143]), .D(n4), 
        .Y(n346) );
  scg10d1_hd U1016 ( .A(n512), .B(r_y_data[91]), .C(r_y_data[123]), .D(n3), 
        .Y(n207) );
  scg10d1_hd U1017 ( .A(n512), .B(r_y_data[92]), .C(r_y_data[124]), .D(n3), 
        .Y(n206) );
  scg10d1_hd U1018 ( .A(n512), .B(r_x_data[110]), .C(r_x_data[142]), .D(n6), 
        .Y(n347) );
  scg10d1_hd U1019 ( .A(n512), .B(r_x_data[109]), .C(r_x_data[141]), .D(n3), 
        .Y(n348) );
  scg10d1_hd U1020 ( .A(n512), .B(r_y_data[93]), .C(r_y_data[125]), .D(n3), 
        .Y(n205) );
  scg10d1_hd U1021 ( .A(n512), .B(r_x_data[108]), .C(r_x_data[140]), .D(n6), 
        .Y(n349) );
  scg10d1_hd U1022 ( .A(n512), .B(r_x_data[107]), .C(r_x_data[139]), .D(n3), 
        .Y(n350) );
  scg10d1_hd U1023 ( .A(n512), .B(r_x_data[106]), .C(r_x_data[138]), .D(n6), 
        .Y(n351) );
  scg10d1_hd U1041 ( .A(n512), .B(r_y_data[94]), .C(r_y_data[126]), .D(n3), 
        .Y(n204) );
  scg10d1_hd U1042 ( .A(n512), .B(r_x_data[105]), .C(r_x_data[137]), .D(n6), 
        .Y(n352) );
  scg10d1_hd U1044 ( .A(n512), .B(r_x_data[104]), .C(r_x_data[136]), .D(n4), 
        .Y(n353) );
  scg10d1_hd U1045 ( .A(n1), .B(r_x_data[30]), .C(r_x_data[62]), .D(n4), .Y(
        n427) );
  scg10d1_hd U1046 ( .A(n512), .B(r_x_data[103]), .C(r_x_data[135]), .D(n6), 
        .Y(n354) );
  scg10d1_hd U1047 ( .A(n1), .B(r_x_data[29]), .C(r_x_data[61]), .D(n4), .Y(
        n428) );
  scg10d1_hd U1048 ( .A(n512), .B(r_y_data[70]), .C(r_y_data[102]), .D(n3), 
        .Y(n228) );
  scg10d1_hd U1049 ( .A(n512), .B(r_y_data[69]), .C(r_y_data[101]), .D(n3), 
        .Y(n229) );
  scg10d1_hd U1050 ( .A(n512), .B(r_y_data[68]), .C(r_y_data[100]), .D(n3), 
        .Y(n230) );
  scg10d1_hd U1052 ( .A(n512), .B(r_y_data[71]), .C(r_y_data[103]), .D(n3), 
        .Y(n227) );
  scg10d1_hd U1053 ( .A(n512), .B(r_y_data[72]), .C(r_y_data[104]), .D(n3), 
        .Y(n226) );
  scg10d1_hd U1054 ( .A(n512), .B(r_y_data[67]), .C(r_y_data[99]), .D(n3), .Y(
        n231) );
  scg10d1_hd U1055 ( .A(n512), .B(r_y_data[66]), .C(r_y_data[98]), .D(n3), .Y(
        n232) );
  scg10d1_hd U1056 ( .A(n512), .B(r_y_data[65]), .C(r_y_data[97]), .D(n3), .Y(
        n233) );
  scg10d1_hd U1057 ( .A(n512), .B(r_y_data[73]), .C(r_y_data[105]), .D(n3), 
        .Y(n225) );
  scg10d1_hd U1058 ( .A(n512), .B(r_x_data[94]), .C(r_x_data[126]), .D(n6), 
        .Y(n363) );
  scg10d1_hd U1059 ( .A(n512), .B(r_y_data[74]), .C(r_y_data[106]), .D(n3), 
        .Y(n224) );
  scg10d1_hd U1060 ( .A(n512), .B(r_x_data[93]), .C(r_x_data[125]), .D(n3), 
        .Y(n364) );
  scg10d1_hd U1061 ( .A(n512), .B(r_y_data[64]), .C(r_y_data[96]), .D(n3), .Y(
        n234) );
  scg10d1_hd U1063 ( .A(n512), .B(r_x_data[127]), .C(r_x_data[159]), .D(n3), 
        .Y(n330) );
  scg10d1_hd U1064 ( .A(n512), .B(r_x_data[92]), .C(r_x_data[124]), .D(n6), 
        .Y(n365) );
  scg10d1_hd U1065 ( .A(n512), .B(r_x_data[126]), .C(r_x_data[158]), .D(n6), 
        .Y(n331) );
  scg10d1_hd U1066 ( .A(n512), .B(r_x_data[91]), .C(r_x_data[123]), .D(n3), 
        .Y(n366) );
  scg10d1_hd U1067 ( .A(n512), .B(r_y_data[75]), .C(r_y_data[107]), .D(n3), 
        .Y(n223) );
  scg10d1_hd U1068 ( .A(n512), .B(r_y_data[76]), .C(r_y_data[108]), .D(n3), 
        .Y(n222) );
  scg10d1_hd U1069 ( .A(n512), .B(r_x_data[90]), .C(r_x_data[122]), .D(n6), 
        .Y(n367) );
  scg10d1_hd U1070 ( .A(n512), .B(r_x_data[89]), .C(r_x_data[121]), .D(n3), 
        .Y(n368) );
  scg10d1_hd U1071 ( .A(n512), .B(r_x_data[88]), .C(r_x_data[120]), .D(n6), 
        .Y(n369) );
  scg10d1_hd U1072 ( .A(n512), .B(r_x_data[87]), .C(r_x_data[119]), .D(n4), 
        .Y(n370) );
  scg10d1_hd U1074 ( .A(n512), .B(r_x_data[125]), .C(r_x_data[157]), .D(n3), 
        .Y(n332) );
  scg10d1_hd U1075 ( .A(n512), .B(r_x_data[86]), .C(r_x_data[118]), .D(n6), 
        .Y(n371) );
  scg10d1_hd U1076 ( .A(n512), .B(r_y_data[77]), .C(r_y_data[109]), .D(n3), 
        .Y(n221) );
  scg10d1_hd U1077 ( .A(n512), .B(r_x_data[85]), .C(r_x_data[117]), .D(n3), 
        .Y(n372) );
  scg10d1_hd U1078 ( .A(n512), .B(r_y_data[78]), .C(r_y_data[110]), .D(n3), 
        .Y(n220) );
  scg10d1_hd U1079 ( .A(n512), .B(r_x_data[124]), .C(r_x_data[156]), .D(n6), 
        .Y(n333) );
  scg10d1_hd U1080 ( .A(n512), .B(r_y_data[79]), .C(r_y_data[111]), .D(n3), 
        .Y(n219) );
  scg10d1_hd U1082 ( .A(n512), .B(r_x_data[123]), .C(r_x_data[155]), .D(n3), 
        .Y(n334) );
  scg10d1_hd U1083 ( .A(n512), .B(r_x_data[84]), .C(r_x_data[116]), .D(n6), 
        .Y(n373) );
  scg10d1_hd U1084 ( .A(n512), .B(r_y_data[80]), .C(r_y_data[112]), .D(n3), 
        .Y(n218) );
  scg10d1_hd U1086 ( .A(n512), .B(r_x_data[83]), .C(r_x_data[115]), .D(n4), 
        .Y(n374) );
  scg10d1_hd U1087 ( .A(n512), .B(r_x_data[82]), .C(r_x_data[114]), .D(n6), 
        .Y(n375) );
  scg10d1_hd U1088 ( .A(n512), .B(r_x_data[115]), .C(r_x_data[147]), .D(n3), 
        .Y(n342) );
  scg10d1_hd U1090 ( .A(n1), .B(r_x_data[25]), .C(r_x_data[57]), .D(n4), .Y(
        n432) );
  scg10d1_hd U1091 ( .A(n1), .B(r_x_data[31]), .C(r_x_data[63]), .D(n4), .Y(
        n426) );
  scg10d1_hd U1093 ( .A(n512), .B(r_x_data[95]), .C(r_x_data[127]), .D(n4), 
        .Y(n362) );
  scg10d1_hd U1094 ( .A(n1), .B(r_x_data[24]), .C(r_x_data[56]), .D(n4), .Y(
        n433) );
  scg10d1_hd U1096 ( .A(n512), .B(r_x_data[102]), .C(r_x_data[134]), .D(n3), 
        .Y(n355) );
  scg10d1_hd U1097 ( .A(n512), .B(r_x_data[101]), .C(r_x_data[133]), .D(n3), 
        .Y(n356) );
  scg10d1_hd U1099 ( .A(n1), .B(r_x_data[28]), .C(r_x_data[60]), .D(n4), .Y(
        n429) );
  scg10d1_hd U1100 ( .A(n512), .B(r_x_data[100]), .C(r_x_data[132]), .D(n6), 
        .Y(n357) );
  scg10d1_hd U1102 ( .A(n512), .B(r_x_data[99]), .C(r_x_data[131]), .D(n3), 
        .Y(n358) );
  scg10d1_hd U1103 ( .A(n1), .B(r_x_data[27]), .C(r_x_data[59]), .D(n4), .Y(
        n430) );
  scg10d1_hd U1105 ( .A(n512), .B(r_x_data[98]), .C(r_x_data[130]), .D(n6), 
        .Y(n359) );
  scg10d1_hd U1106 ( .A(n512), .B(r_x_data[97]), .C(r_x_data[129]), .D(n4), 
        .Y(n360) );
  scg10d1_hd U1108 ( .A(n512), .B(r_x_data[96]), .C(r_x_data[128]), .D(n6), 
        .Y(n361) );
  scg10d1_hd U1109 ( .A(n1), .B(r_x_data[26]), .C(r_x_data[58]), .D(n4), .Y(
        n431) );
  scg10d1_hd U1111 ( .A(n512), .B(r_x_data[79]), .C(r_x_data[111]), .D(n4), 
        .Y(n378) );
  scg10d1_hd U1113 ( .A(n512), .B(r_x_data[80]), .C(r_x_data[112]), .D(n4), 
        .Y(n377) );
  scg10d1_hd U1115 ( .A(n828), .B(r_x_data[73]), .C(r_x_data[105]), .D(n4), 
        .Y(n384) );
  scg10d1_hd U1116 ( .A(n828), .B(r_x_data[74]), .C(r_x_data[106]), .D(n4), 
        .Y(n383) );
  scg10d1_hd U1118 ( .A(n828), .B(r_x_data[72]), .C(r_x_data[104]), .D(n4), 
        .Y(n385) );
  scg10d1_hd U1119 ( .A(n828), .B(r_x_data[75]), .C(r_x_data[107]), .D(n4), 
        .Y(n382) );
  scg10d1_hd U1121 ( .A(n828), .B(r_x_data[76]), .C(r_x_data[108]), .D(n4), 
        .Y(n381) );
  scg10d1_hd U1122 ( .A(n828), .B(r_x_data[71]), .C(r_x_data[103]), .D(n4), 
        .Y(n386) );
  scg10d1_hd U1124 ( .A(n828), .B(r_x_data[70]), .C(r_x_data[102]), .D(n4), 
        .Y(n387) );
  scg10d1_hd U1125 ( .A(n512), .B(r_x_data[81]), .C(r_x_data[113]), .D(n4), 
        .Y(n376) );
  scg10d1_hd U1127 ( .A(n828), .B(r_x_data[77]), .C(r_x_data[109]), .D(n4), 
        .Y(n380) );
  scg10d1_hd U1128 ( .A(n828), .B(r_x_data[69]), .C(r_x_data[101]), .D(n4), 
        .Y(n388) );
  scg10d1_hd U1130 ( .A(n828), .B(r_x_data[68]), .C(r_x_data[100]), .D(n4), 
        .Y(n389) );
  scg10d1_hd U1131 ( .A(n828), .B(r_x_data[67]), .C(r_x_data[99]), .D(n4), .Y(
        n390) );
  scg10d1_hd U1133 ( .A(n828), .B(r_x_data[62]), .C(r_x_data[94]), .D(n4), .Y(
        n395) );
  scg10d1_hd U1134 ( .A(n828), .B(r_x_data[47]), .C(r_x_data[79]), .D(n4), .Y(
        n410) );
  or2d1_hd U1136 ( .A(n517), .B(n833), .Y(n519) );
  scg10d1_hd U1137 ( .A(n512), .B(r_x_data[1]), .C(r_x_data[33]), .D(n4), .Y(
        n456) );
  nr2ad1_hd U1139 ( .A(n884), .B(n515), .Y(n1281) );
  nr2ad1_hd U1140 ( .A(n508), .B(n1396), .Y(n1413) );
  nr2d2_hd U1142 ( .A(r_pstate_0_), .B(n11), .Y(n884) );
  ivd1_hd U1144 ( .A(n521), .Y(n1374) );
  nid2_hd U1146 ( .A(n952), .Y(n505) );
  nid2_hd U1147 ( .A(n1086), .Y(n511) );
  nid2_hd U1149 ( .A(n830), .Y(n13) );
  ivd1_hd U1150 ( .A(n836), .Y(n880) );
  nid2_hd U1152 ( .A(n1275), .Y(n506) );
  oa21d1_hd U1153 ( .A(n883), .B(n882), .C(n881), .Y(n952) );
  ivd1_hd U1155 ( .A(n656), .Y(n883) );
  nd2bd1_hd U1156 ( .AN(n835), .B(n790), .Y(n839) );
  ivd1_hd U1158 ( .A(n792), .Y(n833) );
  nd3bd1_hd U1159 ( .AN(n1401), .B(n884), .C(n654), .Y(n1375) );
  ivd1_hd U1161 ( .A(n831), .Y(n654) );
  nd2d1_hd U1162 ( .A(n521), .B(n834), .Y(n1341) );
  nd2d1_hd U1164 ( .A(n884), .B(n521), .Y(n1403) );
  ao21d1_hd U1165 ( .A(n831), .B(n882), .C(n840), .Y(n830) );
  ivd2_hd U1167 ( .A(n1269), .Y(n509) );
  ivd4_hd U1168 ( .A(n1269), .Y(n507) );
  nid4_hd U1170 ( .A(n948), .Y(n503) );
  oa21d1_hd U1171 ( .A(n516), .B(n522), .C(n836), .Y(n834) );
  ivd2_hd U1173 ( .A(n1269), .Y(n508) );
  nr2d1_hd U1174 ( .A(n880), .B(n516), .Y(n656) );
  nd2bd1_hd U1176 ( .AN(n840), .B(n829), .Y(n950) );
  nr2d1_hd U1178 ( .A(n908), .B(n651), .Y(n836) );
  ivd1_hd U1179 ( .A(r_pstate_0_), .Y(n651) );
  ivd1_hd U1181 ( .A(r_y_data[5]), .Y(n612) );
  ivd1_hd U1182 ( .A(r_y_data[52]), .Y(n566) );
  ivd1_hd U1184 ( .A(r_y_data[20]), .Y(n597) );
  ivd1_hd U1185 ( .A(r_y_data[37]), .Y(n581) );
  ivd1_hd U1186 ( .A(r_y_data[32]), .Y(n586) );
  ivd1_hd U1193 ( .A(r_y_data[27]), .Y(n590) );
  ivd1_hd U1205 ( .A(r_y_data[35]), .Y(n583) );
  ivd1_hd U1217 ( .A(r_y_data[38]), .Y(n580) );
  ivd1_hd U1224 ( .A(r_y_data[34]), .Y(n584) );
  ivd1_hd U1225 ( .A(r_y_data[33]), .Y(n585) );
  ivd1_hd U1230 ( .A(r_y_data[29]), .Y(n588) );
  ivd1_hd U1242 ( .A(r_y_data[28]), .Y(n589) );
  ivd1_hd U1254 ( .A(r_y_data[26]), .Y(n591) );
  ivd1_hd U1264 ( .A(r_y_data[39]), .Y(n579) );
  ivd1_hd U1265 ( .A(r_y_data[57]), .Y(n561) );
  ivd1_hd U1266 ( .A(r_y_data[25]), .Y(n592) );
  ivd1_hd U1267 ( .A(r_y_data[30]), .Y(n587) );
  ivd1_hd U1268 ( .A(r_y_data[36]), .Y(n582) );
  ivd1_hd U1269 ( .A(r_y_data[47]), .Y(n571) );
  ivd1_hd U1270 ( .A(r_y_data[55]), .Y(n563) );
  ivd1_hd U1271 ( .A(r_y_data[23]), .Y(n594) );
  ivd1_hd U1273 ( .A(r_y_data[43]), .Y(n575) );
  ivd1_hd U1274 ( .A(r_y_data[11]), .Y(n606) );
  ivd1_hd U1275 ( .A(r_y_data[41]), .Y(n577) );
  ivd1_hd U1276 ( .A(r_y_data[7]), .Y(n610) );
  ivd1_hd U1277 ( .A(r_y_data[46]), .Y(n572) );
  ivd1_hd U1278 ( .A(r_y_data[14]), .Y(n603) );
  ivd1_hd U1279 ( .A(r_y_data[15]), .Y(n602) );
  ivd1_hd U1280 ( .A(r_y_data[44]), .Y(n574) );
  ivd1_hd U1281 ( .A(r_y_data[6]), .Y(n611) );
  ivd1_hd U1282 ( .A(r_y_data[40]), .Y(n578) );
  ivd1_hd U1283 ( .A(r_y_data[8]), .Y(n609) );
  ivd1_hd U1285 ( .A(r_y_data[4]), .Y(n613) );
  ivd1_hd U1286 ( .A(r_y_data[22]), .Y(n595) );
  ivd1_hd U1287 ( .A(r_y_data[49]), .Y(n569) );
  ivd1_hd U1288 ( .A(r_y_data[17]), .Y(n600) );
  ivd1_hd U1289 ( .A(r_y_data[12]), .Y(n605) );
  ivd1_hd U1290 ( .A(r_y_data[9]), .Y(n608) );
  ivd1_hd U1291 ( .A(r_y_data[2]), .Y(n615) );
  ivd1_hd U1292 ( .A(r_y_data[48]), .Y(n570) );
  ivd1_hd U1293 ( .A(r_y_data[16]), .Y(n601) );
  ivd1_hd U1294 ( .A(r_y_data[50]), .Y(n568) );
  ivd1_hd U1295 ( .A(r_y_data[18]), .Y(n599) );
  ivd1_hd U1297 ( .A(r_y_data[51]), .Y(n567) );
  ivd1_hd U1298 ( .A(r_y_data[19]), .Y(n598) );
  ivd1_hd U1299 ( .A(r_y_data[53]), .Y(n565) );
  ivd1_hd U1300 ( .A(r_y_data[21]), .Y(n596) );
  ivd1_hd U1301 ( .A(r_y_data[42]), .Y(n576) );
  ivd1_hd U1302 ( .A(r_y_data[10]), .Y(n607) );
  ivd1_hd U1303 ( .A(r_y_data[3]), .Y(n614) );
  ivd1_hd U1304 ( .A(r_y_data[56]), .Y(n562) );
  ivd1_hd U1305 ( .A(r_y_data[24]), .Y(n593) );
  ivd1_hd U1306 ( .A(r_y_data[45]), .Y(n573) );
  ivd1_hd U1307 ( .A(r_y_data[13]), .Y(n604) );
  ivd1_hd U1308 ( .A(r_y_data[1]), .Y(n616) );
  ivd1_hd U1309 ( .A(r_y_data[59]), .Y(n559) );
  ivd1_hd U1310 ( .A(r_y_data[0]), .Y(n617) );
  ivd1_hd U1311 ( .A(r_y_data[31]), .Y(n658) );
  ivd1_hd U1312 ( .A(r_y_data[63]), .Y(n555) );
  ivd1_hd U1313 ( .A(r_y_data[62]), .Y(n556) );
  ivd1_hd U1314 ( .A(r_y_data[58]), .Y(n560) );
  ivd1_hd U1316 ( .A(r_y_data[61]), .Y(n557) );
  ivd1_hd U1318 ( .A(r_y_data[54]), .Y(n564) );
  ivd1_hd U1320 ( .A(r_y_data[60]), .Y(n558) );
  nd2d1_hd U1322 ( .A(n521), .B(n520), .Y(n1434) );
  nd2d1_hd U1324 ( .A(n518), .B(n520), .Y(n1262) );
  ivd1_hd U1326 ( .A(r_y_data[79]), .Y(n538) );
  ivd1_hd U1328 ( .A(r_y_data[75]), .Y(n542) );
  ivd1_hd U1330 ( .A(r_y_data[77]), .Y(n540) );
  ivd1_hd U1332 ( .A(r_y_data[81]), .Y(n536) );
  ivd1_hd U1334 ( .A(r_y_data[78]), .Y(n539) );
  ivd1_hd U1336 ( .A(r_y_data[74]), .Y(n543) );
  ivd1_hd U1338 ( .A(r_y_data[76]), .Y(n541) );
  ivd1_hd U1340 ( .A(r_y_data[80]), .Y(n537) );
  ivd1_hd U1342 ( .A(r_y_data[82]), .Y(n535) );
  ivd1_hd U1344 ( .A(r_y_data[73]), .Y(n544) );
  ivd1_hd U1346 ( .A(r_y_data[72]), .Y(n545) );
  ivd1_hd U1348 ( .A(r_y_data[83]), .Y(n534) );
  ivd1_hd U1350 ( .A(r_y_data[93]), .Y(n524) );
  ivd1_hd U1351 ( .A(r_y_data[86]), .Y(n531) );
  ivd1_hd U1354 ( .A(r_y_data[87]), .Y(n530) );
  ivd1_hd U1355 ( .A(r_y_data[88]), .Y(n529) );
  ivd1_hd U1356 ( .A(r_y_data[89]), .Y(n528) );
  ivd1_hd U1358 ( .A(r_y_data[90]), .Y(n527) );
  ivd1_hd U1359 ( .A(r_y_data[91]), .Y(n526) );
  ivd1_hd U1360 ( .A(r_y_data[92]), .Y(n525) );
  ivd1_hd U1361 ( .A(r_y_data[85]), .Y(n532) );
  ivd1_hd U1362 ( .A(r_y_data[84]), .Y(n533) );
  ivd1_hd U1365 ( .A(r_y_data[68]), .Y(n550) );
  ivd1_hd U1368 ( .A(r_y_data[69]), .Y(n549) );
  ivd1_hd U1369 ( .A(r_y_data[65]), .Y(n553) );
  ivd1_hd U1370 ( .A(r_y_data[66]), .Y(n552) );
  ivd1_hd U1371 ( .A(r_y_data[64]), .Y(n554) );
  ivd1_hd U1373 ( .A(r_y_data[67]), .Y(n551) );
  ivd1_hd U1374 ( .A(r_y_data[71]), .Y(n546) );
  ivd1_hd U1375 ( .A(r_y_data[70]), .Y(n547) );
  ivd2_hd U1376 ( .A(n1269), .Y(n510) );
  ivd1_hd U1377 ( .A(o_Y_DATA[1]), .Y(n887) );
  ivd1_hd U1378 ( .A(o_Y_DATA[0]), .Y(n885) );
  ivd1_hd U1379 ( .A(o_Y_DATA[3]), .Y(n891) );
  ivd1_hd U1380 ( .A(o_Y_DATA[4]), .Y(n893) );
  ivd1_hd U1381 ( .A(o_Y_DATA[5]), .Y(n895) );
  ivd1_hd U1382 ( .A(o_Y_DATA[6]), .Y(n897) );
  ivd1_hd U1383 ( .A(o_Y_DATA[2]), .Y(n889) );
  ivd1_hd U1385 ( .A(r_y_data[94]), .Y(n523) );
  ivd1_hd U1386 ( .A(o_Y_DATA[7]), .Y(n899) );
  ivd1_hd U1387 ( .A(o_Y_DATA[30]), .Y(n946) );
  ivd1_hd U1388 ( .A(o_Y_DATA[26]), .Y(n938) );
  ivd1_hd U1389 ( .A(o_Y_DATA[10]), .Y(n905) );
  ivd1_hd U1390 ( .A(o_Y_DATA[29]), .Y(n944) );
  ivd1_hd U1391 ( .A(o_Y_DATA[8]), .Y(n901) );
  ivd1_hd U1392 ( .A(o_Y_DATA[22]), .Y(n930) );
  ivd1_hd U1393 ( .A(o_Y_DATA[9]), .Y(n903) );
  ivd1_hd U1394 ( .A(o_Y_DATA[24]), .Y(n934) );
  ivd1_hd U1395 ( .A(o_Y_DATA[23]), .Y(n932) );
  ivd1_hd U1397 ( .A(o_Y_DATA[25]), .Y(n936) );
  ivd1_hd U1398 ( .A(r_y_data[95]), .Y(n659) );
  oa21d1_hd U1399 ( .A(n517), .B(n522), .C(n880), .Y(n518) );
  ivd1_hd U1400 ( .A(o_Y_DATA[15]), .Y(n916) );
  ivd1_hd U1401 ( .A(o_Y_DATA[16]), .Y(n918) );
  ivd1_hd U1402 ( .A(o_Y_DATA[17]), .Y(n920) );
  ivd1_hd U1403 ( .A(o_Y_DATA[19]), .Y(n924) );
  ivd1_hd U1404 ( .A(o_Y_DATA[18]), .Y(n922) );
  ivd1_hd U1405 ( .A(o_Y_DATA[11]), .Y(n907) );
  ivd1_hd U1406 ( .A(o_Y_DATA[13]), .Y(n912) );
  ivd1_hd U1407 ( .A(o_Y_DATA[31]), .Y(n951) );
  ivd1_hd U1409 ( .A(o_Y_DATA[14]), .Y(n914) );
  ivd1_hd U1410 ( .A(o_Y_DATA[12]), .Y(n910) );
  ivd1_hd U1411 ( .A(o_Y_DATA[28]), .Y(n942) );
  ivd1_hd U1412 ( .A(o_Y_DATA[20]), .Y(n926) );
  ivd1_hd U1413 ( .A(o_Y_DATA[21]), .Y(n928) );
  ivd1_hd U1414 ( .A(o_Y_DATA[27]), .Y(n940) );
  nr2d1_hd U1415 ( .A(n831), .B(n832), .Y(n1275) );
  ivd1_hd U1416 ( .A(w_add_1_Z[21]), .Y(n929) );
  ivd1_hd U1417 ( .A(w_add_1_Z[25]), .Y(n937) );
  ivd1_hd U1418 ( .A(w_add_1_Z[23]), .Y(n933) );
  ivd1_hd U1419 ( .A(w_add_1_Z[26]), .Y(n939) );
  ivd1_hd U1421 ( .A(w_add_1_Z[22]), .Y(n931) );
  ivd1_hd U1422 ( .A(w_add_1_Z[24]), .Y(n935) );
  ivd1_hd U1423 ( .A(w_add_1_Z[27]), .Y(n941) );
  ivd1_hd U1424 ( .A(w_add_1_Z[29]), .Y(n945) );
  ivd1_hd U1425 ( .A(w_add_1_Z[28]), .Y(n943) );
  ivd1_hd U1426 ( .A(w_add_1_Z[30]), .Y(n947) );
  ivd1_hd U1427 ( .A(w_add_1_Z[31]), .Y(n954) );
  ivd1_hd U1428 ( .A(w_add_1_Z[18]), .Y(n923) );
  ivd1_hd U1429 ( .A(w_add_1_Z[14]), .Y(n915) );
  ivd1_hd U1430 ( .A(w_add_1_Z[17]), .Y(n921) );
  ivd1_hd U1431 ( .A(w_add_1_Z[16]), .Y(n919) );
  ivd1_hd U1432 ( .A(w_add_1_Z[15]), .Y(n917) );
  ivd1_hd U1433 ( .A(w_add_1_Z[20]), .Y(n927) );
  ivd1_hd U1434 ( .A(w_add_1_Z[0]), .Y(n886) );
  ivd1_hd U1435 ( .A(w_add_1_Z[1]), .Y(n888) );
  ivd1_hd U1436 ( .A(w_add_1_Z[2]), .Y(n890) );
  ivd1_hd U1437 ( .A(w_add_1_Z[3]), .Y(n892) );
  ivd1_hd U1438 ( .A(w_add_1_Z[4]), .Y(n894) );
  ivd1_hd U1439 ( .A(w_add_1_Z[10]), .Y(n906) );
  ivd1_hd U1440 ( .A(w_add_1_Z[5]), .Y(n896) );
  ivd1_hd U1441 ( .A(w_add_1_Z[6]), .Y(n898) );
  ivd1_hd U1442 ( .A(w_add_1_Z[11]), .Y(n909) );
  ivd1_hd U1444 ( .A(w_add_1_Z[7]), .Y(n900) );
  ivd1_hd U1445 ( .A(w_add_1_Z[13]), .Y(n913) );
  ivd1_hd U1446 ( .A(w_add_1_Z[9]), .Y(n904) );
  ivd1_hd U1447 ( .A(w_add_1_Z[19]), .Y(n925) );
  ivd1_hd U1448 ( .A(w_add_1_Z[12]), .Y(n911) );
  ivd1_hd U1449 ( .A(w_add_1_Z[8]), .Y(n902) );
  nr2d1_hd U1450 ( .A(n10), .B(n874), .Y(n829) );
  nr2d1_hd U1451 ( .A(n10), .B(r_counter_1_), .Y(n792) );
  nd4d1_hd U1452 ( .A(n884), .B(w_add_1_Z_STB), .C(n878), .D(n10), .Y(n881) );
  nr2d1_hd U1453 ( .A(r_counter_1_), .B(n12), .Y(n878) );
  nr2d1_hd U1454 ( .A(n833), .B(n832), .Y(n1086) );
  nd3d1_hd U1456 ( .A(n548), .B(r_counter_1_), .C(n495), .Y(n831) );
  scg2d1_hd U1457 ( .A(w_mult_1_Z[31]), .B(n8), .C(r_mult_1_A[31]), .D(n9), 
        .Y(n14) );
  scg2d1_hd U1458 ( .A(w_mult_1_Z[30]), .B(n8), .C(r_mult_1_A[30]), .D(n9), 
        .Y(n15) );
  scg2d1_hd U1459 ( .A(w_mult_1_Z[20]), .B(n8), .C(r_mult_1_A[20]), .D(n9), 
        .Y(n25) );
  scg2d1_hd U1460 ( .A(w_mult_1_Z[16]), .B(n8), .C(r_mult_1_A[16]), .D(n9), 
        .Y(n29) );
  scg2d1_hd U1461 ( .A(w_mult_1_Z[12]), .B(n8), .C(r_mult_1_A[12]), .D(n9), 
        .Y(n33) );
  scg2d1_hd U1462 ( .A(w_mult_1_Z[9]), .B(n8), .C(r_mult_1_A[9]), .D(n9), .Y(
        n36) );
  scg2d1_hd U1463 ( .A(w_mult_1_Z[8]), .B(n8), .C(r_mult_1_A[8]), .D(n9), .Y(
        n37) );
  scg2d1_hd U1464 ( .A(w_mult_1_Z[6]), .B(n8), .C(r_mult_1_A[6]), .D(n9), .Y(
        n39) );
  scg2d1_hd U1465 ( .A(w_mult_1_Z[1]), .B(n8), .C(r_mult_1_A[1]), .D(n9), .Y(
        n44) );
  nr2d1_hd U1466 ( .A(n880), .B(n833), .Y(N1343) );
  ao211d1_hd U1468 ( .A(o_Y_DATA_VALID), .B(i_Y_ACK), .C(n651), .D(n11), .Y(
        n838) );
  nd4d1_hd U1469 ( .A(n884), .B(n829), .C(w_add_1_Z_STB), .D(w_add_2_Z_STB), 
        .Y(n790) );
  nd4d1_hd U1470 ( .A(n519), .B(n1375), .C(n790), .D(n881), .Y(n879) );
  ao211d1_hd U1471 ( .A(n836), .B(n516), .C(n838), .D(n879), .Y(n513) );
  oa21d1_hd U1472 ( .A(n1), .B(n514), .C(n513), .Y(N1383) );
  nr2d1_hd U1473 ( .A(N23), .B(n514), .Y(N1402) );
  scg20d1_hd U1474 ( .A(n878), .B(n495), .C(n883), .Y(n515) );
  nr2d1_hd U1475 ( .A(n1281), .B(N23), .Y(N1403) );
  ivd1_hd U1476 ( .A(n884), .Y(n652) );
  oa21d1_hd U1477 ( .A(n1261), .B(n523), .C(n1469), .Y(n109) );
  oa21d1_hd U1478 ( .A(n1261), .B(n524), .C(n1468), .Y(n110) );
  oa21d1_hd U1480 ( .A(n1261), .B(n525), .C(n1467), .Y(n111) );
  oa21d1_hd U1481 ( .A(n1261), .B(n526), .C(n1466), .Y(n112) );
  oa21d1_hd U1482 ( .A(n1261), .B(n527), .C(n1465), .Y(n113) );
  oa21d1_hd U1483 ( .A(n1261), .B(n528), .C(n1464), .Y(n114) );
  oa21d1_hd U1484 ( .A(n1261), .B(n529), .C(n1463), .Y(n115) );
  oa21d1_hd U1485 ( .A(n1261), .B(n530), .C(n1462), .Y(n116) );
  oa21d1_hd U1486 ( .A(n1261), .B(n531), .C(n1461), .Y(n117) );
  oa21d1_hd U1487 ( .A(n1261), .B(n532), .C(n1460), .Y(n118) );
  oa21d1_hd U1488 ( .A(n1261), .B(n533), .C(n1459), .Y(n119) );
  oa21d1_hd U1489 ( .A(n1261), .B(n534), .C(n1458), .Y(n120) );
  oa21d1_hd U1490 ( .A(n1261), .B(n535), .C(n1457), .Y(n121) );
  oa21d1_hd U1491 ( .A(n1261), .B(n536), .C(n1456), .Y(n122) );
  oa21d1_hd U1492 ( .A(n1261), .B(n537), .C(n1455), .Y(n123) );
  oa21d1_hd U1493 ( .A(n1261), .B(n538), .C(n1454), .Y(n124) );
  oa21d1_hd U1494 ( .A(n1261), .B(n539), .C(n1453), .Y(n125) );
  oa21d1_hd U1495 ( .A(n1261), .B(n540), .C(n1452), .Y(n126) );
  oa21d1_hd U1496 ( .A(n1261), .B(n541), .C(n1451), .Y(n127) );
  oa21d1_hd U1497 ( .A(n1261), .B(n542), .C(n1450), .Y(n128) );
  oa21d1_hd U1498 ( .A(n1261), .B(n543), .C(n1449), .Y(n129) );
  oa21d1_hd U1499 ( .A(n1261), .B(n544), .C(n1448), .Y(n130) );
  oa21d1_hd U1500 ( .A(n1261), .B(n545), .C(n1447), .Y(n131) );
  oa21d1_hd U1501 ( .A(n1261), .B(n546), .C(n1446), .Y(n132) );
  oa21d1_hd U1503 ( .A(n1261), .B(n547), .C(n1445), .Y(n133) );
  oa21d1_hd U1504 ( .A(n1261), .B(n549), .C(n1444), .Y(n134) );
  oa21d1_hd U1505 ( .A(n1261), .B(n550), .C(n1443), .Y(n135) );
  oa21d1_hd U1506 ( .A(n1261), .B(n551), .C(n1442), .Y(n136) );
  oa21d1_hd U1507 ( .A(n1261), .B(n552), .C(n1441), .Y(n137) );
  oa21d1_hd U1508 ( .A(n1261), .B(n553), .C(n1440), .Y(n138) );
  oa21d1_hd U1509 ( .A(n1261), .B(n554), .C(n1439), .Y(n139) );
  ao22d1_hd U1510 ( .A(n4), .B(n555), .C(n659), .D(n1), .Y(n235) );
  ao22d1_hd U1511 ( .A(n3), .B(n556), .C(n523), .D(n1), .Y(n236) );
  ao22d1_hd U1512 ( .A(n3), .B(n557), .C(n524), .D(n1), .Y(n237) );
  ao22d1_hd U1513 ( .A(n3), .B(n558), .C(n525), .D(n1), .Y(n238) );
  ao22d1_hd U1514 ( .A(n3), .B(n559), .C(n526), .D(n1), .Y(n239) );
  ao22d1_hd U1515 ( .A(n3), .B(n560), .C(n527), .D(n1), .Y(n240) );
  ao22d1_hd U1516 ( .A(n3), .B(n561), .C(n528), .D(n1), .Y(n241) );
  ao22d1_hd U1517 ( .A(n4), .B(n562), .C(n529), .D(n1), .Y(n242) );
  ao22d1_hd U1518 ( .A(n3), .B(n563), .C(n530), .D(n1), .Y(n243) );
  ao22d1_hd U1519 ( .A(n3), .B(n564), .C(n531), .D(n1), .Y(n244) );
  ao22d1_hd U1520 ( .A(n3), .B(n565), .C(n532), .D(n1), .Y(n245) );
  ao22d1_hd U1521 ( .A(n3), .B(n566), .C(n533), .D(n828), .Y(n246) );
  ao22d1_hd U1522 ( .A(n3), .B(n567), .C(n534), .D(n1), .Y(n247) );
  ao22d1_hd U1523 ( .A(n3), .B(n568), .C(n535), .D(n828), .Y(n248) );
  ao22d1_hd U1524 ( .A(n4), .B(n569), .C(n536), .D(n1), .Y(n249) );
  ao22d1_hd U1525 ( .A(n3), .B(n570), .C(n537), .D(n828), .Y(n250) );
  ao22d1_hd U1526 ( .A(n3), .B(n571), .C(n538), .D(n1), .Y(n251) );
  ao22d1_hd U1527 ( .A(n3), .B(n572), .C(n539), .D(n828), .Y(n252) );
  ao22d1_hd U1528 ( .A(n4), .B(n573), .C(n540), .D(n1), .Y(n253) );
  ao22d1_hd U1529 ( .A(n3), .B(n574), .C(n541), .D(n828), .Y(n254) );
  ao22d1_hd U1530 ( .A(n3), .B(n575), .C(n542), .D(n1), .Y(n255) );
  ao22d1_hd U1531 ( .A(n3), .B(n576), .C(n543), .D(n828), .Y(n256) );
  ao22d1_hd U1532 ( .A(n3), .B(n577), .C(n544), .D(n1), .Y(n257) );
  ao22d1_hd U1533 ( .A(n6), .B(n578), .C(n545), .D(n1), .Y(n258) );
  ao22d1_hd U1534 ( .A(n6), .B(n579), .C(n546), .D(n1), .Y(n259) );
  ao22d1_hd U1535 ( .A(n6), .B(n580), .C(n547), .D(n1), .Y(n260) );
  ao22d1_hd U1537 ( .A(n3), .B(n581), .C(n549), .D(n1), .Y(n261) );
  ao22d1_hd U1538 ( .A(n6), .B(n582), .C(n550), .D(n1), .Y(n262) );
  ao22d1_hd U1539 ( .A(n6), .B(n583), .C(n551), .D(n1), .Y(n263) );
  ao22d1_hd U1540 ( .A(n6), .B(n584), .C(n552), .D(n1), .Y(n264) );
  ao22d1_hd U1541 ( .A(n6), .B(n585), .C(n553), .D(n1), .Y(n265) );
  ao22d1_hd U1542 ( .A(n6), .B(n586), .C(n554), .D(n1), .Y(n266) );
  ao22d1_hd U1543 ( .A(n6), .B(n658), .C(n555), .D(n1), .Y(n267) );
  ao22d1_hd U1544 ( .A(n6), .B(n587), .C(n556), .D(n1), .Y(n268) );
  ao22d1_hd U1545 ( .A(n6), .B(n588), .C(n557), .D(n1), .Y(n269) );
  ao22d1_hd U1546 ( .A(n6), .B(n589), .C(n558), .D(n1), .Y(n270) );
  ao22d1_hd U1547 ( .A(n6), .B(n590), .C(n559), .D(n1), .Y(n271) );
  ao22d1_hd U1549 ( .A(n6), .B(n591), .C(n560), .D(n1), .Y(n272) );
  ao22d1_hd U1550 ( .A(n6), .B(n592), .C(n561), .D(n1), .Y(n273) );
  ao22d1_hd U1551 ( .A(n6), .B(n593), .C(n562), .D(n1), .Y(n274) );
  ao22d1_hd U1552 ( .A(n6), .B(n594), .C(n563), .D(n1), .Y(n275) );
  ao22d1_hd U1553 ( .A(n6), .B(n595), .C(n564), .D(n1), .Y(n276) );
  ao22d1_hd U1554 ( .A(n6), .B(n596), .C(n565), .D(n1), .Y(n277) );
  ao22d1_hd U1555 ( .A(n6), .B(n597), .C(n566), .D(n828), .Y(n278) );
  ao22d1_hd U1556 ( .A(n6), .B(n598), .C(n567), .D(n1), .Y(n279) );
  ao22d1_hd U1557 ( .A(n6), .B(n599), .C(n568), .D(n1), .Y(n280) );
  ao22d1_hd U1558 ( .A(n6), .B(n600), .C(n569), .D(n1), .Y(n281) );
  ao22d1_hd U1559 ( .A(n6), .B(n601), .C(n570), .D(n512), .Y(n282) );
  ao22d1_hd U1560 ( .A(n6), .B(n602), .C(n571), .D(n1), .Y(n283) );
  ao22d1_hd U1561 ( .A(n6), .B(n603), .C(n572), .D(n1), .Y(n284) );
  ao22d1_hd U1562 ( .A(n6), .B(n604), .C(n573), .D(n1), .Y(n285) );
  ao22d1_hd U1563 ( .A(n6), .B(n605), .C(n574), .D(n1), .Y(n286) );
  ao22d1_hd U1564 ( .A(n6), .B(n606), .C(n575), .D(n1), .Y(n287) );
  ao22d1_hd U1565 ( .A(n6), .B(n607), .C(n576), .D(n1), .Y(n288) );
  ao22d1_hd U1566 ( .A(n6), .B(n608), .C(n577), .D(n1), .Y(n289) );
  ao22d1_hd U1567 ( .A(n6), .B(n609), .C(n578), .D(n1), .Y(n290) );
  ao22d1_hd U1568 ( .A(n4), .B(n610), .C(n579), .D(n512), .Y(n291) );
  ao22d1_hd U1569 ( .A(n4), .B(n611), .C(n580), .D(n512), .Y(n292) );
  ao22d1_hd U1570 ( .A(n4), .B(n612), .C(n581), .D(n512), .Y(n293) );
  ao22d1_hd U1572 ( .A(n4), .B(n613), .C(n582), .D(n512), .Y(n294) );
  ao22d1_hd U1573 ( .A(n4), .B(n614), .C(n583), .D(n512), .Y(n295) );
  ao22d1_hd U1574 ( .A(n4), .B(n615), .C(n584), .D(n512), .Y(n296) );
  ao22d1_hd U1575 ( .A(n4), .B(n616), .C(n585), .D(n512), .Y(n297) );
  ao22d1_hd U1576 ( .A(n4), .B(n617), .C(n586), .D(n512), .Y(n298) );
  ao22d1_hd U1577 ( .A(n6), .B(n946), .C(n587), .D(n1), .Y(n299) );
  ao22d1_hd U1578 ( .A(n3), .B(n944), .C(n588), .D(n512), .Y(n300) );
  ao22d1_hd U1579 ( .A(n4), .B(n942), .C(n589), .D(n512), .Y(n301) );
  ao22d1_hd U1580 ( .A(n3), .B(n940), .C(n590), .D(n512), .Y(n302) );
  ao22d1_hd U1581 ( .A(n4), .B(n938), .C(n591), .D(n512), .Y(n303) );
  ao22d1_hd U1582 ( .A(n3), .B(n936), .C(n592), .D(n512), .Y(n304) );
  ao22d1_hd U1584 ( .A(n4), .B(n934), .C(n593), .D(n512), .Y(n305) );
  ao22d1_hd U1585 ( .A(n3), .B(n932), .C(n594), .D(n512), .Y(n306) );
  ao22d1_hd U1586 ( .A(n4), .B(n930), .C(n595), .D(n512), .Y(n307) );
  ao22d1_hd U1587 ( .A(n3), .B(n928), .C(n596), .D(n512), .Y(n308) );
  ao22d1_hd U1588 ( .A(n4), .B(n926), .C(n597), .D(n828), .Y(n309) );
  ao22d1_hd U1589 ( .A(n3), .B(n924), .C(n598), .D(n1), .Y(n310) );
  ao22d1_hd U1590 ( .A(n3), .B(n922), .C(n599), .D(n1), .Y(n311) );
  ao22d1_hd U1591 ( .A(n3), .B(n920), .C(n600), .D(n828), .Y(n312) );
  ao22d1_hd U1592 ( .A(n4), .B(n918), .C(n601), .D(n1), .Y(n313) );
  ao22d1_hd U1593 ( .A(n3), .B(n916), .C(n602), .D(n1), .Y(n314) );
  ao22d1_hd U1594 ( .A(n4), .B(n914), .C(n603), .D(n828), .Y(n315) );
  ao22d1_hd U1596 ( .A(n3), .B(n912), .C(n604), .D(n1), .Y(n316) );
  ao22d1_hd U1597 ( .A(n4), .B(n910), .C(n605), .D(n1), .Y(n317) );
  ao22d1_hd U1598 ( .A(n3), .B(n907), .C(n606), .D(n828), .Y(n318) );
  ao22d1_hd U1599 ( .A(n4), .B(n905), .C(n607), .D(n1), .Y(n319) );
  ao22d1_hd U1600 ( .A(n3), .B(n903), .C(n608), .D(n1), .Y(n320) );
  ao22d1_hd U1601 ( .A(n4), .B(n901), .C(n609), .D(n828), .Y(n321) );
  ao22d1_hd U1602 ( .A(n3), .B(n899), .C(n610), .D(n1), .Y(n322) );
  ao22d1_hd U1603 ( .A(n4), .B(n897), .C(n611), .D(n1), .Y(n323) );
  ao22d1_hd U1604 ( .A(n3), .B(n895), .C(n612), .D(n828), .Y(n324) );
  ao22d1_hd U1605 ( .A(n4), .B(n893), .C(n613), .D(n1), .Y(n325) );
  ao22d1_hd U1606 ( .A(n3), .B(n891), .C(n614), .D(n1), .Y(n326) );
  ao22d1_hd U1607 ( .A(n4), .B(n889), .C(n615), .D(n512), .Y(n327) );
  ao22d1_hd U1608 ( .A(n3), .B(n887), .C(n616), .D(n1), .Y(n328) );
  ao22d1_hd U1609 ( .A(n4), .B(n885), .C(n617), .D(n1), .Y(n329) );
  oa21d1_hd U1610 ( .A(n954), .B(n5), .C(n1411), .Y(n45) );
  scg14d1_hd U1611 ( .A(r_x_data[31]), .B(n512), .C(n618), .Y(n458) );
  scg14d1_hd U1612 ( .A(r_x_data[30]), .B(n512), .C(n619), .Y(n459) );
  oa21d1_hd U1613 ( .A(n947), .B(n5), .C(n1410), .Y(n46) );
  scg14d1_hd U1614 ( .A(r_x_data[29]), .B(n512), .C(n620), .Y(n460) );
  scg14d1_hd U1615 ( .A(r_x_data[28]), .B(n512), .C(n621), .Y(n461) );
  scg14d1_hd U1616 ( .A(r_x_data[27]), .B(n512), .C(n622), .Y(n462) );
  scg14d1_hd U1617 ( .A(r_x_data[26]), .B(n512), .C(n623), .Y(n463) );
  scg14d1_hd U1619 ( .A(r_x_data[25]), .B(n512), .C(n624), .Y(n464) );
  scg14d1_hd U1620 ( .A(r_x_data[24]), .B(n512), .C(n625), .Y(n465) );
  scg14d1_hd U1621 ( .A(r_x_data[23]), .B(n512), .C(n626), .Y(n466) );
  scg14d1_hd U1622 ( .A(r_x_data[22]), .B(n512), .C(n627), .Y(n467) );
  scg14d1_hd U1623 ( .A(r_x_data[21]), .B(n512), .C(n628), .Y(n468) );
  scg14d1_hd U1624 ( .A(r_x_data[20]), .B(n512), .C(n629), .Y(n469) );
  oa211d1_hd U1625 ( .A(n5), .B(n945), .C(n1409), .D(n1083), .Y(n47) );
  scg14d1_hd U1626 ( .A(r_x_data[19]), .B(n512), .C(n630), .Y(n470) );
  scg14d1_hd U1627 ( .A(r_x_data[18]), .B(n512), .C(n631), .Y(n471) );
  scg14d1_hd U1628 ( .A(r_x_data[17]), .B(n512), .C(n632), .Y(n472) );
  scg14d1_hd U1629 ( .A(r_x_data[16]), .B(n512), .C(n633), .Y(n473) );
  scg14d1_hd U1631 ( .A(r_x_data[15]), .B(n512), .C(n634), .Y(n474) );
  scg14d1_hd U1632 ( .A(r_x_data[14]), .B(n512), .C(n635), .Y(n475) );
  scg14d1_hd U1633 ( .A(r_x_data[13]), .B(n512), .C(n636), .Y(n476) );
  scg14d1_hd U1634 ( .A(r_x_data[12]), .B(n512), .C(n637), .Y(n477) );
  scg14d1_hd U1635 ( .A(r_x_data[11]), .B(n512), .C(n638), .Y(n478) );
  scg14d1_hd U1636 ( .A(r_x_data[10]), .B(n512), .C(n639), .Y(n479) );
  oa211d1_hd U1637 ( .A(n5), .B(n943), .C(n1408), .D(n1083), .Y(n48) );
  scg14d1_hd U1638 ( .A(r_x_data[9]), .B(n512), .C(n640), .Y(n480) );
  scg14d1_hd U1639 ( .A(r_x_data[8]), .B(n512), .C(n641), .Y(n481) );
  scg14d1_hd U1640 ( .A(r_x_data[7]), .B(n512), .C(n642), .Y(n482) );
  scg14d1_hd U1641 ( .A(r_x_data[6]), .B(n512), .C(n643), .Y(n483) );
  scg14d1_hd U1643 ( .A(r_x_data[5]), .B(n512), .C(n644), .Y(n484) );
  scg14d1_hd U1644 ( .A(r_x_data[4]), .B(n512), .C(n645), .Y(n485) );
  scg14d1_hd U1645 ( .A(r_x_data[3]), .B(n512), .C(n646), .Y(n486) );
  scg14d1_hd U1646 ( .A(r_x_data[2]), .B(n512), .C(n647), .Y(n487) );
  scg14d1_hd U1647 ( .A(r_x_data[1]), .B(n512), .C(n648), .Y(n488) );
  scg14d1_hd U1648 ( .A(r_x_data[0]), .B(n512), .C(n649), .Y(n489) );
  oa211d1_hd U1649 ( .A(n5), .B(n941), .C(n1407), .D(n1083), .Y(n49) );
  ivd1_hd U1650 ( .A(N1343), .Y(n650) );
  nr2d1_hd U1651 ( .A(n1281), .B(n880), .Y(n873) );
  oa22d1_hd U1652 ( .A(n1281), .B(n650), .C(n12), .D(n872), .Y(n1406) );
  oa21d1_hd U1653 ( .A(n11), .B(n879), .C(n651), .Y(n876) );
  nr3d1_hd U1654 ( .A(n10), .B(n652), .C(n876), .Y(n875) );
  ao22d1_hd U1655 ( .A(n875), .B(n829), .C(n10), .D(n876), .Y(n494) );
  ao22d1_hd U1656 ( .A(n548), .B(n875), .C(n876), .D(n12), .Y(n496) );
  ao211d1_hd U1657 ( .A(n1401), .B(n654), .C(n10), .D(n653), .Y(n655) );
  oa21d1_hd U1658 ( .A(r_counter_1_), .B(n1399), .C(n655), .Y(n657) );
  ao211d1_hd U1659 ( .A(n884), .B(n657), .C(n838), .D(n656), .Y(n498) );
  oa211d1_hd U1660 ( .A(n5), .B(n939), .C(n1395), .D(n1083), .Y(n50) );
  ao22d1_hd U1661 ( .A(n4), .B(n951), .C(n658), .D(n1), .Y(n500) );
  oa21d1_hd U1662 ( .A(n1261), .B(n659), .C(n1394), .Y(n501) );
  oa211d1_hd U1663 ( .A(n5), .B(n937), .C(n1392), .D(n1083), .Y(n51) );
  oa211d1_hd U1664 ( .A(n5), .B(n935), .C(n1391), .D(n1083), .Y(n52) );
  oa211d1_hd U1666 ( .A(n5), .B(n933), .C(n1389), .D(n1083), .Y(n53) );
  oa21d1_hd U1667 ( .A(n931), .B(n5), .C(n1388), .Y(n54) );
  oa21d1_hd U1668 ( .A(n929), .B(n5), .C(n1387), .Y(n55) );
  oa21d1_hd U1669 ( .A(n927), .B(n5), .C(n1386), .Y(n56) );
  oa21d1_hd U1670 ( .A(n925), .B(n5), .C(n1385), .Y(n57) );
  oa21d1_hd U1671 ( .A(n923), .B(n5), .C(n1384), .Y(n58) );
  oa21d1_hd U1672 ( .A(n921), .B(n5), .C(n1383), .Y(n59) );
  oa21d1_hd U1673 ( .A(n919), .B(n5), .C(n1382), .Y(n60) );
  oa21d1_hd U1674 ( .A(n917), .B(n5), .C(n1381), .Y(n61) );
  oa21d1_hd U1675 ( .A(n915), .B(n5), .C(n1380), .Y(n62) );
  oa21d1_hd U1676 ( .A(n913), .B(n5), .C(n1379), .Y(n63) );
  oa21d1_hd U1678 ( .A(n911), .B(n5), .C(n1378), .Y(n64) );
  oa21d1_hd U1679 ( .A(n909), .B(n5), .C(n1377), .Y(n65) );
  oa21d1_hd U1680 ( .A(n906), .B(n5), .C(n1376), .Y(n66) );
  scg4d1_hd U1681 ( .A(n503), .B(r_add_1_B[31]), .C(n13), .D(w_add_1_Z[31]), 
        .E(w_add_2_Z[31]), .F(n504), .G(n2), .H(r_x_data[159]), .Y(n660) );
  scg4d1_hd U1682 ( .A(n13), .B(w_add_1_Z[30]), .C(n503), .D(r_add_1_B[30]), 
        .E(w_add_2_Z[30]), .F(n504), .G(r_x_data[158]), .H(n2), .Y(n661) );
  scg4d1_hd U1683 ( .A(n13), .B(w_add_1_Z[29]), .C(n503), .D(r_add_1_B[29]), 
        .E(w_add_2_Z[29]), .F(n504), .G(r_x_data[157]), .H(n507), .Y(n662) );
  scg4d1_hd U1684 ( .A(n13), .B(w_add_1_Z[28]), .C(n503), .D(r_add_1_B[28]), 
        .E(w_add_2_Z[28]), .F(n504), .G(r_x_data[156]), .H(n2), .Y(n663) );
  scg4d1_hd U1685 ( .A(n13), .B(w_add_1_Z[27]), .C(n503), .D(r_add_1_B[27]), 
        .E(w_add_2_Z[27]), .F(n504), .G(r_x_data[155]), .H(n2), .Y(n664) );
  scg4d1_hd U1686 ( .A(n13), .B(w_add_1_Z[26]), .C(n503), .D(r_add_1_B[26]), 
        .E(w_add_2_Z[26]), .F(n504), .G(r_x_data[154]), .H(n2), .Y(n665) );
  scg4d1_hd U1687 ( .A(n13), .B(w_add_1_Z[25]), .C(n503), .D(r_add_1_B[25]), 
        .E(w_add_2_Z[25]), .F(n504), .G(r_x_data[153]), .H(n507), .Y(n666) );
  scg4d1_hd U1688 ( .A(n13), .B(w_add_1_Z[24]), .C(n503), .D(r_add_1_B[24]), 
        .E(w_add_2_Z[24]), .F(n504), .G(r_x_data[152]), .H(n2), .Y(n667) );
  scg4d1_hd U1690 ( .A(n13), .B(w_add_1_Z[23]), .C(n503), .D(r_add_1_B[23]), 
        .E(w_add_2_Z[23]), .F(n504), .G(r_x_data[151]), .H(n507), .Y(n668) );
  scg4d1_hd U1691 ( .A(n13), .B(w_add_1_Z[22]), .C(n503), .D(r_add_1_B[22]), 
        .E(w_add_2_Z[22]), .F(n504), .G(r_x_data[150]), .H(n2), .Y(n669) );
  oa21d1_hd U1692 ( .A(n904), .B(n5), .C(n1370), .Y(n67) );
  scg4d1_hd U1693 ( .A(n830), .B(w_add_1_Z[21]), .C(n503), .D(r_add_1_B[21]), 
        .E(w_add_2_Z[21]), .F(n504), .G(r_x_data[149]), .H(n507), .Y(n670) );
  scg4d1_hd U1694 ( .A(n830), .B(w_add_1_Z[20]), .C(n503), .D(r_add_1_B[20]), 
        .E(w_add_2_Z[20]), .F(n504), .G(r_x_data[148]), .H(n507), .Y(n671) );
  scg4d1_hd U1695 ( .A(n830), .B(w_add_1_Z[19]), .C(n503), .D(r_add_1_B[19]), 
        .E(w_add_2_Z[19]), .F(n504), .G(r_x_data[147]), .H(n507), .Y(n672) );
  scg4d1_hd U1696 ( .A(n830), .B(w_add_1_Z[18]), .C(n503), .D(r_add_1_B[18]), 
        .E(w_add_2_Z[18]), .F(n504), .G(r_x_data[146]), .H(n507), .Y(n673) );
  scg4d1_hd U1697 ( .A(n830), .B(w_add_1_Z[17]), .C(n503), .D(r_add_1_B[17]), 
        .E(w_add_2_Z[17]), .F(n504), .G(r_x_data[145]), .H(n507), .Y(n674) );
  scg4d1_hd U1698 ( .A(n13), .B(w_add_1_Z[16]), .C(n503), .D(r_add_1_B[16]), 
        .E(w_add_2_Z[16]), .F(n504), .G(r_x_data[144]), .H(n507), .Y(n675) );
  scg4d1_hd U1699 ( .A(n13), .B(w_add_1_Z[15]), .C(n503), .D(r_add_1_B[15]), 
        .E(w_add_2_Z[15]), .F(n504), .G(r_x_data[143]), .H(n2), .Y(n676) );
  scg4d1_hd U1700 ( .A(n13), .B(w_add_1_Z[14]), .C(n503), .D(r_add_1_B[14]), 
        .E(w_add_2_Z[14]), .F(n504), .G(r_x_data[142]), .H(n507), .Y(n677) );
  scg4d1_hd U1702 ( .A(n13), .B(w_add_1_Z[13]), .C(n503), .D(r_add_1_B[13]), 
        .E(w_add_2_Z[13]), .F(n504), .G(r_x_data[141]), .H(n507), .Y(n678) );
  scg4d1_hd U1703 ( .A(n13), .B(w_add_1_Z[12]), .C(n503), .D(r_add_1_B[12]), 
        .E(w_add_2_Z[12]), .F(n504), .G(r_x_data[140]), .H(n2), .Y(n679) );
  oa21d1_hd U1704 ( .A(n902), .B(n5), .C(n1369), .Y(n68) );
  scg4d1_hd U1705 ( .A(n13), .B(w_add_1_Z[11]), .C(n503), .D(r_add_1_B[11]), 
        .E(w_add_2_Z[11]), .F(n504), .G(r_x_data[139]), .H(n2), .Y(n680) );
  scg4d1_hd U1706 ( .A(n13), .B(w_add_1_Z[10]), .C(n503), .D(r_add_1_B[10]), 
        .E(w_add_2_Z[10]), .F(n504), .G(r_x_data[138]), .H(n507), .Y(n681) );
  scg4d1_hd U1707 ( .A(n13), .B(w_add_1_Z[9]), .C(n503), .D(r_add_1_B[9]), .E(
        w_add_2_Z[9]), .F(n504), .G(r_x_data[137]), .H(n2), .Y(n682) );
  scg4d1_hd U1708 ( .A(n13), .B(w_add_1_Z[8]), .C(n503), .D(r_add_1_B[8]), .E(
        w_add_2_Z[8]), .F(n504), .G(r_x_data[136]), .H(n507), .Y(n683) );
  scg4d1_hd U1712 ( .A(n13), .B(w_add_1_Z[7]), .C(n503), .D(r_add_1_B[7]), .E(
        w_add_2_Z[7]), .F(n504), .G(r_x_data[135]), .H(n2), .Y(n684) );
  scg4d1_hd U1724 ( .A(n13), .B(w_add_1_Z[6]), .C(n503), .D(r_add_1_B[6]), .E(
        w_add_2_Z[6]), .F(n504), .G(r_x_data[134]), .H(n507), .Y(n685) );
  scg4d1_hd U1736 ( .A(n13), .B(w_add_1_Z[5]), .C(n503), .D(r_add_1_B[5]), .E(
        w_add_2_Z[5]), .F(n504), .G(r_x_data[133]), .H(n2), .Y(n686) );
  scg4d1_hd U1748 ( .A(n13), .B(w_add_1_Z[4]), .C(n503), .D(r_add_1_B[4]), .E(
        w_add_2_Z[4]), .F(n504), .G(r_x_data[132]), .H(n507), .Y(n687) );
  scg4d1_hd U1760 ( .A(n13), .B(w_add_1_Z[3]), .C(n503), .D(r_add_1_B[3]), .E(
        w_add_2_Z[3]), .F(n504), .G(r_x_data[131]), .H(n2), .Y(n688) );
  scg4d1_hd U1772 ( .A(n13), .B(w_add_1_Z[2]), .C(n503), .D(r_add_1_B[2]), .E(
        w_add_2_Z[2]), .F(n504), .G(r_x_data[130]), .H(n2), .Y(n689) );
  oa21d1_hd U1773 ( .A(n900), .B(n5), .C(n1368), .Y(n69) );
  scg4d1_hd U1774 ( .A(n13), .B(w_add_1_Z[1]), .C(n503), .D(r_add_1_B[1]), .E(
        w_add_2_Z[1]), .F(n504), .G(r_x_data[129]), .H(n2), .Y(n690) );
  scg4d1_hd U1783 ( .A(n13), .B(w_add_1_Z[0]), .C(n503), .D(r_add_1_B[0]), .E(
        w_add_2_Z[0]), .F(n504), .G(r_x_data[128]), .H(n2), .Y(n691) );
  oa21d1_hd U1786 ( .A(n898), .B(n5), .C(n1362), .Y(n70) );
  oa21d1_hd U1787 ( .A(n896), .B(n5), .C(n1361), .Y(n71) );
  oa21d1_hd U1788 ( .A(n894), .B(n5), .C(n1360), .Y(n72) );
  oa21d1_hd U1789 ( .A(n836), .B(n884), .C(o_Y_DATA_VALID), .Y(n837) );
  nd2bd1_hd U1790 ( .AN(n838), .B(n837), .Y(n724) );
  oa21d1_hd U1791 ( .A(n892), .B(n5), .C(n1353), .Y(n73) );
  oa21d1_hd U1792 ( .A(n890), .B(n5), .C(n1352), .Y(n74) );
  oa21d1_hd U1793 ( .A(n888), .B(n5), .C(n1351), .Y(n75) );
  scg16d1_hd U1794 ( .A(r_add_2_Z_ACK), .B(n839), .C(n840), .Y(n756) );
  ao22d1_hd U1796 ( .A(n507), .B(r_x_data[30]), .C(r_add_1_A[30]), .D(n503), 
        .Y(n841) );
  oa211d1_hd U1798 ( .A(n7), .B(n947), .C(n1347), .D(n841), .Y(n757) );
  ao22d1_hd U1800 ( .A(n507), .B(r_x_data[29]), .C(r_add_1_A[29]), .D(n503), 
        .Y(n842) );
  oa211d1_hd U1802 ( .A(n7), .B(n945), .C(n1345), .D(n842), .Y(n758) );
  ao22d1_hd U1804 ( .A(n509), .B(r_x_data[28]), .C(r_add_1_A[28]), .D(n503), 
        .Y(n843) );
  oa211d1_hd U1806 ( .A(n7), .B(n943), .C(n1343), .D(n843), .Y(n759) );
  oa21d1_hd U1808 ( .A(n886), .B(n5), .C(n1340), .Y(n76) );
  ao22d1_hd U1810 ( .A(n508), .B(r_x_data[27]), .C(r_add_1_A[27]), .D(n503), 
        .Y(n844) );
  oa211d1_hd U1812 ( .A(n7), .B(n941), .C(n1339), .D(n844), .Y(n760) );
  ao22d1_hd U1814 ( .A(n509), .B(r_x_data[26]), .C(r_add_1_A[26]), .D(n503), 
        .Y(n845) );
  oa211d1_hd U1816 ( .A(n7), .B(n939), .C(n1337), .D(n845), .Y(n761) );
  ao22d1_hd U1818 ( .A(n508), .B(r_x_data[25]), .C(r_add_1_A[25]), .D(n503), 
        .Y(n846) );
  oa211d1_hd U1820 ( .A(n7), .B(n937), .C(n1335), .D(n846), .Y(n762) );
  ao22d1_hd U1822 ( .A(n507), .B(r_x_data[24]), .C(r_add_1_A[24]), .D(n503), 
        .Y(n847) );
  oa211d1_hd U1824 ( .A(n7), .B(n935), .C(n1333), .D(n847), .Y(n763) );
  ao22d1_hd U1826 ( .A(n2), .B(r_x_data[23]), .C(r_add_1_A[23]), .D(n503), .Y(
        n848) );
  oa211d1_hd U1828 ( .A(n7), .B(n933), .C(n1331), .D(n848), .Y(n764) );
  ao22d1_hd U1830 ( .A(n509), .B(r_x_data[22]), .C(r_add_1_A[22]), .D(n503), 
        .Y(n849) );
  oa211d1_hd U1832 ( .A(n7), .B(n931), .C(n1329), .D(n849), .Y(n765) );
  ao22d1_hd U1834 ( .A(n508), .B(r_x_data[21]), .C(r_add_1_A[21]), .D(n503), 
        .Y(n850) );
  oa211d1_hd U1836 ( .A(n7), .B(n929), .C(n1327), .D(n850), .Y(n766) );
  ao22d1_hd U1838 ( .A(n507), .B(r_x_data[20]), .C(r_add_1_A[20]), .D(n503), 
        .Y(n851) );
  oa211d1_hd U1840 ( .A(n7), .B(n927), .C(n1325), .D(n851), .Y(n767) );
  ao22d1_hd U1842 ( .A(n507), .B(r_x_data[19]), .C(r_add_1_A[19]), .D(n503), 
        .Y(n852) );
  oa211d1_hd U1844 ( .A(n7), .B(n925), .C(n1323), .D(n852), .Y(n768) );
  ao22d1_hd U1846 ( .A(n2), .B(r_x_data[18]), .C(r_add_1_A[18]), .D(n503), .Y(
        n853) );
  oa211d1_hd U1848 ( .A(n7), .B(n923), .C(n1321), .D(n853), .Y(n769) );
  ao22d1_hd U1850 ( .A(n507), .B(r_x_data[17]), .C(r_add_1_A[17]), .D(n503), 
        .Y(n854) );
  oa211d1_hd U1852 ( .A(n7), .B(n921), .C(n1319), .D(n854), .Y(n770) );
  ao22d1_hd U1854 ( .A(n507), .B(r_x_data[16]), .C(r_add_1_A[16]), .D(n503), 
        .Y(n855) );
  oa211d1_hd U1863 ( .A(n7), .B(n919), .C(n1317), .D(n855), .Y(n771) );
  ao22d1_hd U1865 ( .A(n508), .B(r_x_data[15]), .C(r_add_1_A[15]), .D(n503), 
        .Y(n856) );
  oa211d1_hd U1866 ( .A(n7), .B(n917), .C(n1315), .D(n856), .Y(n772) );
  ao22d1_hd U1868 ( .A(n2), .B(r_x_data[14]), .C(r_add_1_A[14]), .D(n503), .Y(
        n857) );
  oa211d1_hd U1869 ( .A(n7), .B(n915), .C(n1313), .D(n857), .Y(n773) );
  ao22d1_hd U1870 ( .A(n507), .B(r_x_data[13]), .C(r_add_1_A[13]), .D(n503), 
        .Y(n858) );
  oa211d1_hd U1871 ( .A(n7), .B(n913), .C(n1311), .D(n858), .Y(n774) );
  ao22d1_hd U1872 ( .A(n507), .B(r_x_data[12]), .C(r_add_1_A[12]), .D(n503), 
        .Y(n859) );
  oa211d1_hd U1873 ( .A(n7), .B(n911), .C(n1309), .D(n859), .Y(n775) );
  ao22d1_hd U1874 ( .A(n2), .B(r_x_data[11]), .C(r_add_1_A[11]), .D(n503), .Y(
        n860) );
  oa211d1_hd U1875 ( .A(n7), .B(n909), .C(n1307), .D(n860), .Y(n776) );
  ao22d1_hd U1876 ( .A(n507), .B(r_x_data[10]), .C(r_add_1_A[10]), .D(n503), 
        .Y(n861) );
  oa211d1_hd U1877 ( .A(n7), .B(n906), .C(n1305), .D(n861), .Y(n777) );
  ao22d1_hd U1878 ( .A(n509), .B(r_x_data[9]), .C(r_add_1_A[9]), .D(n503), .Y(
        n862) );
  oa211d1_hd U1879 ( .A(n7), .B(n904), .C(n1303), .D(n862), .Y(n778) );
  ao22d1_hd U1880 ( .A(n508), .B(r_x_data[8]), .C(r_add_1_A[8]), .D(n503), .Y(
        n863) );
  oa211d1_hd U1881 ( .A(n7), .B(n902), .C(n1301), .D(n863), .Y(n779) );
  ao22d1_hd U1882 ( .A(n507), .B(r_x_data[7]), .C(r_add_1_A[7]), .D(n503), .Y(
        n864) );
  oa211d1_hd U1883 ( .A(n7), .B(n900), .C(n1299), .D(n864), .Y(n780) );
  ao22d1_hd U1884 ( .A(n510), .B(r_x_data[6]), .C(r_add_1_A[6]), .D(n503), .Y(
        n865) );
  oa211d1_hd U1885 ( .A(n7), .B(n898), .C(n1297), .D(n865), .Y(n781) );
  ao22d1_hd U1886 ( .A(n2), .B(r_x_data[5]), .C(r_add_1_A[5]), .D(n503), .Y(
        n866) );
  oa211d1_hd U1887 ( .A(n7), .B(n896), .C(n1295), .D(n866), .Y(n782) );
  ao22d1_hd U1888 ( .A(n509), .B(r_x_data[4]), .C(r_add_1_A[4]), .D(n503), .Y(
        n867) );
  oa211d1_hd U1889 ( .A(n7), .B(n894), .C(n1293), .D(n867), .Y(n783) );
  ao22d1_hd U1890 ( .A(n509), .B(r_x_data[3]), .C(r_add_1_A[3]), .D(n503), .Y(
        n868) );
  oa211d1_hd U1891 ( .A(n7), .B(n892), .C(n1291), .D(n868), .Y(n784) );
  ao22d1_hd U1894 ( .A(n509), .B(r_x_data[2]), .C(r_add_1_A[2]), .D(n503), .Y(
        n869) );
  oa211d1_hd U1896 ( .A(n7), .B(n890), .C(n1289), .D(n869), .Y(n785) );
  ao22d1_hd U1897 ( .A(n509), .B(r_x_data[1]), .C(r_add_1_A[1]), .D(n503), .Y(
        n870) );
  oa211d1_hd U1898 ( .A(n7), .B(n888), .C(n1287), .D(n870), .Y(n786) );
  ao22d1_hd U1899 ( .A(n509), .B(r_x_data[0]), .C(r_add_1_A[0]), .D(n503), .Y(
        n871) );
  oa211d1_hd U1900 ( .A(n7), .B(n886), .C(n1285), .D(n871), .Y(n787) );
  scg14d1_hd U1901 ( .A(n1281), .B(r_add_2_AB_STB), .C(n872), .Y(n788) );
  scg6d1_hd U1902 ( .A(n1281), .B(r_add_1_AB_STB), .C(n873), .Y(n789) );
  oa22ad1_hd U1903 ( .A(n878), .B(n877), .C(n876), .D(r_counter_1_), .Y(n791)
         );
  scg6d1_hd U1904 ( .A(r_add_1_Z_ACK), .B(n880), .C(n879), .Y(n793) );
  oa22d1_hd U1905 ( .A(n886), .B(n953), .C(n505), .D(n885), .Y(n795) );
  oa22d1_hd U1906 ( .A(n888), .B(n953), .C(n505), .D(n887), .Y(n796) );
  oa22d1_hd U1907 ( .A(n890), .B(n953), .C(n505), .D(n889), .Y(n797) );
  oa22d1_hd U1908 ( .A(n892), .B(n953), .C(n505), .D(n891), .Y(n798) );
  oa22d1_hd U1909 ( .A(n894), .B(n953), .C(n505), .D(n893), .Y(n799) );
  oa22d1_hd U1910 ( .A(n896), .B(n953), .C(n505), .D(n895), .Y(n800) );
  oa22d1_hd U1911 ( .A(n898), .B(n953), .C(n505), .D(n897), .Y(n801) );
  oa22d1_hd U1912 ( .A(n900), .B(n953), .C(n505), .D(n899), .Y(n802) );
  oa22d1_hd U1913 ( .A(n902), .B(n953), .C(n505), .D(n901), .Y(n803) );
  oa22d1_hd U1914 ( .A(n904), .B(n953), .C(n505), .D(n903), .Y(n804) );
  oa22d1_hd U1915 ( .A(n906), .B(n953), .C(n505), .D(n905), .Y(n805) );
  oa22d1_hd U1916 ( .A(n909), .B(n953), .C(n505), .D(n907), .Y(n806) );
  oa22d1_hd U1917 ( .A(n911), .B(n953), .C(n505), .D(n910), .Y(n807) );
  oa22d1_hd U1918 ( .A(n913), .B(n953), .C(n505), .D(n912), .Y(n808) );
  oa22d1_hd U1919 ( .A(n915), .B(n953), .C(n505), .D(n914), .Y(n809) );
  oa22d1_hd U1920 ( .A(n917), .B(n953), .C(n952), .D(n916), .Y(n810) );
  oa22d1_hd U1921 ( .A(n919), .B(n953), .C(n952), .D(n918), .Y(n811) );
  oa22d1_hd U1922 ( .A(n921), .B(n953), .C(n952), .D(n920), .Y(n812) );
  oa22d1_hd U1923 ( .A(n923), .B(n953), .C(n952), .D(n922), .Y(n813) );
  oa22d1_hd U1924 ( .A(n925), .B(n953), .C(n952), .D(n924), .Y(n814) );
  oa22d1_hd U1925 ( .A(n927), .B(n953), .C(n505), .D(n926), .Y(n815) );
  oa22d1_hd U1926 ( .A(n929), .B(n953), .C(n505), .D(n928), .Y(n816) );
  oa22d1_hd U1927 ( .A(n931), .B(n953), .C(n505), .D(n930), .Y(n817) );
  oa22d1_hd U1928 ( .A(n933), .B(n953), .C(n505), .D(n932), .Y(n818) );
  oa22d1_hd U1929 ( .A(n935), .B(n953), .C(n505), .D(n934), .Y(n819) );
  oa22d1_hd U1930 ( .A(n937), .B(n953), .C(n505), .D(n936), .Y(n820) );
  oa22d1_hd U1931 ( .A(n939), .B(n953), .C(n505), .D(n938), .Y(n821) );
  oa22d1_hd U1932 ( .A(n941), .B(n953), .C(n505), .D(n940), .Y(n822) );
  oa22d1_hd U1933 ( .A(n943), .B(n953), .C(n505), .D(n942), .Y(n823) );
  oa22d1_hd U1934 ( .A(n945), .B(n953), .C(n505), .D(n944), .Y(n824) );
  oa22d1_hd U1935 ( .A(n947), .B(n953), .C(n505), .D(n946), .Y(n825) );
  ao22d1_hd U1936 ( .A(n509), .B(r_x_data[31]), .C(r_add_1_A[31]), .D(n503), 
        .Y(n949) );
  oa211d1_hd U1937 ( .A(n954), .B(n7), .C(n1266), .D(n949), .Y(n826) );
  oa22d1_hd U1938 ( .A(n954), .B(n953), .C(n505), .D(n951), .Y(n827) );
endmodule


module float_adder_2 ( i_A, i_B, i_AB_STB, o_AB_ACK, o_Z, o_Z_STB, i_Z_ACK, 
        i_CLK, i_RST );
  input [31:0] i_A;
  input [31:0] i_B;
  output [31:0] o_Z;
  input i_AB_STB, i_Z_ACK, i_CLK, i_RST;
  output o_AB_ACK, o_Z_STB;
  wire   N41, a_s, b_s, guard, round_bit, sticky, z_s, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, C91_DATA2_1, C91_DATA2_2, C91_DATA2_3, C91_DATA2_4,
         C91_DATA2_5, C91_DATA2_6, C91_DATA2_7, C91_DATA2_8, n1, n2, n27, n265,
         n266, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n509, C2_Z_26, C2_Z_25, C2_Z_24, C2_Z_23,
         C2_Z_22, C2_Z_21, C2_Z_20, C2_Z_19, C2_Z_18, C2_Z_17, C2_Z_16,
         C2_Z_15, C2_Z_14, C2_Z_13, C2_Z_12, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_43J4_124_6938_n58, DP_OP_43J4_124_6938_n57,
         DP_OP_43J4_124_6938_n56, DP_OP_43J4_124_6938_n55,
         DP_OP_43J4_124_6938_n54, DP_OP_43J4_124_6938_n53,
         DP_OP_43J4_124_6938_n52, DP_OP_43J4_124_6938_n51,
         DP_OP_43J4_124_6938_n50, DP_OP_43J4_124_6938_n49,
         DP_OP_43J4_124_6938_n48, DP_OP_43J4_124_6938_n47,
         DP_OP_43J4_124_6938_n46, DP_OP_43J4_124_6938_n45,
         DP_OP_43J4_124_6938_n44, DP_OP_43J4_124_6938_n43,
         DP_OP_43J4_124_6938_n42, DP_OP_43J4_124_6938_n41,
         DP_OP_43J4_124_6938_n40, DP_OP_43J4_124_6938_n39,
         DP_OP_43J4_124_6938_n38, DP_OP_43J4_124_6938_n37,
         DP_OP_43J4_124_6938_n36, DP_OP_43J4_124_6938_n35,
         DP_OP_43J4_124_6938_n34, DP_OP_43J4_124_6938_n33,
         DP_OP_43J4_124_6938_n32, DP_OP_43J4_124_6938_n27,
         DP_OP_43J4_124_6938_n26, DP_OP_43J4_124_6938_n25,
         DP_OP_43J4_124_6938_n24, DP_OP_43J4_124_6938_n23,
         DP_OP_43J4_124_6938_n22, DP_OP_43J4_124_6938_n21,
         DP_OP_43J4_124_6938_n20, DP_OP_43J4_124_6938_n19,
         DP_OP_43J4_124_6938_n18, DP_OP_43J4_124_6938_n17,
         DP_OP_43J4_124_6938_n16, DP_OP_43J4_124_6938_n15,
         DP_OP_43J4_124_6938_n14, DP_OP_43J4_124_6938_n13,
         DP_OP_43J4_124_6938_n12, DP_OP_43J4_124_6938_n11,
         DP_OP_43J4_124_6938_n10, DP_OP_43J4_124_6938_n9,
         DP_OP_43J4_124_6938_n8, DP_OP_43J4_124_6938_n7,
         DP_OP_43J4_124_6938_n6, DP_OP_43J4_124_6938_n5,
         DP_OP_43J4_124_6938_n4, DP_OP_43J4_124_6938_n3,
         DP_OP_43J4_124_6938_n2, DP_OP_43J4_124_6938_n1,
         DP_OP_154J4_137_6175_n9, DP_OP_154J4_137_6175_n8,
         DP_OP_154J4_137_6175_n7, DP_OP_154J4_137_6175_n6,
         DP_OP_154J4_137_6175_n5, DP_OP_154J4_137_6175_n4,
         DP_OP_154J4_137_6175_n3, DP_OP_154J4_137_6175_n2, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
  wire   [3:0] state;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [9:0] a_e;
  wire   [26:0] a_m;
  wire   [9:0] b_e;
  wire   [26:0] b_m;
  wire   [27:0] sum;
  wire   [9:0] z_e;
  wire   [23:0] z_m;
  wire   [31:0] z;

  ivd1_hd U485 ( .A(i_RST), .Y(N41) );
  fad1_hd DP_OP_154J4_137_6175_U10 ( .A(n2266), .B(z_e[1]), .CI(z_e[0]), .CO(
        DP_OP_154J4_137_6175_n9), .S(C91_DATA2_1) );
  fad1_hd DP_OP_154J4_137_6175_U9 ( .A(n2266), .B(z_e[2]), .CI(
        DP_OP_154J4_137_6175_n9), .CO(DP_OP_154J4_137_6175_n8), .S(C91_DATA2_2) );
  fad1_hd DP_OP_154J4_137_6175_U8 ( .A(n2266), .B(z_e[3]), .CI(
        DP_OP_154J4_137_6175_n8), .CO(DP_OP_154J4_137_6175_n7), .S(C91_DATA2_3) );
  fad1_hd DP_OP_154J4_137_6175_U7 ( .A(n2266), .B(z_e[4]), .CI(
        DP_OP_154J4_137_6175_n7), .CO(DP_OP_154J4_137_6175_n6), .S(C91_DATA2_4) );
  fad1_hd DP_OP_154J4_137_6175_U6 ( .A(n2266), .B(z_e[5]), .CI(
        DP_OP_154J4_137_6175_n6), .CO(DP_OP_154J4_137_6175_n5), .S(C91_DATA2_5) );
  fad1_hd DP_OP_154J4_137_6175_U5 ( .A(n2266), .B(z_e[6]), .CI(
        DP_OP_154J4_137_6175_n5), .CO(DP_OP_154J4_137_6175_n4), .S(C91_DATA2_6) );
  fad1_hd DP_OP_154J4_137_6175_U4 ( .A(n2266), .B(z_e[7]), .CI(
        DP_OP_154J4_137_6175_n4), .CO(DP_OP_154J4_137_6175_n3), .S(C91_DATA2_7) );
  fad1_hd DP_OP_154J4_137_6175_U3 ( .A(n2266), .B(z_e[8]), .CI(
        DP_OP_154J4_137_6175_n3), .CO(DP_OP_154J4_137_6175_n2), .S(C91_DATA2_8) );
  fd1qd1_hd z_e_reg_0_ ( .D(n427), .CK(i_CLK), .Q(z_e[0]) );
  fd1qd1_hd b_e_reg_4_ ( .D(n494), .CK(i_CLK), .Q(b_e[4]) );
  fd1qd1_hd a_e_reg_6_ ( .D(n482), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd b_e_reg_2_ ( .D(n496), .CK(i_CLK), .Q(b_e[2]) );
  fd1qd1_hd a_e_reg_4_ ( .D(n484), .CK(i_CLK), .Q(a_e[4]) );
  fd1qd1_hd a_e_reg_2_ ( .D(n486), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1581), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n509), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n509), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n509), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1581), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1581), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1581), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1581), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1581), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_0_ ( .D(z[0]), .E(n1581), .CK(i_CLK), .Q(o_Z[0]) );
  fd1eqd1_hd o_Z_reg_1_ ( .D(z[1]), .E(n1581), .CK(i_CLK), .Q(o_Z[1]) );
  fd1eqd1_hd o_Z_reg_2_ ( .D(z[2]), .E(n1581), .CK(i_CLK), .Q(o_Z[2]) );
  fd1eqd1_hd o_Z_reg_3_ ( .D(z[3]), .E(n1581), .CK(i_CLK), .Q(o_Z[3]) );
  fd1eqd1_hd o_Z_reg_4_ ( .D(z[4]), .E(n1581), .CK(i_CLK), .Q(o_Z[4]) );
  fd1eqd1_hd o_Z_reg_5_ ( .D(z[5]), .E(n1581), .CK(i_CLK), .Q(o_Z[5]) );
  fd1eqd1_hd o_Z_reg_6_ ( .D(z[6]), .E(n1581), .CK(i_CLK), .Q(o_Z[6]) );
  fd1eqd1_hd o_Z_reg_7_ ( .D(z[7]), .E(n1581), .CK(i_CLK), .Q(o_Z[7]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1581), .CK(i_CLK), .Q(o_Z[8]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1581), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1581), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1581), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1581), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n509), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n509), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n509), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n509), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1581), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1581), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n1581), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1581), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1581), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1581), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd b_reg_31_ ( .D(i_B[31]), .E(n1571), .CK(i_CLK), .Q(b[31]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n1571), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n1571), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd b_reg_30_ ( .D(i_B[30]), .E(n1571), .CK(i_CLK), .Q(b[30]) );
  fd1eqd1_hd z_s_reg ( .D(N338), .E(n1570), .CK(i_CLK), .Q(z_s) );
  fd1eqd1_hd sum_reg_0_ ( .D(N310), .E(n1570), .CK(i_CLK), .Q(sum[0]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n1571), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n1571), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n1571), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n1571), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n1571), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n1571), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n1571), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n1571), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n1571), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n1571), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n1571), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n1571), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n1571), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n1571), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n1571), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n1571), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n1571), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n1571), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n1571), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n1571), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n1571), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n1571), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n1571), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd b_reg_0_ ( .D(i_B[0]), .E(n1571), .CK(i_CLK), .Q(b[0]) );
  fd1eqd1_hd b_reg_1_ ( .D(i_B[1]), .E(n1571), .CK(i_CLK), .Q(b[1]) );
  fd1eqd1_hd b_reg_2_ ( .D(i_B[2]), .E(n1571), .CK(i_CLK), .Q(b[2]) );
  fd1eqd1_hd b_reg_3_ ( .D(i_B[3]), .E(n1571), .CK(i_CLK), .Q(b[3]) );
  fd1eqd1_hd b_reg_4_ ( .D(i_B[4]), .E(n1571), .CK(i_CLK), .Q(b[4]) );
  fd1eqd1_hd b_reg_5_ ( .D(i_B[5]), .E(n1571), .CK(i_CLK), .Q(b[5]) );
  fd1eqd1_hd b_reg_6_ ( .D(i_B[6]), .E(n1571), .CK(i_CLK), .Q(b[6]) );
  fd1eqd1_hd b_reg_7_ ( .D(i_B[7]), .E(n1571), .CK(i_CLK), .Q(b[7]) );
  fd1eqd1_hd b_reg_8_ ( .D(i_B[8]), .E(n1571), .CK(i_CLK), .Q(b[8]) );
  fd1eqd1_hd b_reg_9_ ( .D(i_B[9]), .E(n1571), .CK(i_CLK), .Q(b[9]) );
  fd1eqd1_hd b_reg_10_ ( .D(i_B[10]), .E(n1571), .CK(i_CLK), .Q(b[10]) );
  fd1eqd1_hd b_reg_11_ ( .D(i_B[11]), .E(n1571), .CK(i_CLK), .Q(b[11]) );
  fd1eqd1_hd b_reg_12_ ( .D(i_B[12]), .E(n1571), .CK(i_CLK), .Q(b[12]) );
  fd1eqd1_hd b_reg_13_ ( .D(i_B[13]), .E(n1571), .CK(i_CLK), .Q(b[13]) );
  fd1eqd1_hd b_reg_14_ ( .D(i_B[14]), .E(n1571), .CK(i_CLK), .Q(b[14]) );
  fd1eqd1_hd b_reg_15_ ( .D(i_B[15]), .E(n1571), .CK(i_CLK), .Q(b[15]) );
  fd1eqd1_hd b_reg_16_ ( .D(i_B[16]), .E(n1571), .CK(i_CLK), .Q(b[16]) );
  fd1eqd1_hd b_reg_17_ ( .D(i_B[17]), .E(n1571), .CK(i_CLK), .Q(b[17]) );
  fd1eqd1_hd b_reg_18_ ( .D(i_B[18]), .E(n1571), .CK(i_CLK), .Q(b[18]) );
  fd1eqd1_hd b_reg_19_ ( .D(i_B[19]), .E(n1571), .CK(i_CLK), .Q(b[19]) );
  fd1eqd1_hd b_reg_20_ ( .D(i_B[20]), .E(n1571), .CK(i_CLK), .Q(b[20]) );
  fd1eqd1_hd b_reg_21_ ( .D(i_B[21]), .E(n1571), .CK(i_CLK), .Q(b[21]) );
  fd1eqd1_hd b_reg_22_ ( .D(i_B[22]), .E(n1571), .CK(i_CLK), .Q(b[22]) );
  fd1qd1_hd z_reg_1_ ( .D(n391), .CK(i_CLK), .Q(z[1]) );
  fd1qd1_hd z_reg_2_ ( .D(n390), .CK(i_CLK), .Q(z[2]) );
  fd1qd1_hd z_reg_3_ ( .D(n389), .CK(i_CLK), .Q(z[3]) );
  fd1qd1_hd z_reg_5_ ( .D(n387), .CK(i_CLK), .Q(z[5]) );
  fd1qd1_hd z_reg_12_ ( .D(n380), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_13_ ( .D(n379), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_14_ ( .D(n378), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_15_ ( .D(n377), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_16_ ( .D(n376), .CK(i_CLK), .Q(z[16]) );
  fd1eqd1_hd sum_reg_3_ ( .D(N313), .E(n1570), .CK(i_CLK), .Q(sum[3]) );
  fd1qd1_hd z_reg_31_ ( .D(n361), .CK(i_CLK), .Q(z[31]) );
  fd1eqd1_hd sum_reg_2_ ( .D(N312), .E(n1570), .CK(i_CLK), .Q(sum[2]) );
  fd1qd1_hd z_reg_22_ ( .D(n370), .CK(i_CLK), .Q(z[22]) );
  fd1eqd1_hd sum_reg_26_ ( .D(N336), .E(n1570), .CK(i_CLK), .Q(sum[26]) );
  fd1eqd1_hd sum_reg_4_ ( .D(N314), .E(n1570), .CK(i_CLK), .Q(sum[4]) );
  fd1eqd1_hd sum_reg_5_ ( .D(N315), .E(n1570), .CK(i_CLK), .Q(sum[5]) );
  fd1eqd1_hd sum_reg_6_ ( .D(N316), .E(n1570), .CK(i_CLK), .Q(sum[6]) );
  fd1eqd1_hd sum_reg_7_ ( .D(N317), .E(n1570), .CK(i_CLK), .Q(sum[7]) );
  fd1eqd1_hd sum_reg_8_ ( .D(N318), .E(n1570), .CK(i_CLK), .Q(sum[8]) );
  fd1eqd1_hd sum_reg_9_ ( .D(N319), .E(n1570), .CK(i_CLK), .Q(sum[9]) );
  fd1eqd1_hd sum_reg_10_ ( .D(N320), .E(n1570), .CK(i_CLK), .Q(sum[10]) );
  fd1eqd1_hd sum_reg_11_ ( .D(N321), .E(n1570), .CK(i_CLK), .Q(sum[11]) );
  fd1eqd1_hd sum_reg_12_ ( .D(N322), .E(n1570), .CK(i_CLK), .Q(sum[12]) );
  fd1eqd1_hd sum_reg_13_ ( .D(N323), .E(n1570), .CK(i_CLK), .Q(sum[13]) );
  fd1eqd1_hd sum_reg_14_ ( .D(N324), .E(n1570), .CK(i_CLK), .Q(sum[14]) );
  fd1eqd1_hd sum_reg_15_ ( .D(N325), .E(n1570), .CK(i_CLK), .Q(sum[15]) );
  fd1eqd1_hd sum_reg_16_ ( .D(N326), .E(n1570), .CK(i_CLK), .Q(sum[16]) );
  fd1eqd1_hd sum_reg_17_ ( .D(N327), .E(n1570), .CK(i_CLK), .Q(sum[17]) );
  fd1eqd1_hd sum_reg_18_ ( .D(N328), .E(n1570), .CK(i_CLK), .Q(sum[18]) );
  fd1eqd1_hd sum_reg_19_ ( .D(N329), .E(n1570), .CK(i_CLK), .Q(sum[19]) );
  fd1eqd1_hd sum_reg_20_ ( .D(N330), .E(n1570), .CK(i_CLK), .Q(sum[20]) );
  fd1eqd1_hd sum_reg_21_ ( .D(N331), .E(n1570), .CK(i_CLK), .Q(sum[21]) );
  fd1eqd1_hd sum_reg_22_ ( .D(N332), .E(n1570), .CK(i_CLK), .Q(sum[22]) );
  fd1eqd1_hd sum_reg_23_ ( .D(N333), .E(n1570), .CK(i_CLK), .Q(sum[23]) );
  fd1eqd1_hd sum_reg_24_ ( .D(N334), .E(n1570), .CK(i_CLK), .Q(sum[24]) );
  fd1eqd1_hd sum_reg_25_ ( .D(N335), .E(n1570), .CK(i_CLK), .Q(sum[25]) );
  fd1eqd1_hd sum_reg_1_ ( .D(N311), .E(n1570), .CK(i_CLK), .Q(sum[1]) );
  fd1qd1_hd z_reg_30_ ( .D(n362), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_28_ ( .D(n364), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_26_ ( .D(n366), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_24_ ( .D(n368), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n369), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_29_ ( .D(n363), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_27_ ( .D(n365), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_25_ ( .D(n367), .CK(i_CLK), .Q(z[25]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n1571), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n1571), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd b_reg_27_ ( .D(i_B[27]), .E(n1571), .CK(i_CLK), .Q(b[27]) );
  fd1eqd1_hd b_reg_29_ ( .D(i_B[29]), .E(n1571), .CK(i_CLK), .Q(b[29]) );
  fd1eqd1_hd sum_reg_27_ ( .D(N337), .E(n1570), .CK(i_CLK), .Q(sum[27]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n1571), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd b_reg_28_ ( .D(i_B[28]), .E(n1571), .CK(i_CLK), .Q(b[28]) );
  fd1qd1_hd z_m_reg_18_ ( .D(n399), .CK(i_CLK), .Q(z_m[18]) );
  fd1qd1_hd z_m_reg_21_ ( .D(n396), .CK(i_CLK), .Q(z_m[21]) );
  fd1qd1_hd z_m_reg_22_ ( .D(n395), .CK(i_CLK), .Q(z_m[22]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n1571), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd b_reg_25_ ( .D(i_B[25]), .E(n1571), .CK(i_CLK), .Q(b[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n1571), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd b_reg_24_ ( .D(i_B[24]), .E(n1571), .CK(i_CLK), .Q(b[24]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n1571), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd b_reg_26_ ( .D(i_B[26]), .E(n1571), .CK(i_CLK), .Q(b[26]) );
  fd1qd1_hd z_m_reg_20_ ( .D(n397), .CK(i_CLK), .Q(z_m[20]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n1571), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd b_reg_23_ ( .D(i_B[23]), .E(n1571), .CK(i_CLK), .Q(b[23]) );
  fd1qd1_hd z_m_reg_16_ ( .D(n401), .CK(i_CLK), .Q(z_m[16]) );
  fd1eqd1_hd guard_reg ( .D(n266), .E(n265), .CK(i_CLK), .Q(guard) );
  fd1qd1_hd z_m_reg_14_ ( .D(n403), .CK(i_CLK), .Q(z_m[14]) );
  fd1qd1_hd z_m_reg_19_ ( .D(n398), .CK(i_CLK), .Q(z_m[19]) );
  fd1qd1_hd z_m_reg_15_ ( .D(n402), .CK(i_CLK), .Q(z_m[15]) );
  fd1qd1_hd z_m_reg_17_ ( .D(n400), .CK(i_CLK), .Q(z_m[17]) );
  fd1qd1_hd z_m_reg_13_ ( .D(n404), .CK(i_CLK), .Q(z_m[13]) );
  fd1qd1_hd z_m_reg_12_ ( .D(n405), .CK(i_CLK), .Q(z_m[12]) );
  fd1qd1_hd z_m_reg_8_ ( .D(n409), .CK(i_CLK), .Q(z_m[8]) );
  fd1qd1_hd z_m_reg_10_ ( .D(n407), .CK(i_CLK), .Q(z_m[10]) );
  fd1qd1_hd z_m_reg_6_ ( .D(n411), .CK(i_CLK), .Q(z_m[6]) );
  fd1qd1_hd z_m_reg_11_ ( .D(n406), .CK(i_CLK), .Q(z_m[11]) );
  fd1qd1_hd z_m_reg_7_ ( .D(n410), .CK(i_CLK), .Q(z_m[7]) );
  fd1qd1_hd z_m_reg_23_ ( .D(n418), .CK(i_CLK), .Q(z_m[23]) );
  fd1qd1_hd z_m_reg_9_ ( .D(n408), .CK(i_CLK), .Q(z_m[9]) );
  fd1qd1_hd z_e_reg_1_ ( .D(n426), .CK(i_CLK), .Q(z_e[1]) );
  fd1qd1_hd z_e_reg_8_ ( .D(n419), .CK(i_CLK), .Q(z_e[8]) );
  fd1qd1_hd z_e_reg_9_ ( .D(n428), .CK(i_CLK), .Q(z_e[9]) );
  fd1qd1_hd z_m_reg_5_ ( .D(n412), .CK(i_CLK), .Q(z_m[5]) );
  fd1qd1_hd z_e_reg_7_ ( .D(n420), .CK(i_CLK), .Q(z_e[7]) );
  fd1qd1_hd z_m_reg_4_ ( .D(n413), .CK(i_CLK), .Q(z_m[4]) );
  fd1qd1_hd z_m_reg_0_ ( .D(n417), .CK(i_CLK), .Q(z_m[0]) );
  fd1qd1_hd z_m_reg_2_ ( .D(n415), .CK(i_CLK), .Q(z_m[2]) );
  fd1qd1_hd z_e_reg_5_ ( .D(n422), .CK(i_CLK), .Q(z_e[5]) );
  fd1qd1_hd z_m_reg_3_ ( .D(n414), .CK(i_CLK), .Q(z_m[3]) );
  fd1qd1_hd z_e_reg_2_ ( .D(n425), .CK(i_CLK), .Q(z_e[2]) );
  fd1qd1_hd z_e_reg_3_ ( .D(n424), .CK(i_CLK), .Q(z_e[3]) );
  fd1qd1_hd z_e_reg_4_ ( .D(n423), .CK(i_CLK), .Q(z_e[4]) );
  fd1qd1_hd z_e_reg_6_ ( .D(n421), .CK(i_CLK), .Q(z_e[6]) );
  fd1qd1_hd z_m_reg_1_ ( .D(n416), .CK(i_CLK), .Q(z_m[1]) );
  fd1qd1_hd state_reg_1_ ( .D(n501), .CK(i_CLK), .Q(state[1]) );
  fd1qd1_hd state_reg_2_ ( .D(n500), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd b_e_reg_6_ ( .D(n492), .CK(i_CLK), .Q(b_e[6]) );
  fd1qd1_hd b_e_reg_9_ ( .D(n504), .CK(i_CLK), .Q(b_e[9]) );
  fd1qd1_hd a_e_reg_9_ ( .D(n489), .CK(i_CLK), .Q(a_e[9]) );
  fd1qd1_hd b_e_reg_8_ ( .D(n490), .CK(i_CLK), .Q(b_e[8]) );
  fd1qd1_hd a_e_reg_8_ ( .D(n480), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_3_ ( .D(n505), .CK(i_CLK), .Q(state[3]) );
  fd1qd1_hd a_e_reg_5_ ( .D(n483), .CK(i_CLK), .Q(a_e[5]) );
  fd1qd1_hd a_e_reg_7_ ( .D(n481), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_e_reg_1_ ( .D(n487), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_e_reg_3_ ( .D(n485), .CK(i_CLK), .Q(a_e[3]) );
  fd1qd1_hd b_e_reg_3_ ( .D(n495), .CK(i_CLK), .Q(b_e[3]) );
  fd1qd1_hd b_e_reg_5_ ( .D(n493), .CK(i_CLK), .Q(b_e[5]) );
  fd1qd1_hd b_e_reg_1_ ( .D(n497), .CK(i_CLK), .Q(b_e[1]) );
  fd1qd1_hd state_reg_0_ ( .D(n502), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd a_e_reg_0_ ( .D(n488), .CK(i_CLK), .Q(a_e[0]) );
  fd1qd1_hd b_e_reg_7_ ( .D(n491), .CK(i_CLK), .Q(b_e[7]) );
  fd1qd1_hd b_e_reg_0_ ( .D(n498), .CK(i_CLK), .Q(b_e[0]) );
  fd1eqd1_hd b_s_reg ( .D(b[31]), .E(n1578), .CK(i_CLK), .Q(b_s) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n1578), .CK(i_CLK), .Q(a_s) );
  fd1qd1_hd a_m_reg_25_ ( .D(n479), .CK(i_CLK), .Q(a_m[25]) );
  fd1eqd1_hd a_m_reg_26_ ( .D(n2267), .E(n1), .CK(i_CLK), .Q(a_m[26]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n454), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd b_m_reg_24_ ( .D(n429), .CK(i_CLK), .Q(b_m[24]) );
  fd1qd1_hd b_m_reg_21_ ( .D(n432), .CK(i_CLK), .Q(b_m[21]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n455), .CK(i_CLK), .Q(a_m[23]) );
  fd1eqd1_hd b_m_reg_26_ ( .D(n2267), .E(n2), .CK(i_CLK), .Q(b_m[26]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n461), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd b_m_reg_15_ ( .D(n438), .CK(i_CLK), .Q(b_m[15]) );
  fd1qd1_hd b_m_reg_16_ ( .D(n437), .CK(i_CLK), .Q(b_m[16]) );
  fd1qd1_hd b_m_reg_13_ ( .D(n440), .CK(i_CLK), .Q(b_m[13]) );
  fd1qd1_hd b_m_reg_10_ ( .D(n443), .CK(i_CLK), .Q(b_m[10]) );
  fd1qd1_hd b_m_reg_18_ ( .D(n435), .CK(i_CLK), .Q(b_m[18]) );
  fd1qd1_hd b_m_reg_25_ ( .D(n503), .CK(i_CLK), .Q(b_m[25]) );
  fd1qd1_hd b_m_reg_19_ ( .D(n434), .CK(i_CLK), .Q(b_m[19]) );
  fd1qd1_hd b_m_reg_17_ ( .D(n436), .CK(i_CLK), .Q(b_m[17]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n457), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n469), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd b_m_reg_14_ ( .D(n439), .CK(i_CLK), .Q(b_m[14]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n459), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n465), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd b_m_reg_8_ ( .D(n445), .CK(i_CLK), .Q(b_m[8]) );
  fd1qd1_hd b_m_reg_11_ ( .D(n442), .CK(i_CLK), .Q(b_m[11]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n456), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n467), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd b_m_reg_23_ ( .D(n430), .CK(i_CLK), .Q(b_m[23]) );
  fd1qd1_hd b_m_reg_12_ ( .D(n441), .CK(i_CLK), .Q(b_m[12]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n463), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n458), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd b_m_reg_7_ ( .D(n446), .CK(i_CLK), .Q(b_m[7]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n466), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd b_m_reg_22_ ( .D(n431), .CK(i_CLK), .Q(b_m[22]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n468), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n460), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n464), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n462), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n470), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd b_m_reg_20_ ( .D(n433), .CK(i_CLK), .Q(b_m[20]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n478), .CK(i_CLK), .Q(a_m[0]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n477), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n476), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n471), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd b_m_reg_0_ ( .D(n453), .CK(i_CLK), .Q(b_m[0]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n473), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n475), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd b_m_reg_3_ ( .D(n450), .CK(i_CLK), .Q(b_m[3]) );
  fd1qd1_hd b_m_reg_6_ ( .D(n447), .CK(i_CLK), .Q(b_m[6]) );
  fd1qd1_hd b_m_reg_4_ ( .D(n449), .CK(i_CLK), .Q(b_m[4]) );
  fd1qd1_hd b_m_reg_9_ ( .D(n444), .CK(i_CLK), .Q(b_m[9]) );
  fd1qd1_hd b_m_reg_1_ ( .D(n452), .CK(i_CLK), .Q(b_m[1]) );
  fd1qd1_hd b_m_reg_2_ ( .D(n451), .CK(i_CLK), .Q(b_m[2]) );
  fd1qd1_hd b_m_reg_5_ ( .D(n448), .CK(i_CLK), .Q(b_m[5]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n474), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n472), .CK(i_CLK), .Q(a_m[6]) );
  fad1_hd DP_OP_43J4_124_6938_U28 ( .A(C2_Z_0), .B(n2265), .CI(
        DP_OP_43J4_124_6938_n58), .CO(DP_OP_43J4_124_6938_n27), .S(N310) );
  fad1_hd DP_OP_43J4_124_6938_U27 ( .A(DP_OP_43J4_124_6938_n57), .B(C2_Z_1), 
        .CI(DP_OP_43J4_124_6938_n27), .CO(DP_OP_43J4_124_6938_n26), .S(N311)
         );
  fad1_hd DP_OP_43J4_124_6938_U26 ( .A(DP_OP_43J4_124_6938_n56), .B(C2_Z_2), 
        .CI(DP_OP_43J4_124_6938_n26), .CO(DP_OP_43J4_124_6938_n25), .S(N312)
         );
  fad1_hd DP_OP_43J4_124_6938_U25 ( .A(DP_OP_43J4_124_6938_n55), .B(C2_Z_3), 
        .CI(DP_OP_43J4_124_6938_n25), .CO(DP_OP_43J4_124_6938_n24), .S(N313)
         );
  fad1_hd DP_OP_43J4_124_6938_U24 ( .A(DP_OP_43J4_124_6938_n54), .B(C2_Z_4), 
        .CI(DP_OP_43J4_124_6938_n24), .CO(DP_OP_43J4_124_6938_n23), .S(N314)
         );
  fad1_hd DP_OP_43J4_124_6938_U23 ( .A(DP_OP_43J4_124_6938_n53), .B(C2_Z_5), 
        .CI(DP_OP_43J4_124_6938_n23), .CO(DP_OP_43J4_124_6938_n22), .S(N315)
         );
  fad1_hd DP_OP_43J4_124_6938_U2 ( .A(DP_OP_43J4_124_6938_n32), .B(C2_Z_26), 
        .CI(DP_OP_43J4_124_6938_n2), .CO(DP_OP_43J4_124_6938_n1), .S(N336) );
  fad1_hd DP_OP_43J4_124_6938_U3 ( .A(DP_OP_43J4_124_6938_n33), .B(C2_Z_25), 
        .CI(DP_OP_43J4_124_6938_n3), .CO(DP_OP_43J4_124_6938_n2), .S(N335) );
  fad1_hd DP_OP_43J4_124_6938_U4 ( .A(DP_OP_43J4_124_6938_n34), .B(C2_Z_24), 
        .CI(DP_OP_43J4_124_6938_n4), .CO(DP_OP_43J4_124_6938_n3), .S(N334) );
  fad1_hd DP_OP_43J4_124_6938_U14 ( .A(DP_OP_43J4_124_6938_n44), .B(C2_Z_14), 
        .CI(DP_OP_43J4_124_6938_n14), .CO(DP_OP_43J4_124_6938_n13), .S(N324)
         );
  fad1_hd DP_OP_43J4_124_6938_U15 ( .A(DP_OP_43J4_124_6938_n45), .B(C2_Z_13), 
        .CI(DP_OP_43J4_124_6938_n15), .CO(DP_OP_43J4_124_6938_n14), .S(N323)
         );
  fad1_hd DP_OP_43J4_124_6938_U16 ( .A(DP_OP_43J4_124_6938_n46), .B(C2_Z_12), 
        .CI(DP_OP_43J4_124_6938_n16), .CO(DP_OP_43J4_124_6938_n15), .S(N322)
         );
  fad1_hd DP_OP_43J4_124_6938_U17 ( .A(DP_OP_43J4_124_6938_n47), .B(C2_Z_11), 
        .CI(DP_OP_43J4_124_6938_n17), .CO(DP_OP_43J4_124_6938_n16), .S(N321)
         );
  fad1_hd DP_OP_43J4_124_6938_U18 ( .A(DP_OP_43J4_124_6938_n48), .B(C2_Z_10), 
        .CI(DP_OP_43J4_124_6938_n18), .CO(DP_OP_43J4_124_6938_n17), .S(N320)
         );
  fad1_hd DP_OP_43J4_124_6938_U19 ( .A(DP_OP_43J4_124_6938_n49), .B(C2_Z_9), 
        .CI(DP_OP_43J4_124_6938_n19), .CO(DP_OP_43J4_124_6938_n18), .S(N319)
         );
  fad1_hd DP_OP_43J4_124_6938_U20 ( .A(DP_OP_43J4_124_6938_n50), .B(C2_Z_8), 
        .CI(DP_OP_43J4_124_6938_n20), .CO(DP_OP_43J4_124_6938_n19), .S(N318)
         );
  fad1_hd DP_OP_43J4_124_6938_U21 ( .A(DP_OP_43J4_124_6938_n51), .B(C2_Z_7), 
        .CI(DP_OP_43J4_124_6938_n21), .CO(DP_OP_43J4_124_6938_n20), .S(N317)
         );
  fad1_hd DP_OP_43J4_124_6938_U22 ( .A(DP_OP_43J4_124_6938_n52), .B(C2_Z_6), 
        .CI(DP_OP_43J4_124_6938_n22), .CO(DP_OP_43J4_124_6938_n21), .S(N316)
         );
  fad1_hd DP_OP_43J4_124_6938_U13 ( .A(DP_OP_43J4_124_6938_n43), .B(C2_Z_15), 
        .CI(DP_OP_43J4_124_6938_n13), .CO(DP_OP_43J4_124_6938_n12), .S(N325)
         );
  fad1_hd DP_OP_43J4_124_6938_U12 ( .A(DP_OP_43J4_124_6938_n42), .B(C2_Z_16), 
        .CI(DP_OP_43J4_124_6938_n12), .CO(DP_OP_43J4_124_6938_n11), .S(N326)
         );
  fad1_hd DP_OP_43J4_124_6938_U11 ( .A(DP_OP_43J4_124_6938_n41), .B(C2_Z_17), 
        .CI(DP_OP_43J4_124_6938_n11), .CO(DP_OP_43J4_124_6938_n10), .S(N327)
         );
  fad1_hd DP_OP_43J4_124_6938_U10 ( .A(DP_OP_43J4_124_6938_n40), .B(C2_Z_18), 
        .CI(DP_OP_43J4_124_6938_n10), .CO(DP_OP_43J4_124_6938_n9), .S(N328) );
  fad1_hd DP_OP_43J4_124_6938_U9 ( .A(DP_OP_43J4_124_6938_n39), .B(C2_Z_19), 
        .CI(DP_OP_43J4_124_6938_n9), .CO(DP_OP_43J4_124_6938_n8), .S(N329) );
  fad1_hd DP_OP_43J4_124_6938_U8 ( .A(DP_OP_43J4_124_6938_n38), .B(C2_Z_20), 
        .CI(DP_OP_43J4_124_6938_n8), .CO(DP_OP_43J4_124_6938_n7), .S(N330) );
  fad1_hd DP_OP_43J4_124_6938_U7 ( .A(DP_OP_43J4_124_6938_n37), .B(C2_Z_21), 
        .CI(DP_OP_43J4_124_6938_n7), .CO(DP_OP_43J4_124_6938_n6), .S(N331) );
  fad1_hd DP_OP_43J4_124_6938_U6 ( .A(DP_OP_43J4_124_6938_n36), .B(C2_Z_22), 
        .CI(DP_OP_43J4_124_6938_n6), .CO(DP_OP_43J4_124_6938_n5), .S(N332) );
  fad1_hd DP_OP_43J4_124_6938_U5 ( .A(DP_OP_43J4_124_6938_n35), .B(C2_Z_23), 
        .CI(DP_OP_43J4_124_6938_n5), .CO(DP_OP_43J4_124_6938_n4), .S(N333) );
  fd1qd1_hd o_AB_ACK_reg ( .D(n499), .CK(i_CLK), .Q(o_AB_ACK) );
  fd1qd1_hd sticky_reg ( .D(n393), .CK(i_CLK), .Q(sticky) );
  fd1qd1_hd round_bit_reg ( .D(n394), .CK(i_CLK), .Q(round_bit) );
  fd1qd1_hd o_Z_STB_reg ( .D(n506), .CK(i_CLK), .Q(o_Z_STB) );
  fd1qd1_hd z_reg_11_ ( .D(n381), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n382), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_9_ ( .D(n383), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n384), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_7_ ( .D(n385), .CK(i_CLK), .Q(z[7]) );
  fd1qd1_hd z_reg_6_ ( .D(n386), .CK(i_CLK), .Q(z[6]) );
  fd1qd1_hd z_reg_0_ ( .D(n392), .CK(i_CLK), .Q(z[0]) );
  fd1qd1_hd z_reg_4_ ( .D(n388), .CK(i_CLK), .Q(z[4]) );
  fd1qd1_hd z_reg_21_ ( .D(n371), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n372), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n373), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n374), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_17_ ( .D(n375), .CK(i_CLK), .Q(z[17]) );
  nr2d1_hd U523 ( .A(n1988), .B(n1932), .Y(n1949) );
  clknd2d1_hd U524 ( .A(b_m[5]), .B(n2081), .Y(n1588) );
  clknd2d1_hd U525 ( .A(n1596), .B(n1595), .Y(n1597) );
  clknd2d1_hd U526 ( .A(b_m[18]), .B(n1612), .Y(n1613) );
  clknd2d1_hd U527 ( .A(b_m[8]), .B(n2075), .Y(n1593) );
  clknd2d1_hd U528 ( .A(n1591), .B(b_m[7]), .Y(n1592) );
  clknd2d1_hd U529 ( .A(b_m[12]), .B(n2067), .Y(n1601) );
  clknd2d1_hd U530 ( .A(b_m[11]), .B(n1599), .Y(n1600) );
  clknd2d1_hd U531 ( .A(b_m[17]), .B(n2057), .Y(n1611) );
  clknd2d1_hd U532 ( .A(b_e[8]), .B(n2099), .Y(n1697) );
  clknd2d1_hd U533 ( .A(n1680), .B(n1679), .Y(n1688) );
  clknd2d1_hd U534 ( .A(b_e[6]), .B(n2097), .Y(n1679) );
  clknd2d1_hd U535 ( .A(a_e[9]), .B(n1683), .Y(n1700) );
  clknd2d1_hd U536 ( .A(b_m[19]), .B(n2053), .Y(n1614) );
  clknd2d1_hd U537 ( .A(n1717), .B(n1715), .Y(n1719) );
  clknd2d1_hd U538 ( .A(n1750), .B(n1792), .Y(n1716) );
  clknd2d1_hd U539 ( .A(n1700), .B(n1699), .Y(n1701) );
  clknd2d1_hd U540 ( .A(a_e[8]), .B(n2166), .Y(n1694) );
  clknd2d1_hd U541 ( .A(n2186), .B(n1701), .Y(n2232) );
  clknd2d1_hd U542 ( .A(n1705), .B(n1727), .Y(n2228) );
  clknd2d1_hd U543 ( .A(n1712), .B(n2094), .Y(n1715) );
  clknd2d1_hd U544 ( .A(n2160), .B(n1711), .Y(n1717) );
  clknd2d1_hd U545 ( .A(n1703), .B(z_e[1]), .Y(n1727) );
  clknd2d1_hd U546 ( .A(a_e[4]), .B(n2118), .Y(n2096) );
  clknd2d1_hd U547 ( .A(state[0]), .B(n2240), .Y(n2225) );
  clknd2d1_hd U548 ( .A(n1971), .B(guard), .Y(n1963) );
  clknd2d1_hd U549 ( .A(n1576), .B(n2186), .Y(n2249) );
  clknd2d1_hd U550 ( .A(n1718), .B(n2260), .Y(n1707) );
  clknd2d1_hd U551 ( .A(n1574), .B(n2186), .Y(n2091) );
  clknd2d1_hd U552 ( .A(n2185), .B(n2163), .Y(n2170) );
  clknd2d1_hd U553 ( .A(n2246), .B(n2240), .Y(n2243) );
  clknd2d1_hd U554 ( .A(n2202), .B(n2212), .Y(n2210) );
  clknd2d1_hd U555 ( .A(b_e[2]), .B(n2201), .Y(n2195) );
  clknd2d1_hd U556 ( .A(a_e[2]), .B(n2133), .Y(n2127) );
  clknd2d1_hd U557 ( .A(n2136), .B(n2128), .Y(n2126) );
  clknd2d1_hd U558 ( .A(n2136), .B(n2145), .Y(n2143) );
  clknd2d1_hd U559 ( .A(n2117), .B(n2095), .Y(n2103) );
  clknd2d1_hd U560 ( .A(n2177), .B(n2173), .Y(n2253) );
  clknd2d1_hd U561 ( .A(b_e[5]), .B(n2180), .Y(n2179) );
  clknd2d1_hd U562 ( .A(n2191), .B(b_e[4]), .Y(n2162) );
  clknd2d1_hd U563 ( .A(n2187), .B(b[28]), .Y(n2181) );
  clknd2d1_hd U564 ( .A(state[2]), .B(n2260), .Y(n2244) );
  clknd2d1_hd U565 ( .A(N41), .B(n2259), .Y(n2261) );
  clknd2d1_hd U566 ( .A(n1955), .B(n1946), .Y(n1937) );
  clknd2d1_hd U567 ( .A(n1942), .B(n1937), .Y(n1933) );
  clknd2d1_hd U568 ( .A(n1955), .B(n1918), .Y(n1925) );
  clknd2d1_hd U569 ( .A(z_m[21]), .B(n1964), .Y(n1957) );
  clknd2d1_hd U570 ( .A(n1972), .B(sum[27]), .Y(n1969) );
  clknd2d1_hd U571 ( .A(n1955), .B(n1893), .Y(n1900) );
  clknd2d1_hd U572 ( .A(n1955), .B(n1869), .Y(n1876) );
  clknd2d1_hd U573 ( .A(n1955), .B(n1967), .Y(n1827) );
  clknd2d1_hd U574 ( .A(n1955), .B(n1845), .Y(n1852) );
  clknd2d1_hd U575 ( .A(z_m[20]), .B(n1823), .Y(n1958) );
  clknd2d1_hd U576 ( .A(z_m[19]), .B(z_m[20]), .Y(n1813) );
  clknd2d1_hd U577 ( .A(n2190), .B(n2121), .Y(n1758) );
  clknd2d1_hd U578 ( .A(n2164), .B(n2097), .Y(n1743) );
  clknd2d1_hd U579 ( .A(b_e[0]), .B(a_e[0]), .Y(n1786) );
  clknd2d1_hd U580 ( .A(n1751), .B(n1750), .Y(n1779) );
  clknd2d1_hd U581 ( .A(n1778), .B(n1773), .Y(n1772) );
  clknd2d1_hd U582 ( .A(n1764), .B(n1760), .Y(n1759) );
  clknd2d1_hd U583 ( .A(b_e[7]), .B(a_e[7]), .Y(n1738) );
  clknd2d1_hd U584 ( .A(n1749), .B(n1745), .Y(n1744) );
  clknd2d1_hd U585 ( .A(n1796), .B(n1735), .Y(n1790) );
  clknd2d1_hd U586 ( .A(n1726), .B(n1725), .Y(n1729) );
  nid1_hd U587 ( .A(n1802), .Y(n1572) );
  clknd2d1_hd U588 ( .A(state[1]), .B(n2246), .Y(n2222) );
  clknd2d1_hd U589 ( .A(state[3]), .B(n1718), .Y(n2221) );
  clknd2d1_hd U590 ( .A(a[23]), .B(a[24]), .Y(n2147) );
  clknd2d1_hd U591 ( .A(n2134), .B(a[26]), .Y(n2130) );
  clknd2d1_hd U592 ( .A(b[23]), .B(b[24]), .Y(n2214) );
  clknd2d1_hd U593 ( .A(n2213), .B(n2210), .Y(n2206) );
  clknd2d1_hd U594 ( .A(a_e[5]), .B(n2112), .Y(n2111) );
  clknd2d1_hd U595 ( .A(n2119), .B(a[28]), .Y(n2113) );
  clknd2d1_hd U596 ( .A(b_e[4]), .B(n2202), .Y(n2194) );
  clknd2d1_hd U597 ( .A(n2203), .B(b[26]), .Y(n2198) );
  clknd2d1_hd U598 ( .A(n1808), .B(n1807), .Y(n393) );
  clknd2d1_hd U599 ( .A(n1580), .B(n2167), .Y(n2172) );
  clknd2d1_hd U600 ( .A(n2200), .B(n2199), .Y(n495) );
  clknd2d1_hd U601 ( .A(a[30]), .B(n2100), .Y(n2105) );
  clknd2d1_hd U602 ( .A(n2181), .B(n2174), .Y(n2176) );
  clknd2d1_hd U603 ( .A(n1956), .B(n1937), .Y(n1939) );
  clknd2d1_hd U604 ( .A(n1993), .B(n1992), .Y(n428) );
  clknd2d1_hd U605 ( .A(DP_OP_154J4_137_6175_n2), .B(n1991), .Y(n1989) );
  clknd2d1_hd U606 ( .A(n1970), .B(n1805), .Y(n265) );
  clknd2d1_hd U607 ( .A(n1789), .B(n1741), .Y(n362) );
  clknd2d1_hd U608 ( .A(n2136), .B(n2133), .Y(n2142) );
  clknd2d1_hd U609 ( .A(n2136), .B(n2118), .Y(n2125) );
  clknd2d1_hd U610 ( .A(n2202), .B(n2201), .Y(n2209) );
  clknd2d1_hd U611 ( .A(n2113), .B(n2106), .Y(n2107) );
  ad2d4_hd U612 ( .A(n2265), .B(n1627), .Y(n1568) );
  ivd4_hd U613 ( .A(n1568), .Y(n1569) );
  ivd2_hd U614 ( .A(n1791), .Y(n2265) );
  ivd1_hd U615 ( .A(b_m[2]), .Y(n2039) );
  ivd1_hd U616 ( .A(b_m[1]), .Y(n2040) );
  ivd1_hd U617 ( .A(b_m[23]), .Y(n1997) );
  nr2d4_hd U618 ( .A(n1568), .B(n1791), .Y(n1655) );
  oa21d1_hd U619 ( .A(n1624), .B(n1623), .C(n1622), .Y(n1625) );
  ao21d1_hd U620 ( .A(a_m[23]), .B(n1997), .C(n1621), .Y(n1624) );
  ivd3_hd U621 ( .A(n2269), .Y(n1570) );
  ivd1_hd U622 ( .A(b_m[26]), .Y(n2250) );
  xo2d1_hd U623 ( .A(n2265), .B(DP_OP_43J4_124_6938_n1), .Y(N337) );
  nid6_hd U624 ( .A(n27), .Y(n1571) );
  ad3d1_hd U625 ( .A(n2220), .B(i_AB_STB), .C(o_AB_ACK), .Y(n27) );
  or2d2_hd U626 ( .A(n1707), .B(n2225), .Y(n2268) );
  scg9d1_hd U627 ( .A(n2238), .B(n1701), .C(n2268), .Y(n2158) );
  ad3d1_hd U628 ( .A(n2258), .B(n1577), .C(n2256), .Y(n2262) );
  scg2d1_hd U629 ( .A(b_e[9]), .B(n1698), .C(n1697), .D(n1696), .Y(n1699) );
  ivd2_hd U630 ( .A(n1779), .Y(n1804) );
  ivd2_hd U631 ( .A(n1969), .Y(n1943) );
  or4d1_hd U632 ( .A(z_m[23]), .B(z_e[0]), .C(n1728), .D(n1727), .Y(n1735) );
  or2d1_hd U633 ( .A(n2243), .B(n2244), .Y(n2269) );
  or4d1_hd U634 ( .A(n1678), .B(a_e[9]), .C(a_e[0]), .D(a_e[8]), .Y(n1792) );
  oa22d4_hd U635 ( .A(n1657), .B(n1709), .C(a_s), .D(b_s), .Y(n1791) );
  ivd1_hd U636 ( .A(b_m[0]), .Y(n2041) );
  or2d1_hd U637 ( .A(b_e[2]), .B(a_e[2]), .Y(n1771) );
  nr2d2_hd U638 ( .A(n1797), .B(n2224), .Y(n1803) );
  ivd2_hd U639 ( .A(n1949), .Y(n1956) );
  nr2ad1_hd U640 ( .A(n1973), .B(n1986), .Y(n1990) );
  nr2ad1_hd U641 ( .A(n2256), .B(n1932), .Y(n1938) );
  nr2ad1_hd U642 ( .A(n2222), .B(n2244), .Y(n2266) );
  oa22ad1_hd U643 ( .A(n1590), .B(a_m[6]), .C(n1589), .D(b_m[6]), .Y(n1591) );
  ivd1_hd U644 ( .A(b_m[3]), .Y(n2038) );
  ivd1_hd U645 ( .A(b_m[4]), .Y(n2035) );
  ao22d1_hd U646 ( .A(a_m[26]), .B(n2250), .C(n1626), .D(n1625), .Y(n1627) );
  ivd1_hd U647 ( .A(a_m[3]), .Y(n2086) );
  ivd1_hd U648 ( .A(a_m[5]), .Y(n2081) );
  ivd1_hd U649 ( .A(b_m[5]), .Y(n2033) );
  nid2_hd U650 ( .A(n2257), .Y(n1577) );
  ivd1_hd U651 ( .A(n1955), .Y(n1931) );
  ivd1_hd U652 ( .A(n1984), .Y(n1986) );
  ivd1_hd U653 ( .A(n2093), .Y(n1575) );
  oa21d1_hd U654 ( .A(a_m[21]), .B(n2001), .C(n1618), .Y(n1619) );
  ivd1_hd U655 ( .A(a_m[4]), .Y(n2083) );
  ivd1_hd U656 ( .A(n1787), .Y(n1800) );
  ivd1_hd U657 ( .A(n2268), .Y(n1578) );
  nr2d1_hd U658 ( .A(n2258), .B(n1932), .Y(n1955) );
  ivd1_hd U659 ( .A(n1971), .Y(n2258) );
  nid2_hd U660 ( .A(n1944), .Y(n1573) );
  ivd1_hd U661 ( .A(n1938), .Y(n1945) );
  nr2d1_hd U662 ( .A(n2221), .B(n2243), .Y(n1971) );
  ivd1_hd U663 ( .A(n2266), .Y(n1988) );
  ivd2_hd U664 ( .A(n2158), .Y(n1576) );
  ivd2_hd U665 ( .A(n1575), .Y(n1574) );
  ivd1_hd U666 ( .A(n2267), .Y(n2223) );
  ivd1_hd U667 ( .A(n2238), .Y(n2186) );
  nd2bd1_hd U668 ( .AN(n1707), .B(n2234), .Y(n2238) );
  ivd1_hd U669 ( .A(b_m[24]), .Y(n1995) );
  ivd1_hd U670 ( .A(a_m[16]), .Y(n2059) );
  ivd1_hd U671 ( .A(b_m[10]), .Y(n2023) );
  ivd1_hd U672 ( .A(b_m[13]), .Y(n2017) );
  ivd1_hd U673 ( .A(a_m[15]), .Y(n2061) );
  ivd1_hd U674 ( .A(b_m[14]), .Y(n2015) );
  ivd1_hd U675 ( .A(a_m[17]), .Y(n2057) );
  ivd1_hd U676 ( .A(b_m[17]), .Y(n2009) );
  ivd1_hd U677 ( .A(b_m[21]), .Y(n2001) );
  nid2_hd U678 ( .A(n509), .Y(n1581) );
  nr3d1_hd U679 ( .A(n1751), .B(n1717), .C(n1716), .Y(n1802) );
  ivd1_hd U680 ( .A(n1715), .Y(n1751) );
  ivd2_hd U681 ( .A(n2249), .Y(n2036) );
  scg20d2_hd U682 ( .A(n1812), .B(n1963), .C(n265), .Y(n1932) );
  ivd1_hd U683 ( .A(n1972), .Y(n1805) );
  ivd2_hd U684 ( .A(n2268), .Y(n1579) );
  ivd2_hd U685 ( .A(n2091), .Y(n2084) );
  nr2d1_hd U686 ( .A(n2225), .B(n2244), .Y(n1972) );
  nd2bd1_hd U687 ( .AN(n2244), .B(n2234), .Y(n2256) );
  ivd1_hd U688 ( .A(n2202), .Y(n2252) );
  nr2d1_hd U689 ( .A(n2218), .B(n2238), .Y(n2202) );
  ao21d1_hd U690 ( .A(n2160), .B(n2159), .C(n1576), .Y(n2218) );
  ivd1_hd U691 ( .A(n2268), .Y(n1580) );
  ivd1_hd U692 ( .A(n2136), .Y(n2154) );
  nr2d1_hd U693 ( .A(n2151), .B(n2238), .Y(n2136) );
  ao21d1_hd U694 ( .A(n2094), .B(n2159), .C(n1574), .Y(n2151) );
  scg16d1_hd U695 ( .A(n2233), .B(n2232), .C(n2268), .Y(n2093) );
  ivd1_hd U696 ( .A(b_e[1]), .Y(n2212) );
  nr2d1_hd U697 ( .A(n1719), .B(n1716), .Y(n2159) );
  nr2d1_hd U698 ( .A(n1707), .B(n2222), .Y(n2267) );
  ivd1_hd U699 ( .A(b_e[6]), .Y(n2164) );
  ivd1_hd U700 ( .A(a_e[8]), .Y(n2099) );
  ivd1_hd U701 ( .A(a_e[5]), .Y(n2116) );
  ivd1_hd U702 ( .A(a_e[6]), .Y(n2097) );
  nr2d1_hd U703 ( .A(n2246), .B(n2240), .Y(n2234) );
  ivd1_hd U704 ( .A(state[0]), .Y(n2246) );
  ivd1_hd U705 ( .A(state[1]), .Y(n2240) );
  ivd1_hd U706 ( .A(state[3]), .Y(n2260) );
  ivd1_hd U707 ( .A(b_m[25]), .Y(n1629) );
  ivd1_hd U708 ( .A(b_m[19]), .Y(n2005) );
  ivd1_hd U709 ( .A(b_m[20]), .Y(n2003) );
  ivd1_hd U710 ( .A(a_m[20]), .Y(n2051) );
  ivd1_hd U711 ( .A(b_m[22]), .Y(n1999) );
  ivd1_hd U712 ( .A(a_m[22]), .Y(n2047) );
  ivd1_hd U713 ( .A(a_m[25]), .Y(n1668) );
  ivd1_hd U714 ( .A(n2159), .Y(n2242) );
  nr2d1_hd U715 ( .A(n2222), .B(n2221), .Y(n509) );
  ivd1_hd U716 ( .A(n1796), .Y(n2224) );
  ivd1_hd U717 ( .A(z_m[1]), .Y(n1946) );
  ao21d1_hd U718 ( .A(n1796), .B(n1797), .C(n1734), .Y(n1789) );
  ivd1_hd U719 ( .A(n1710), .Y(n1793) );
  nr2d1_hd U720 ( .A(n2225), .B(n2221), .Y(n1796) );
  ivd1_hd U721 ( .A(z_m[20]), .Y(n1832) );
  ivd1_hd U722 ( .A(z_m[21]), .Y(n1826) );
  ivd1_hd U723 ( .A(n1932), .Y(n1952) );
  ivd1_hd U724 ( .A(z_m[22]), .Y(n1965) );
  ivd1_hd U725 ( .A(z_m[17]), .Y(n1850) );
  ivd1_hd U726 ( .A(z_m[18]), .Y(n1838) );
  ivd1_hd U727 ( .A(z_m[13]), .Y(n1874) );
  ivd1_hd U728 ( .A(z_m[14]), .Y(n1862) );
  ivd1_hd U729 ( .A(z_m[10]), .Y(n1886) );
  ivd1_hd U730 ( .A(z_m[9]), .Y(n1898) );
  ivd1_hd U731 ( .A(z_m[5]), .Y(n1923) );
  ivd1_hd U732 ( .A(z_m[6]), .Y(n1910) );
  ivd1_hd U733 ( .A(z_m[23]), .Y(n1964) );
  ivd1_hd U734 ( .A(z_e[0]), .Y(n1985) );
  ivd1_hd U735 ( .A(z_e[7]), .Y(n1733) );
  ivd1_hd U736 ( .A(z_e[8]), .Y(n1975) );
  ivd1_hd U737 ( .A(n2254), .Y(n2207) );
  nr2d1_hd U738 ( .A(n2223), .B(n2218), .Y(n2254) );
  ivd1_hd U739 ( .A(b[30]), .Y(n2173) );
  ivd1_hd U740 ( .A(n2156), .Y(n2140) );
  nr2d1_hd U741 ( .A(n2223), .B(n2151), .Y(n2156) );
  ivd1_hd U742 ( .A(a_e[7]), .Y(n2101) );
  ivd1_hd U743 ( .A(a_e[4]), .Y(n2121) );
  ivd1_hd U744 ( .A(a_e[2]), .Y(n2137) );
  ivd1_hd U745 ( .A(b_e[7]), .Y(n2168) );
  nr3d1_hd U746 ( .A(n1676), .B(n1675), .C(n1674), .Y(n1712) );
  ivd1_hd U747 ( .A(b_e[9]), .Y(n1683) );
  ivd1_hd U748 ( .A(b_e[0]), .Y(n2211) );
  ivd1_hd U749 ( .A(b_e[5]), .Y(n2184) );
  ivd1_hd U750 ( .A(b_e[8]), .Y(n2166) );
  ivd1_hd U751 ( .A(a_e[0]), .Y(n2144) );
  ivd1_hd U752 ( .A(a_e[1]), .Y(n2145) );
  ivd1_hd U753 ( .A(a_e[3]), .Y(n2128) );
  ivd1_hd U754 ( .A(state[2]), .Y(n1718) );
  ivd1_hd U755 ( .A(a_m[1]), .Y(n2088) );
  ivd1_hd U756 ( .A(a_m[2]), .Y(n2087) );
  ivd1_hd U757 ( .A(a_m[6]), .Y(n2079) );
  ivd1_hd U758 ( .A(b_m[6]), .Y(n2031) );
  ivd1_hd U759 ( .A(a_m[7]), .Y(n2077) );
  ivd1_hd U760 ( .A(b_m[7]), .Y(n2029) );
  ivd1_hd U761 ( .A(a_m[11]), .Y(n2069) );
  ivd1_hd U762 ( .A(b_m[11]), .Y(n2021) );
  ivd1_hd U763 ( .A(a_m[13]), .Y(n2065) );
  ivd1_hd U764 ( .A(a_m[14]), .Y(n2063) );
  ivd1_hd U765 ( .A(a_m[18]), .Y(n2055) );
  ivd1_hd U766 ( .A(b_m[18]), .Y(n2007) );
  ivd1_hd U767 ( .A(a_m[21]), .Y(n2049) );
  ivd1_hd U768 ( .A(a_m[23]), .Y(n2045) );
  ivd1_hd U769 ( .A(a_m[24]), .Y(n2043) );
  ivd1_hd U770 ( .A(a_m[19]), .Y(n2053) );
  ivd1_hd U771 ( .A(b_m[15]), .Y(n2013) );
  ivd1_hd U772 ( .A(b_m[16]), .Y(n2011) );
  ivd1_hd U773 ( .A(a_m[12]), .Y(n2067) );
  ivd1_hd U774 ( .A(a_m[8]), .Y(n2075) );
  ivd1_hd U775 ( .A(b_m[8]), .Y(n2027) );
  ivd1_hd U776 ( .A(b_m[9]), .Y(n2025) );
  ivd1_hd U777 ( .A(a_m[10]), .Y(n2071) );
  ivd1_hd U778 ( .A(a_m[9]), .Y(n2073) );
  ivd1_hd U779 ( .A(b_m[12]), .Y(n2019) );
  ivd1_hd U780 ( .A(a_m[26]), .Y(n2092) );
  ivd1_hd U781 ( .A(a_s), .Y(n1709) );
  ivd1_hd U782 ( .A(b_s), .Y(n1657) );
  ivd1_hd U783 ( .A(z_m[0]), .Y(n1953) );
  nr2d1_hd U784 ( .A(n1577), .B(n2223), .Y(n1787) );
  nd2bd1_hd U785 ( .AN(a[30]), .B(n2108), .Y(n2155) );
  ivd1_hd U786 ( .A(a_e[9]), .Y(n1698) );
  nr2d1_hd U787 ( .A(sum[27]), .B(n1805), .Y(n1944) );
  ao22d1_hd U788 ( .A(b_m[25]), .B(n1668), .C(b_m[26]), .D(n2092), .Y(n1626)
         );
  ao22d1_hd U789 ( .A(a_m[21]), .B(n2001), .C(a_m[22]), .D(n1999), .Y(n1620)
         );
  ao22d1_hd U790 ( .A(a_m[20]), .B(n2003), .C(a_m[19]), .D(n2005), .Y(n1617)
         );
  nr2d1_hd U791 ( .A(b_m[15]), .B(n2061), .Y(n1607) );
  ao22d1_hd U792 ( .A(a_m[13]), .B(n2017), .C(a_m[12]), .D(n2019), .Y(n1605)
         );
  ao22d1_hd U793 ( .A(b_m[9]), .B(n2073), .C(b_m[10]), .D(n2071), .Y(n1598) );
  ao22d1_hd U794 ( .A(a_m[9]), .B(n2025), .C(a_m[8]), .D(n2027), .Y(n1596) );
  ao211d1_hd U795 ( .A(a_m[1]), .B(n2040), .C(a_m[0]), .D(n2041), .Y(n1583) );
  oa22d1_hd U796 ( .A(a_m[1]), .B(n2040), .C(a_m[2]), .D(n2039), .Y(n1582) );
  oa22d1_hd U797 ( .A(b_m[3]), .B(n2086), .C(n1583), .D(n1582), .Y(n1584) );
  ao21d1_hd U798 ( .A(a_m[2]), .B(n2039), .C(n1584), .Y(n1586) );
  oa22d1_hd U799 ( .A(a_m[4]), .B(n2035), .C(a_m[3]), .D(n2038), .Y(n1585) );
  oa22d1_hd U800 ( .A(n1586), .B(n1585), .C(b_m[4]), .D(n2083), .Y(n1587) );
  ao22d1_hd U801 ( .A(a_m[5]), .B(n2033), .C(n1588), .D(n1587), .Y(n1589) );
  nr2d1_hd U802 ( .A(n1589), .B(b_m[6]), .Y(n1590) );
  nr2d1_hd U803 ( .A(n1591), .B(b_m[7]), .Y(n1594) );
  oa211d1_hd U804 ( .A(a_m[7]), .B(n1594), .C(n1593), .D(n1592), .Y(n1595) );
  ao22d1_hd U805 ( .A(a_m[10]), .B(n2023), .C(n1598), .D(n1597), .Y(n1599) );
  nr2d1_hd U806 ( .A(b_m[11]), .B(n1599), .Y(n1602) );
  oa211d1_hd U807 ( .A(a_m[11]), .B(n1602), .C(n1601), .D(n1600), .Y(n1604) );
  oa22d1_hd U808 ( .A(a_m[13]), .B(n2017), .C(a_m[14]), .D(n2015), .Y(n1603)
         );
  ao21d1_hd U809 ( .A(n1605), .B(n1604), .C(n1603), .Y(n1606) );
  ao211d1_hd U810 ( .A(a_m[14]), .B(n2015), .C(n1607), .D(n1606), .Y(n1609) );
  oa22d1_hd U811 ( .A(a_m[16]), .B(n2011), .C(a_m[15]), .D(n2013), .Y(n1608)
         );
  oa22d1_hd U812 ( .A(n1609), .B(n1608), .C(b_m[16]), .D(n2059), .Y(n1610) );
  ao22d1_hd U813 ( .A(a_m[17]), .B(n2009), .C(n1611), .D(n1610), .Y(n1612) );
  nr2d1_hd U814 ( .A(b_m[18]), .B(n1612), .Y(n1615) );
  oa211d1_hd U815 ( .A(a_m[18]), .B(n1615), .C(n1614), .D(n1613), .Y(n1616) );
  ao22d1_hd U816 ( .A(b_m[20]), .B(n2051), .C(n1617), .D(n1616), .Y(n1618) );
  ao22d1_hd U817 ( .A(b_m[22]), .B(n2047), .C(n1620), .D(n1619), .Y(n1621) );
  oa22d1_hd U818 ( .A(a_m[23]), .B(n1997), .C(a_m[24]), .D(n1995), .Y(n1623)
         );
  ao22d1_hd U819 ( .A(a_m[24]), .B(n1995), .C(a_m[25]), .D(n1629), .Y(n1622)
         );
  ivd1_hd U820 ( .A(a_m[0]), .Y(n2089) );
  ao22d1_hd U821 ( .A(n1568), .B(n2041), .C(n2089), .D(n1569), .Y(C2_Z_0) );
  ao22d1_hd U822 ( .A(n1568), .B(n2040), .C(n2088), .D(n1569), .Y(C2_Z_1) );
  ao22d1_hd U823 ( .A(n1568), .B(n2023), .C(n2071), .D(n1569), .Y(C2_Z_10) );
  ao22d1_hd U824 ( .A(n1568), .B(n2021), .C(n2069), .D(n1569), .Y(C2_Z_11) );
  ao22d1_hd U825 ( .A(n1568), .B(n2019), .C(n2067), .D(n1569), .Y(C2_Z_12) );
  ao22d1_hd U826 ( .A(n1568), .B(n2017), .C(n2065), .D(n1569), .Y(C2_Z_13) );
  ao22d1_hd U827 ( .A(n1568), .B(n2015), .C(n2063), .D(n1569), .Y(C2_Z_14) );
  ao22d1_hd U828 ( .A(n1568), .B(n2013), .C(n2061), .D(n1569), .Y(C2_Z_15) );
  ao22d1_hd U829 ( .A(n1568), .B(n2011), .C(n2059), .D(n1569), .Y(C2_Z_16) );
  ao22d1_hd U830 ( .A(n1568), .B(n2009), .C(n2057), .D(n1569), .Y(C2_Z_17) );
  ao22d1_hd U831 ( .A(n1568), .B(n2007), .C(n2055), .D(n1569), .Y(C2_Z_18) );
  ao22d1_hd U832 ( .A(n1568), .B(n2005), .C(n2053), .D(n1569), .Y(C2_Z_19) );
  ao22d1_hd U833 ( .A(n1568), .B(n2039), .C(n2087), .D(n1569), .Y(C2_Z_2) );
  ao22d1_hd U834 ( .A(n1568), .B(n2003), .C(n2051), .D(n1569), .Y(C2_Z_20) );
  ao22d1_hd U835 ( .A(n1568), .B(n2001), .C(n2049), .D(n1569), .Y(C2_Z_21) );
  ao22d1_hd U836 ( .A(n1568), .B(n1999), .C(n2047), .D(n1569), .Y(C2_Z_22) );
  ao22d1_hd U837 ( .A(n1568), .B(n1997), .C(n2045), .D(n1569), .Y(C2_Z_23) );
  ao22d1_hd U838 ( .A(n1568), .B(n1995), .C(n2043), .D(n1569), .Y(C2_Z_24) );
  ao22d1_hd U839 ( .A(n1568), .B(n1629), .C(n1668), .D(n1569), .Y(C2_Z_25) );
  oa21d1_hd U840 ( .A(n2250), .B(n1791), .C(n2092), .Y(C2_Z_26) );
  ao22d1_hd U841 ( .A(n1568), .B(n2038), .C(n2086), .D(n1569), .Y(C2_Z_3) );
  ao22d1_hd U842 ( .A(n1568), .B(n2035), .C(n2083), .D(n1569), .Y(C2_Z_4) );
  ao22d1_hd U843 ( .A(n1568), .B(n2033), .C(n2081), .D(n1569), .Y(C2_Z_5) );
  ao22d1_hd U844 ( .A(n1568), .B(n2031), .C(n2079), .D(n1569), .Y(C2_Z_6) );
  ao22d1_hd U845 ( .A(n1568), .B(n2029), .C(n2077), .D(n1569), .Y(C2_Z_7) );
  ao22d1_hd U846 ( .A(n1568), .B(n2027), .C(n2075), .D(n1569), .Y(C2_Z_8) );
  ao22d1_hd U847 ( .A(n1568), .B(n2025), .C(n2073), .D(n1569), .Y(C2_Z_9) );
  nr2d1_hd U848 ( .A(n2250), .B(n2092), .Y(n1628) );
  ao22d1_hd U849 ( .A(n2265), .B(n1628), .C(n2250), .D(n1791), .Y(
        DP_OP_43J4_124_6938_n32) );
  ao22d1_hd U850 ( .A(b_m[25]), .B(n1791), .C(n1655), .D(n1629), .Y(n1630) );
  oa21d1_hd U851 ( .A(a_m[25]), .B(n1569), .C(n1630), .Y(
        DP_OP_43J4_124_6938_n33) );
  ao22d1_hd U852 ( .A(b_m[24]), .B(n1791), .C(n1655), .D(n1995), .Y(n1631) );
  oa21d1_hd U853 ( .A(a_m[24]), .B(n1569), .C(n1631), .Y(
        DP_OP_43J4_124_6938_n34) );
  ao22d1_hd U854 ( .A(b_m[23]), .B(n1791), .C(n1655), .D(n1997), .Y(n1632) );
  oa21d1_hd U855 ( .A(a_m[23]), .B(n1569), .C(n1632), .Y(
        DP_OP_43J4_124_6938_n35) );
  ao22d1_hd U856 ( .A(n1568), .B(n2047), .C(n1655), .D(n1999), .Y(n1633) );
  oa21d1_hd U857 ( .A(n2265), .B(n1999), .C(n1633), .Y(DP_OP_43J4_124_6938_n36) );
  ao22d1_hd U858 ( .A(b_m[21]), .B(n1791), .C(n1655), .D(n2001), .Y(n1634) );
  oa21d1_hd U859 ( .A(a_m[21]), .B(n1569), .C(n1634), .Y(
        DP_OP_43J4_124_6938_n37) );
  ao22d1_hd U860 ( .A(n1568), .B(n2051), .C(n1655), .D(n2003), .Y(n1635) );
  oa21d1_hd U861 ( .A(n2265), .B(n2003), .C(n1635), .Y(DP_OP_43J4_124_6938_n38) );
  ao22d1_hd U862 ( .A(n1568), .B(n2053), .C(n1655), .D(n2005), .Y(n1636) );
  oa21d1_hd U863 ( .A(n2265), .B(n2005), .C(n1636), .Y(DP_OP_43J4_124_6938_n39) );
  ao22d1_hd U864 ( .A(b_m[18]), .B(n1791), .C(n1655), .D(n2007), .Y(n1637) );
  oa21d1_hd U865 ( .A(a_m[18]), .B(n1569), .C(n1637), .Y(
        DP_OP_43J4_124_6938_n40) );
  ao22d1_hd U866 ( .A(n1568), .B(n2057), .C(n1655), .D(n2009), .Y(n1638) );
  oa21d1_hd U867 ( .A(n2265), .B(n2009), .C(n1638), .Y(DP_OP_43J4_124_6938_n41) );
  ao22d1_hd U868 ( .A(n1568), .B(n2059), .C(n1655), .D(n2011), .Y(n1639) );
  oa21d1_hd U869 ( .A(n2265), .B(n2011), .C(n1639), .Y(DP_OP_43J4_124_6938_n42) );
  ao22d1_hd U870 ( .A(n1568), .B(n2061), .C(n1655), .D(n2013), .Y(n1640) );
  oa21d1_hd U871 ( .A(n2265), .B(n2013), .C(n1640), .Y(DP_OP_43J4_124_6938_n43) );
  ao22d1_hd U872 ( .A(b_m[14]), .B(n1791), .C(n1655), .D(n2015), .Y(n1641) );
  oa21d1_hd U873 ( .A(a_m[14]), .B(n1569), .C(n1641), .Y(
        DP_OP_43J4_124_6938_n44) );
  ao22d1_hd U874 ( .A(b_m[13]), .B(n1791), .C(n1655), .D(n2017), .Y(n1642) );
  oa21d1_hd U875 ( .A(a_m[13]), .B(n1569), .C(n1642), .Y(
        DP_OP_43J4_124_6938_n45) );
  ao22d1_hd U876 ( .A(n1568), .B(n2067), .C(n1655), .D(n2019), .Y(n1643) );
  oa21d1_hd U877 ( .A(n2265), .B(n2019), .C(n1643), .Y(DP_OP_43J4_124_6938_n46) );
  ao22d1_hd U878 ( .A(b_m[11]), .B(n1791), .C(n1655), .D(n2021), .Y(n1644) );
  oa21d1_hd U879 ( .A(a_m[11]), .B(n1569), .C(n1644), .Y(
        DP_OP_43J4_124_6938_n47) );
  ao22d1_hd U880 ( .A(n1568), .B(n2071), .C(n1655), .D(n2023), .Y(n1645) );
  oa21d1_hd U881 ( .A(n2265), .B(n2023), .C(n1645), .Y(DP_OP_43J4_124_6938_n48) );
  ao22d1_hd U882 ( .A(n1568), .B(n2073), .C(n1655), .D(n2025), .Y(n1646) );
  oa21d1_hd U883 ( .A(n2265), .B(n2025), .C(n1646), .Y(DP_OP_43J4_124_6938_n49) );
  ao22d1_hd U884 ( .A(n1568), .B(n2075), .C(n1655), .D(n2027), .Y(n1647) );
  oa21d1_hd U885 ( .A(n2265), .B(n2027), .C(n1647), .Y(DP_OP_43J4_124_6938_n50) );
  ao22d1_hd U886 ( .A(b_m[7]), .B(n1791), .C(n1655), .D(n2029), .Y(n1648) );
  oa21d1_hd U887 ( .A(a_m[7]), .B(n1569), .C(n1648), .Y(
        DP_OP_43J4_124_6938_n51) );
  ao22d1_hd U888 ( .A(b_m[6]), .B(n1791), .C(n1655), .D(n2031), .Y(n1649) );
  oa21d1_hd U889 ( .A(a_m[6]), .B(n1569), .C(n1649), .Y(
        DP_OP_43J4_124_6938_n52) );
  ao22d1_hd U890 ( .A(n1568), .B(n2081), .C(n1655), .D(n2033), .Y(n1650) );
  oa21d1_hd U891 ( .A(n2265), .B(n2033), .C(n1650), .Y(DP_OP_43J4_124_6938_n53) );
  ao22d1_hd U892 ( .A(n1568), .B(n2083), .C(n1655), .D(n2035), .Y(n1651) );
  oa21d1_hd U893 ( .A(n2265), .B(n2035), .C(n1651), .Y(DP_OP_43J4_124_6938_n54) );
  ao22d1_hd U894 ( .A(n1568), .B(n2086), .C(n1655), .D(n2038), .Y(n1652) );
  oa21d1_hd U895 ( .A(n2265), .B(n2038), .C(n1652), .Y(DP_OP_43J4_124_6938_n55) );
  ao22d1_hd U896 ( .A(b_m[2]), .B(n1791), .C(n1655), .D(n2039), .Y(n1653) );
  oa21d1_hd U897 ( .A(a_m[2]), .B(n1569), .C(n1653), .Y(
        DP_OP_43J4_124_6938_n56) );
  ao22d1_hd U898 ( .A(b_m[1]), .B(n1791), .C(n1655), .D(n2040), .Y(n1654) );
  oa21d1_hd U899 ( .A(a_m[1]), .B(n1569), .C(n1654), .Y(
        DP_OP_43J4_124_6938_n57) );
  ao22d1_hd U900 ( .A(b_m[0]), .B(n1791), .C(n1655), .D(n2041), .Y(n1656) );
  oa21d1_hd U901 ( .A(a_m[0]), .B(n1569), .C(n1656), .Y(
        DP_OP_43J4_124_6938_n58) );
  ao22d1_hd U902 ( .A(n1568), .B(n1657), .C(n1709), .D(n1569), .Y(N338) );
  nr4d1_hd U903 ( .A(a_e[1]), .B(a_e[2]), .C(a_e[3]), .D(a_e[4]), .Y(n1658) );
  nd4d1_hd U904 ( .A(a_e[7]), .B(n1658), .C(n2097), .D(n2116), .Y(n1678) );
  nr4d1_hd U905 ( .A(n1678), .B(n2144), .C(n1698), .D(n2099), .Y(n2094) );
  nr4d1_hd U906 ( .A(b_e[2]), .B(b_e[1]), .C(b_e[3]), .D(b_e[4]), .Y(n1659) );
  nd4d1_hd U907 ( .A(b_e[7]), .B(n1659), .C(n2184), .D(n2164), .Y(n1677) );
  nr4d1_hd U908 ( .A(n2166), .B(n1677), .C(n2211), .D(n1683), .Y(n2160) );
  nd4d1_hd U909 ( .A(n2033), .B(n2035), .C(n2025), .D(n2013), .Y(n1667) );
  nr4d1_hd U910 ( .A(b_m[0]), .B(b_m[1]), .C(b_m[2]), .D(b_m[3]), .Y(n1660) );
  nd4d1_hd U911 ( .A(n1660), .B(n2011), .C(n2031), .D(n2017), .Y(n1666) );
  nr4d1_hd U912 ( .A(b_m[25]), .B(b_m[23]), .C(b_m[22]), .D(b_m[26]), .Y(n1664) );
  nr4d1_hd U913 ( .A(b_m[18]), .B(b_m[11]), .C(b_m[14]), .D(b_m[24]), .Y(n1663) );
  nr4d1_hd U914 ( .A(b_m[8]), .B(b_m[7]), .C(b_m[10]), .D(b_m[12]), .Y(n1662)
         );
  nr4d1_hd U915 ( .A(b_m[17]), .B(b_m[19]), .C(b_m[20]), .D(b_m[21]), .Y(n1661) );
  nd4d1_hd U916 ( .A(n1664), .B(n1663), .C(n1662), .D(n1661), .Y(n1665) );
  nr3d1_hd U917 ( .A(n1667), .B(n1666), .C(n1665), .Y(n1711) );
  nd4d1_hd U918 ( .A(n2057), .B(n2075), .C(n2049), .D(n2043), .Y(n1676) );
  nr4d1_hd U919 ( .A(a_m[18]), .B(a_m[12]), .C(a_m[20]), .D(a_m[26]), .Y(n1669) );
  nd4d1_hd U920 ( .A(n1669), .B(n2045), .C(n2047), .D(n1668), .Y(n1675) );
  nr4d1_hd U921 ( .A(a_m[11]), .B(a_m[6]), .C(a_m[9]), .D(a_m[10]), .Y(n1673)
         );
  nr4d1_hd U922 ( .A(a_m[13]), .B(a_m[14]), .C(a_m[15]), .D(a_m[19]), .Y(n1672) );
  nr4d1_hd U923 ( .A(a_m[16]), .B(a_m[5]), .C(a_m[4]), .D(a_m[7]), .Y(n1671)
         );
  nr4d1_hd U924 ( .A(a_m[0]), .B(a_m[1]), .C(a_m[2]), .D(a_m[3]), .Y(n1670) );
  nd4d1_hd U925 ( .A(n1673), .B(n1672), .C(n1671), .D(n1670), .Y(n1674) );
  nr4d1_hd U926 ( .A(b_e[8]), .B(b_e[0]), .C(b_e[9]), .D(n1677), .Y(n1710) );
  nr2d1_hd U927 ( .A(n1710), .B(n2223), .Y(n1750) );
  ao22d1_hd U928 ( .A(b_e[2]), .B(n2137), .C(b_e[3]), .D(n2128), .Y(n1685) );
  nr2d1_hd U929 ( .A(a_e[1]), .B(n2212), .Y(n1681) );
  ao22d1_hd U930 ( .A(b_e[4]), .B(n2121), .C(b_e[5]), .D(n2116), .Y(n1680) );
  ao211d1_hd U931 ( .A(b_e[0]), .B(n2144), .C(n1681), .D(n1688), .Y(n1682) );
  oa211d1_hd U932 ( .A(a_e[7]), .B(n2168), .C(n1685), .D(n1682), .Y(n1684) );
  nd3bd1_hd U933 ( .AN(n1684), .B(n1697), .C(n1700), .Y(n2233) );
  ao211d1_hd U934 ( .A(b_e[6]), .B(n2097), .C(b_e[5]), .D(n2116), .Y(n1692) );
  ivd1_hd U935 ( .A(b_e[4]), .Y(n2190) );
  ivd1_hd U936 ( .A(b_e[3]), .Y(n2161) );
  ao22d1_hd U937 ( .A(a_e[4]), .B(n2190), .C(a_e[3]), .D(n2161), .Y(n1690) );
  ao211d1_hd U938 ( .A(b_e[1]), .B(n2145), .C(b_e[0]), .D(n2144), .Y(n1687) );
  oa22d1_hd U939 ( .A(b_e[1]), .B(n2145), .C(b_e[2]), .D(n2137), .Y(n1686) );
  oa21d1_hd U940 ( .A(n1687), .B(n1686), .C(n1685), .Y(n1689) );
  ao21d1_hd U941 ( .A(n1690), .B(n1689), .C(n1688), .Y(n1691) );
  ao211d1_hd U942 ( .A(a_e[6]), .B(n2164), .C(n1692), .D(n1691), .Y(n1695) );
  scg6d1_hd U943 ( .A(b_e[7]), .B(n1695), .C(n2101), .Y(n1693) );
  oa211d1_hd U944 ( .A(b_e[7]), .B(n1695), .C(n1694), .D(n1693), .Y(n1696) );
  oa21d1_hd U945 ( .A(n2094), .B(n2242), .C(n1575), .Y(n1) );
  oa21d1_hd U946 ( .A(n2160), .B(n2242), .C(n2158), .Y(n2) );
  nr2d1_hd U947 ( .A(n1733), .B(n1975), .Y(n1703) );
  nr4d1_hd U948 ( .A(z_e[2]), .B(z_e[3]), .C(z_e[4]), .D(z_e[5]), .Y(n1702) );
  ivd1_hd U949 ( .A(z_e[6]), .Y(n1745) );
  nd3d1_hd U950 ( .A(z_e[9]), .B(n1702), .C(n1745), .Y(n1728) );
  ivd1_hd U951 ( .A(z_e[9]), .Y(n1987) );
  ao21d1_hd U952 ( .A(n1703), .B(n1728), .C(n1987), .Y(n1705) );
  nr2d1_hd U953 ( .A(n2256), .B(n2228), .Y(n1806) );
  nr2d1_hd U954 ( .A(n1727), .B(n1985), .Y(n1704) );
  scg16d1_hd U955 ( .A(n1705), .B(n1704), .C(n1964), .Y(n2227) );
  nr2d1_hd U956 ( .A(n2227), .B(n1988), .Y(n1706) );
  nr2d1_hd U957 ( .A(n1806), .B(n1706), .Y(n1970) );
  ivd1_hd U958 ( .A(n2256), .Y(n2229) );
  scg4d1_hd U959 ( .A(n2229), .B(z_m[0]), .C(n2266), .D(round_bit), .E(n1573), 
        .F(sum[2]), .G(sum[3]), .H(n1943), .Y(n266) );
  nr2d1_hd U960 ( .A(n1707), .B(n2243), .Y(n2220) );
  nr2d1_hd U961 ( .A(a_s), .B(n1717), .Y(n1708) );
  oa21d1_hd U962 ( .A(n1715), .B(n1708), .C(n1793), .Y(n1714) );
  nr3d1_hd U963 ( .A(n1710), .B(n1792), .C(n1709), .Y(n1713) );
  oa22d1_hd U964 ( .A(n1712), .B(n1792), .C(n1711), .D(n1793), .Y(n1794) );
  ao211d1_hd U965 ( .A(b_s), .B(n1714), .C(n1713), .D(n1794), .Y(n1732) );
  ao21d1_hd U966 ( .A(n1792), .B(n1793), .C(n2223), .Y(n1734) );
  ao211d1_hd U967 ( .A(n2267), .B(n1719), .C(n1734), .D(n1796), .Y(n2257) );
  ao22d1_hd U968 ( .A(a_s), .B(n1572), .C(n1577), .D(z[31]), .Y(n1731) );
  ivd1_hd U969 ( .A(z_m[4]), .Y(n1916) );
  ivd1_hd U970 ( .A(z_m[3]), .Y(n1924) );
  nd4d1_hd U971 ( .A(n1946), .B(n1916), .C(n1924), .D(n1910), .Y(n1720) );
  nr4d1_hd U972 ( .A(z_m[0]), .B(z_m[19]), .C(z_m[2]), .D(n1720), .Y(n1726) );
  ivd1_hd U973 ( .A(z_m[12]), .Y(n1868) );
  ivd1_hd U974 ( .A(z_m[11]), .Y(n1875) );
  nd4d1_hd U975 ( .A(n1886), .B(n1868), .C(n1875), .D(n1862), .Y(n1724) );
  ivd1_hd U976 ( .A(z_m[8]), .Y(n1892) );
  ivd1_hd U977 ( .A(z_m[7]), .Y(n1899) );
  nd4d1_hd U978 ( .A(n1923), .B(n1892), .C(n1899), .D(n1898), .Y(n1723) );
  nd4d1_hd U979 ( .A(n1965), .B(n1826), .C(n1832), .D(n1850), .Y(n1722) );
  ivd1_hd U980 ( .A(z_m[16]), .Y(n1844) );
  ivd1_hd U981 ( .A(z_m[15]), .Y(n1851) );
  nd4d1_hd U982 ( .A(n1874), .B(n1844), .C(n1851), .D(n1838), .Y(n1721) );
  nr4d1_hd U983 ( .A(n1724), .B(n1723), .C(n1722), .D(n1721), .Y(n1725) );
  oa211d1_hd U984 ( .A(n1729), .B(n1735), .C(n1796), .D(z_s), .Y(n1730) );
  oa211d1_hd U985 ( .A(n1732), .B(n2223), .C(n1731), .D(n1730), .Y(n361) );
  ao21d1_hd U986 ( .A(n1733), .B(n1975), .C(z_e[9]), .Y(n1797) );
  nr2d1_hd U987 ( .A(z_e[1]), .B(z_e[0]), .Y(n1778) );
  ivd1_hd U988 ( .A(z_e[2]), .Y(n1773) );
  nr2d1_hd U989 ( .A(z_e[3]), .B(n1772), .Y(n1764) );
  ivd1_hd U990 ( .A(z_e[4]), .Y(n1760) );
  nr2d1_hd U991 ( .A(z_e[5]), .B(n1759), .Y(n1749) );
  nr2d1_hd U992 ( .A(z_e[7]), .B(n1744), .Y(n1736) );
  ao211d1_hd U993 ( .A(z_e[7]), .B(n1744), .C(n1790), .D(n1736), .Y(n1740) );
  nd3d1_hd U994 ( .A(n2212), .B(n2145), .C(n1786), .Y(n1780) );
  nr2d1_hd U995 ( .A(n1780), .B(n1771), .Y(n1770) );
  nd3d1_hd U996 ( .A(n1770), .B(n2161), .C(n2128), .Y(n1765) );
  nr2d1_hd U997 ( .A(n1765), .B(n1758), .Y(n1757) );
  nd3d1_hd U998 ( .A(n1757), .B(n2184), .C(n2116), .Y(n1752) );
  nr2d1_hd U999 ( .A(n1752), .B(n1743), .Y(n1742) );
  nr2d1_hd U1000 ( .A(n1742), .B(n1738), .Y(n1737) );
  ao211d1_hd U1001 ( .A(n1742), .B(n1738), .C(n1800), .D(n1737), .Y(n1739) );
  ao211d1_hd U1002 ( .A(n1577), .B(z[30]), .C(n1740), .D(n1739), .Y(n1741) );
  ao21d1_hd U1003 ( .A(n1752), .B(n1743), .C(n1742), .Y(n1748) );
  ivd1_hd U1004 ( .A(n1790), .Y(n1775) );
  oa21d1_hd U1005 ( .A(n1749), .B(n1745), .C(n1744), .Y(n1746) );
  ao22d1_hd U1006 ( .A(n1577), .B(z[29]), .C(n1775), .D(n1746), .Y(n1747) );
  oa211d1_hd U1007 ( .A(n1748), .B(n1800), .C(n1789), .D(n1747), .Y(n363) );
  ao21d1_hd U1008 ( .A(z_e[5]), .B(n1759), .C(n1749), .Y(n1756) );
  ao22d1_hd U1009 ( .A(b_e[5]), .B(n1804), .C(a_e[5]), .D(n1787), .Y(n1753) );
  oa22d1_hd U1010 ( .A(n1757), .B(n1753), .C(n1800), .D(n1752), .Y(n1754) );
  ao21d1_hd U1011 ( .A(n1577), .B(z[28]), .C(n1754), .Y(n1755) );
  oa211d1_hd U1012 ( .A(n1756), .B(n1790), .C(n1789), .D(n1755), .Y(n364) );
  ao21d1_hd U1013 ( .A(n1765), .B(n1758), .C(n1757), .Y(n1763) );
  oa21d1_hd U1014 ( .A(n1764), .B(n1760), .C(n1759), .Y(n1761) );
  ao22d1_hd U1015 ( .A(n1577), .B(z[27]), .C(n1775), .D(n1761), .Y(n1762) );
  oa211d1_hd U1016 ( .A(n1763), .B(n1800), .C(n1789), .D(n1762), .Y(n365) );
  ao21d1_hd U1017 ( .A(z_e[3]), .B(n1772), .C(n1764), .Y(n1769) );
  ao22d1_hd U1018 ( .A(b_e[3]), .B(n1804), .C(a_e[3]), .D(n1787), .Y(n1766) );
  oa22d1_hd U1019 ( .A(n1770), .B(n1766), .C(n1800), .D(n1765), .Y(n1767) );
  ao21d1_hd U1020 ( .A(n1577), .B(z[26]), .C(n1767), .Y(n1768) );
  oa211d1_hd U1021 ( .A(n1769), .B(n1790), .C(n1789), .D(n1768), .Y(n366) );
  ao21d1_hd U1022 ( .A(n1780), .B(n1771), .C(n1770), .Y(n1777) );
  oa21d1_hd U1023 ( .A(n1778), .B(n1773), .C(n1772), .Y(n1774) );
  ao22d1_hd U1024 ( .A(n1577), .B(z[25]), .C(n1775), .D(n1774), .Y(n1776) );
  oa211d1_hd U1025 ( .A(n1777), .B(n1800), .C(n1789), .D(n1776), .Y(n367) );
  ao21d1_hd U1026 ( .A(z_e[0]), .B(z_e[1]), .C(n1778), .Y(n1785) );
  nr3d1_hd U1027 ( .A(n2212), .B(n1786), .C(n1779), .Y(n1783) );
  nd2bd1_hd U1028 ( .AN(n1786), .B(a_e[1]), .Y(n1781) );
  ao21d1_hd U1029 ( .A(n1781), .B(n1780), .C(n1800), .Y(n1782) );
  ao211d1_hd U1030 ( .A(n1577), .B(z[24]), .C(n1783), .D(n1782), .Y(n1784) );
  oa211d1_hd U1031 ( .A(n1785), .B(n1790), .C(n1789), .D(n1784), .Y(n368) );
  ao22d1_hd U1032 ( .A(n1577), .B(z[23]), .C(n1787), .D(n1786), .Y(n1788) );
  oa211d1_hd U1033 ( .A(z_e[0]), .B(n1790), .C(n1789), .D(n1788), .Y(n369) );
  nr3d1_hd U1034 ( .A(n1793), .B(n1792), .C(n1791), .Y(n1795) );
  nr2d1_hd U1035 ( .A(n1795), .B(n1794), .Y(n1801) );
  ao22d1_hd U1036 ( .A(b_m[25]), .B(n1804), .C(z_m[22]), .D(n1803), .Y(n1799)
         );
  ao22d1_hd U1037 ( .A(a_m[25]), .B(n1572), .C(n1577), .D(z[22]), .Y(n1798) );
  oa211d1_hd U1038 ( .A(n1801), .B(n1800), .C(n1799), .D(n1798), .Y(n370) );
  scg4d1_hd U1039 ( .A(b_m[24]), .B(n1804), .C(z_m[21]), .D(n1803), .E(a_m[24]), .F(n1572), .G(n1577), .H(z[21]), .Y(n371) );
  scg4d1_hd U1040 ( .A(b_m[23]), .B(n1804), .C(z_m[20]), .D(n1803), .E(a_m[23]), .F(n1572), .G(n1577), .H(z[20]), .Y(n372) );
  scg4d1_hd U1041 ( .A(b_m[22]), .B(n1804), .C(z_m[19]), .D(n1803), .E(a_m[22]), .F(n1572), .G(n1577), .H(z[19]), .Y(n373) );
  scg4d1_hd U1042 ( .A(b_m[21]), .B(n1804), .C(z_m[18]), .D(n1803), .E(a_m[21]), .F(n1572), .G(n1577), .H(z[18]), .Y(n374) );
  scg4d1_hd U1043 ( .A(b_m[20]), .B(n1804), .C(z_m[17]), .D(n1803), .E(a_m[20]), .F(n1572), .G(n1577), .H(z[17]), .Y(n375) );
  scg4d1_hd U1044 ( .A(b_m[19]), .B(n1804), .C(z_m[16]), .D(n1803), .E(a_m[19]), .F(n1572), .G(n1577), .H(z[16]), .Y(n376) );
  scg4d1_hd U1045 ( .A(b_m[18]), .B(n1804), .C(z_m[15]), .D(n1803), .E(a_m[18]), .F(n1572), .G(n1577), .H(z[15]), .Y(n377) );
  scg4d1_hd U1046 ( .A(b_m[17]), .B(n1804), .C(z_m[14]), .D(n1803), .E(a_m[17]), .F(n1572), .G(n1577), .H(z[14]), .Y(n378) );
  scg4d1_hd U1047 ( .A(b_m[16]), .B(n1804), .C(z_m[13]), .D(n1803), .E(a_m[16]), .F(n1572), .G(n1577), .H(z[13]), .Y(n379) );
  scg4d1_hd U1048 ( .A(b_m[15]), .B(n1804), .C(z_m[12]), .D(n1803), .E(a_m[15]), .F(n1572), .G(n1577), .H(z[12]), .Y(n380) );
  scg4d1_hd U1049 ( .A(b_m[14]), .B(n1804), .C(z_m[11]), .D(n1803), .E(a_m[14]), .F(n1802), .G(n1577), .H(z[11]), .Y(n381) );
  scg4d1_hd U1050 ( .A(b_m[13]), .B(n1804), .C(z_m[10]), .D(n1803), .E(a_m[13]), .F(n1802), .G(n1577), .H(z[10]), .Y(n382) );
  scg4d1_hd U1051 ( .A(b_m[12]), .B(n1804), .C(z_m[9]), .D(n1803), .E(a_m[12]), 
        .F(n1802), .G(n1577), .H(z[9]), .Y(n383) );
  scg4d1_hd U1052 ( .A(b_m[11]), .B(n1804), .C(z_m[8]), .D(n1803), .E(a_m[11]), 
        .F(n1802), .G(n1577), .H(z[8]), .Y(n384) );
  scg4d1_hd U1053 ( .A(b_m[10]), .B(n1804), .C(z_m[7]), .D(n1803), .E(a_m[10]), 
        .F(n1802), .G(n1577), .H(z[7]), .Y(n385) );
  scg4d1_hd U1054 ( .A(b_m[9]), .B(n1804), .C(z_m[6]), .D(n1803), .E(a_m[9]), 
        .F(n1802), .G(n1577), .H(z[6]), .Y(n386) );
  scg4d1_hd U1055 ( .A(b_m[8]), .B(n1804), .C(z_m[5]), .D(n1803), .E(a_m[8]), 
        .F(n1572), .G(n1577), .H(z[5]), .Y(n387) );
  scg4d1_hd U1056 ( .A(b_m[7]), .B(n1804), .C(z_m[4]), .D(n1803), .E(a_m[7]), 
        .F(n1572), .G(n2257), .H(z[4]), .Y(n388) );
  scg4d1_hd U1057 ( .A(b_m[6]), .B(n1804), .C(z_m[3]), .D(n1803), .E(a_m[6]), 
        .F(n1572), .G(n1577), .H(z[3]), .Y(n389) );
  scg4d1_hd U1058 ( .A(b_m[5]), .B(n1804), .C(z_m[2]), .D(n1803), .E(a_m[5]), 
        .F(n1572), .G(n1577), .H(z[2]), .Y(n390) );
  scg4d1_hd U1059 ( .A(b_m[4]), .B(n1804), .C(z_m[1]), .D(n1803), .E(a_m[4]), 
        .F(n1572), .G(n1577), .H(z[1]), .Y(n391) );
  scg4d1_hd U1060 ( .A(b_m[3]), .B(n1804), .C(z_m[0]), .D(n1803), .E(a_m[3]), 
        .F(n1802), .G(n1577), .H(z[0]), .Y(n392) );
  ao22d1_hd U1061 ( .A(n1972), .B(sum[0]), .C(sticky), .D(n1805), .Y(n1808) );
  ao22d1_hd U1062 ( .A(n1806), .B(round_bit), .C(n1943), .D(sum[1]), .Y(n1807)
         );
  ivd1_hd U1063 ( .A(round_bit), .Y(n1811) );
  ao22d1_hd U1064 ( .A(n1573), .B(sum[1]), .C(n1943), .D(sum[2]), .Y(n1810) );
  nd3d1_hd U1065 ( .A(n2229), .B(guard), .C(n265), .Y(n1809) );
  oa211d1_hd U1066 ( .A(n1811), .B(n265), .C(n1810), .D(n1809), .Y(n394) );
  nr3d1_hd U1067 ( .A(z_m[0]), .B(sticky), .C(round_bit), .Y(n1812) );
  ao22d1_hd U1068 ( .A(n1573), .B(sum[25]), .C(n1943), .D(sum[26]), .Y(n1816)
         );
  nd3d1_hd U1069 ( .A(z_m[0]), .B(z_m[2]), .C(z_m[1]), .Y(n1917) );
  ivd1_hd U1070 ( .A(n1917), .Y(n1918) );
  nd3d1_hd U1071 ( .A(n1918), .B(z_m[4]), .C(z_m[3]), .Y(n1905) );
  nr3d1_hd U1072 ( .A(n1905), .B(n1910), .C(n1923), .Y(n1893) );
  nd3d1_hd U1073 ( .A(n1893), .B(z_m[8]), .C(z_m[7]), .Y(n1881) );
  nr3d1_hd U1074 ( .A(n1881), .B(n1898), .C(n1886), .Y(n1869) );
  nd3d1_hd U1075 ( .A(n1869), .B(z_m[12]), .C(z_m[11]), .Y(n1857) );
  nr3d1_hd U1076 ( .A(n1857), .B(n1862), .C(n1874), .Y(n1845) );
  nd3d1_hd U1077 ( .A(n1845), .B(z_m[16]), .C(z_m[15]), .Y(n1833) );
  nr3d1_hd U1078 ( .A(n1833), .B(n1838), .C(n1850), .Y(n1967) );
  oa21d1_hd U1079 ( .A(n1967), .B(n2258), .C(n1952), .Y(n1829) );
  ao21d1_hd U1080 ( .A(n1971), .B(n1813), .C(n1829), .Y(n1817) );
  oa21d1_hd U1081 ( .A(z_m[21]), .B(n1931), .C(n1817), .Y(n1954) );
  ivd1_hd U1082 ( .A(z_m[19]), .Y(n1962) );
  nr2d1_hd U1083 ( .A(n1962), .B(n1827), .Y(n1823) );
  oa21d1_hd U1084 ( .A(z_m[22]), .B(n1958), .C(n1956), .Y(n1814) );
  ao22d1_hd U1085 ( .A(z_m[22]), .B(n1954), .C(z_m[21]), .D(n1814), .Y(n1815)
         );
  oa211d1_hd U1086 ( .A(n1964), .B(n1945), .C(n1816), .D(n1815), .Y(n395) );
  ao22d1_hd U1087 ( .A(n1573), .B(sum[24]), .C(sum[25]), .D(n1943), .Y(n1820)
         );
  ao22d1_hd U1088 ( .A(z_m[21]), .B(n1817), .C(n1958), .D(n1826), .Y(n1818) );
  ao21d1_hd U1089 ( .A(z_m[20]), .B(n1949), .C(n1818), .Y(n1819) );
  oa211d1_hd U1090 ( .A(n1965), .B(n1945), .C(n1820), .D(n1819), .Y(n396) );
  ao22d1_hd U1091 ( .A(n1573), .B(sum[23]), .C(n1943), .D(sum[24]), .Y(n1825)
         );
  ao21d1_hd U1092 ( .A(n1955), .B(n1962), .C(n1829), .Y(n1821) );
  oa22d1_hd U1093 ( .A(n1821), .B(n1832), .C(n1962), .D(n1956), .Y(n1822) );
  ao21d1_hd U1094 ( .A(n1823), .B(n1832), .C(n1822), .Y(n1824) );
  oa211d1_hd U1095 ( .A(n1826), .B(n1945), .C(n1825), .D(n1824), .Y(n397) );
  ao22d1_hd U1096 ( .A(n1573), .B(sum[22]), .C(n1943), .D(sum[23]), .Y(n1831)
         );
  oa22d1_hd U1097 ( .A(z_m[19]), .B(n1827), .C(n1956), .D(n1838), .Y(n1828) );
  ao21d1_hd U1098 ( .A(z_m[19]), .B(n1829), .C(n1828), .Y(n1830) );
  oa211d1_hd U1099 ( .A(n1832), .B(n1945), .C(n1831), .D(n1830), .Y(n398) );
  nr2d1_hd U1100 ( .A(n1931), .B(n1833), .Y(n1841) );
  ao21d1_hd U1101 ( .A(n1841), .B(n1838), .C(n1949), .Y(n1837) );
  ao22d1_hd U1102 ( .A(n1573), .B(sum[21]), .C(n1943), .D(sum[22]), .Y(n1836)
         );
  ao21d1_hd U1103 ( .A(n1971), .B(n1833), .C(n1932), .Y(n1839) );
  oa21d1_hd U1104 ( .A(z_m[17]), .B(n1931), .C(n1839), .Y(n1834) );
  ao22d1_hd U1105 ( .A(z_m[19]), .B(n1938), .C(z_m[18]), .D(n1834), .Y(n1835)
         );
  oa211d1_hd U1106 ( .A(n1837), .B(n1850), .C(n1836), .D(n1835), .Y(n399) );
  ao22d1_hd U1107 ( .A(n1573), .B(sum[20]), .C(n1943), .D(sum[21]), .Y(n1843)
         );
  oa22d1_hd U1108 ( .A(n1839), .B(n1850), .C(n1838), .D(n1945), .Y(n1840) );
  ao21d1_hd U1109 ( .A(n1841), .B(n1850), .C(n1840), .Y(n1842) );
  oa211d1_hd U1110 ( .A(n1844), .B(n1956), .C(n1843), .D(n1842), .Y(n400) );
  ao22d1_hd U1111 ( .A(n1573), .B(sum[19]), .C(n1943), .D(sum[20]), .Y(n1849)
         );
  scg20d1_hd U1112 ( .A(n2258), .B(n1845), .C(n1932), .Y(n1853) );
  oa21d1_hd U1113 ( .A(z_m[15]), .B(n1931), .C(n1853), .Y(n1847) );
  oa21d1_hd U1114 ( .A(z_m[16]), .B(n1852), .C(n1956), .Y(n1846) );
  ao22d1_hd U1115 ( .A(z_m[16]), .B(n1847), .C(z_m[15]), .D(n1846), .Y(n1848)
         );
  oa211d1_hd U1116 ( .A(n1850), .B(n1945), .C(n1849), .D(n1848), .Y(n401) );
  ao22d1_hd U1117 ( .A(n1573), .B(sum[18]), .C(n1943), .D(sum[19]), .Y(n1856)
         );
  ao22d1_hd U1118 ( .A(z_m[15]), .B(n1853), .C(n1852), .D(n1851), .Y(n1854) );
  ao21d1_hd U1119 ( .A(z_m[16]), .B(n1938), .C(n1854), .Y(n1855) );
  oa211d1_hd U1120 ( .A(n1862), .B(n1956), .C(n1856), .D(n1855), .Y(n402) );
  nr2d1_hd U1121 ( .A(n1931), .B(n1857), .Y(n1865) );
  ao21d1_hd U1122 ( .A(n1865), .B(n1862), .C(n1949), .Y(n1861) );
  ao22d1_hd U1123 ( .A(n1573), .B(sum[17]), .C(n1943), .D(sum[18]), .Y(n1860)
         );
  ao21d1_hd U1124 ( .A(n1971), .B(n1857), .C(n1932), .Y(n1863) );
  oa21d1_hd U1125 ( .A(z_m[13]), .B(n1931), .C(n1863), .Y(n1858) );
  ao22d1_hd U1126 ( .A(z_m[14]), .B(n1858), .C(z_m[15]), .D(n1938), .Y(n1859)
         );
  oa211d1_hd U1127 ( .A(n1861), .B(n1874), .C(n1860), .D(n1859), .Y(n403) );
  ao22d1_hd U1128 ( .A(n1573), .B(sum[16]), .C(n1943), .D(sum[17]), .Y(n1867)
         );
  oa22d1_hd U1129 ( .A(n1863), .B(n1874), .C(n1862), .D(n1945), .Y(n1864) );
  ao21d1_hd U1130 ( .A(n1865), .B(n1874), .C(n1864), .Y(n1866) );
  oa211d1_hd U1131 ( .A(n1868), .B(n1956), .C(n1867), .D(n1866), .Y(n404) );
  ao22d1_hd U1132 ( .A(n1573), .B(sum[15]), .C(n1943), .D(sum[16]), .Y(n1873)
         );
  scg20d1_hd U1133 ( .A(n2258), .B(n1869), .C(n1932), .Y(n1877) );
  oa21d1_hd U1134 ( .A(z_m[11]), .B(n1931), .C(n1877), .Y(n1871) );
  oa21d1_hd U1135 ( .A(z_m[12]), .B(n1876), .C(n1956), .Y(n1870) );
  ao22d1_hd U1136 ( .A(z_m[12]), .B(n1871), .C(z_m[11]), .D(n1870), .Y(n1872)
         );
  oa211d1_hd U1137 ( .A(n1874), .B(n1945), .C(n1873), .D(n1872), .Y(n405) );
  ao22d1_hd U1138 ( .A(n1573), .B(sum[14]), .C(n1943), .D(sum[15]), .Y(n1880)
         );
  ao22d1_hd U1139 ( .A(z_m[11]), .B(n1877), .C(n1876), .D(n1875), .Y(n1878) );
  ao21d1_hd U1140 ( .A(z_m[12]), .B(n1938), .C(n1878), .Y(n1879) );
  oa211d1_hd U1141 ( .A(n1886), .B(n1956), .C(n1880), .D(n1879), .Y(n406) );
  nr2d1_hd U1142 ( .A(n1931), .B(n1881), .Y(n1889) );
  ao21d1_hd U1143 ( .A(n1889), .B(n1886), .C(n1949), .Y(n1885) );
  ao22d1_hd U1144 ( .A(n1573), .B(sum[13]), .C(n1943), .D(sum[14]), .Y(n1884)
         );
  ao21d1_hd U1145 ( .A(n1971), .B(n1881), .C(n1932), .Y(n1887) );
  oa21d1_hd U1146 ( .A(z_m[9]), .B(n1931), .C(n1887), .Y(n1882) );
  ao22d1_hd U1147 ( .A(z_m[10]), .B(n1882), .C(z_m[11]), .D(n1938), .Y(n1883)
         );
  oa211d1_hd U1148 ( .A(n1885), .B(n1898), .C(n1884), .D(n1883), .Y(n407) );
  ao22d1_hd U1149 ( .A(n1573), .B(sum[12]), .C(n1943), .D(sum[13]), .Y(n1891)
         );
  oa22d1_hd U1150 ( .A(n1887), .B(n1898), .C(n1886), .D(n1945), .Y(n1888) );
  ao21d1_hd U1151 ( .A(n1889), .B(n1898), .C(n1888), .Y(n1890) );
  oa211d1_hd U1152 ( .A(n1892), .B(n1956), .C(n1891), .D(n1890), .Y(n408) );
  ao22d1_hd U1153 ( .A(n1573), .B(sum[11]), .C(n1943), .D(sum[12]), .Y(n1897)
         );
  scg20d1_hd U1154 ( .A(n2258), .B(n1893), .C(n1932), .Y(n1901) );
  oa21d1_hd U1155 ( .A(z_m[7]), .B(n1931), .C(n1901), .Y(n1895) );
  oa21d1_hd U1156 ( .A(z_m[8]), .B(n1900), .C(n1956), .Y(n1894) );
  ao22d1_hd U1157 ( .A(z_m[8]), .B(n1895), .C(z_m[7]), .D(n1894), .Y(n1896) );
  oa211d1_hd U1158 ( .A(n1898), .B(n1945), .C(n1897), .D(n1896), .Y(n409) );
  ao22d1_hd U1159 ( .A(n1573), .B(sum[10]), .C(n1943), .D(sum[11]), .Y(n1904)
         );
  ao22d1_hd U1160 ( .A(z_m[7]), .B(n1901), .C(n1900), .D(n1899), .Y(n1902) );
  ao21d1_hd U1161 ( .A(z_m[8]), .B(n1938), .C(n1902), .Y(n1903) );
  oa211d1_hd U1162 ( .A(n1910), .B(n1956), .C(n1904), .D(n1903), .Y(n410) );
  nr2d1_hd U1163 ( .A(n1931), .B(n1905), .Y(n1913) );
  ao21d1_hd U1164 ( .A(n1913), .B(n1910), .C(n1949), .Y(n1909) );
  ao22d1_hd U1165 ( .A(n1573), .B(sum[9]), .C(n1943), .D(sum[10]), .Y(n1908)
         );
  ao21d1_hd U1166 ( .A(n1971), .B(n1905), .C(n1932), .Y(n1911) );
  oa21d1_hd U1167 ( .A(z_m[5]), .B(n1931), .C(n1911), .Y(n1906) );
  ao22d1_hd U1168 ( .A(z_m[6]), .B(n1906), .C(z_m[7]), .D(n1938), .Y(n1907) );
  oa211d1_hd U1169 ( .A(n1909), .B(n1923), .C(n1908), .D(n1907), .Y(n411) );
  ao22d1_hd U1170 ( .A(n1573), .B(sum[8]), .C(n1943), .D(sum[9]), .Y(n1915) );
  oa22d1_hd U1171 ( .A(n1911), .B(n1923), .C(n1910), .D(n1945), .Y(n1912) );
  ao21d1_hd U1172 ( .A(n1913), .B(n1923), .C(n1912), .Y(n1914) );
  oa211d1_hd U1173 ( .A(n1916), .B(n1956), .C(n1915), .D(n1914), .Y(n412) );
  ao22d1_hd U1174 ( .A(n1573), .B(sum[7]), .C(n1943), .D(sum[8]), .Y(n1922) );
  ao21d1_hd U1175 ( .A(n1971), .B(n1917), .C(n1932), .Y(n1926) );
  oa21d1_hd U1176 ( .A(z_m[3]), .B(n1931), .C(n1926), .Y(n1920) );
  oa21d1_hd U1177 ( .A(z_m[4]), .B(n1925), .C(n1956), .Y(n1919) );
  ao22d1_hd U1178 ( .A(z_m[4]), .B(n1920), .C(z_m[3]), .D(n1919), .Y(n1921) );
  oa211d1_hd U1179 ( .A(n1923), .B(n1945), .C(n1922), .D(n1921), .Y(n413) );
  ao22d1_hd U1180 ( .A(n1573), .B(sum[6]), .C(n1943), .D(sum[7]), .Y(n1929) );
  ao22d1_hd U1181 ( .A(z_m[3]), .B(n1926), .C(n1925), .D(n1924), .Y(n1927) );
  ao21d1_hd U1182 ( .A(z_m[4]), .B(n1938), .C(n1927), .Y(n1928) );
  scg15d1_hd U1183 ( .A(z_m[2]), .B(n1949), .C(n1929), .D(n1928), .Y(n414) );
  nr3d1_hd U1184 ( .A(z_m[2]), .B(n1931), .C(n1953), .Y(n1930) );
  nr2d1_hd U1185 ( .A(n1930), .B(n1949), .Y(n1936) );
  ao22d1_hd U1186 ( .A(n1573), .B(sum[5]), .C(n1943), .D(sum[6]), .Y(n1935) );
  nr2d1_hd U1187 ( .A(z_m[0]), .B(n1931), .Y(n1948) );
  nr2d1_hd U1188 ( .A(n1932), .B(n1948), .Y(n1942) );
  ao22d1_hd U1189 ( .A(z_m[2]), .B(n1933), .C(z_m[3]), .D(n1938), .Y(n1934) );
  oa211d1_hd U1190 ( .A(n1936), .B(n1946), .C(n1935), .D(n1934), .Y(n415) );
  ao22d1_hd U1191 ( .A(n1573), .B(sum[4]), .C(n1943), .D(sum[5]), .Y(n1941) );
  ao22d1_hd U1192 ( .A(z_m[0]), .B(n1939), .C(z_m[2]), .D(n1938), .Y(n1940) );
  oa211d1_hd U1193 ( .A(n1942), .B(n1946), .C(n1941), .D(n1940), .Y(n416) );
  ao22d1_hd U1194 ( .A(n1573), .B(sum[3]), .C(n1943), .D(sum[4]), .Y(n1951) );
  nr2d1_hd U1195 ( .A(n1946), .B(n1945), .Y(n1947) );
  ao211d1_hd U1196 ( .A(n1949), .B(guard), .C(n1948), .D(n1947), .Y(n1950) );
  oa211d1_hd U1197 ( .A(n1953), .B(n1952), .C(n1951), .D(n1950), .Y(n417) );
  ao21d1_hd U1198 ( .A(n1955), .B(n1965), .C(n1954), .Y(n1961) );
  oa21d1_hd U1199 ( .A(n1958), .B(n1957), .C(n1956), .Y(n1959) );
  ao22d1_hd U1200 ( .A(z_m[22]), .B(n1959), .C(n1972), .D(sum[26]), .Y(n1960)
         );
  oa211d1_hd U1201 ( .A(n1961), .B(n1964), .C(n1960), .D(n1969), .Y(n418) );
  nr4d1_hd U1202 ( .A(n1965), .B(n1964), .C(n1963), .D(n1962), .Y(n1966) );
  nd4d1_hd U1203 ( .A(z_m[21]), .B(z_m[20]), .C(n1967), .D(n1966), .Y(n1968)
         );
  nd4d1_hd U1204 ( .A(n1970), .B(n2269), .C(n1969), .D(n1968), .Y(n1984) );
  nr3d1_hd U1205 ( .A(n1972), .B(state[1]), .C(n1971), .Y(n1973) );
  ao22d1_hd U1206 ( .A(a_e[8]), .B(n1570), .C(n1990), .D(C91_DATA2_8), .Y(
        n1974) );
  oa21d1_hd U1207 ( .A(n1975), .B(n1984), .C(n1974), .Y(n419) );
  ao22d1_hd U1208 ( .A(z_e[7]), .B(n1986), .C(n1990), .D(C91_DATA2_7), .Y(
        n1976) );
  oa21d1_hd U1209 ( .A(n2101), .B(n2269), .C(n1976), .Y(n420) );
  ao22d1_hd U1210 ( .A(z_e[6]), .B(n1986), .C(n1990), .D(C91_DATA2_6), .Y(
        n1977) );
  oa21d1_hd U1211 ( .A(n2097), .B(n2269), .C(n1977), .Y(n421) );
  ao22d1_hd U1212 ( .A(z_e[5]), .B(n1986), .C(n1990), .D(C91_DATA2_5), .Y(
        n1978) );
  oa21d1_hd U1213 ( .A(n2116), .B(n2269), .C(n1978), .Y(n422) );
  ao22d1_hd U1214 ( .A(z_e[4]), .B(n1986), .C(n1990), .D(C91_DATA2_4), .Y(
        n1979) );
  oa21d1_hd U1215 ( .A(n2121), .B(n2269), .C(n1979), .Y(n423) );
  ao22d1_hd U1216 ( .A(z_e[3]), .B(n1986), .C(n1990), .D(C91_DATA2_3), .Y(
        n1980) );
  oa21d1_hd U1217 ( .A(n2128), .B(n2269), .C(n1980), .Y(n424) );
  ao22d1_hd U1218 ( .A(z_e[2]), .B(n1986), .C(n1990), .D(C91_DATA2_2), .Y(
        n1981) );
  oa21d1_hd U1219 ( .A(n2137), .B(n2269), .C(n1981), .Y(n425) );
  ao22d1_hd U1220 ( .A(z_e[1]), .B(n1986), .C(n1990), .D(C91_DATA2_1), .Y(
        n1982) );
  oa21d1_hd U1221 ( .A(n2145), .B(n2269), .C(n1982), .Y(n426) );
  ao22d1_hd U1222 ( .A(a_e[0]), .B(n1570), .C(n1990), .D(n1985), .Y(n1983) );
  oa21d1_hd U1223 ( .A(n1985), .B(n1984), .C(n1983), .Y(n427) );
  ao22d1_hd U1224 ( .A(a_e[9]), .B(n1570), .C(z_e[9]), .D(n1986), .Y(n1993) );
  ao22d1_hd U1225 ( .A(z_e[9]), .B(n2266), .C(n1988), .D(n1987), .Y(n1991) );
  oa211d1_hd U1226 ( .A(DP_OP_154J4_137_6175_n2), .B(n1991), .C(n1990), .D(
        n1989), .Y(n1992) );
  ao22d1_hd U1227 ( .A(b_m[25]), .B(n2036), .C(n1578), .D(b[21]), .Y(n1994) );
  oa21d1_hd U1228 ( .A(n1995), .B(n1576), .C(n1994), .Y(n429) );
  ao22d1_hd U1229 ( .A(b_m[24]), .B(n2036), .C(n1579), .D(b[20]), .Y(n1996) );
  oa21d1_hd U1230 ( .A(n1997), .B(n1576), .C(n1996), .Y(n430) );
  ao22d1_hd U1231 ( .A(b_m[23]), .B(n2036), .C(n1580), .D(b[19]), .Y(n1998) );
  oa21d1_hd U1232 ( .A(n1999), .B(n1576), .C(n1998), .Y(n431) );
  ao22d1_hd U1233 ( .A(b_m[22]), .B(n2036), .C(n1579), .D(b[18]), .Y(n2000) );
  oa21d1_hd U1234 ( .A(n2001), .B(n1576), .C(n2000), .Y(n432) );
  ao22d1_hd U1235 ( .A(b_m[21]), .B(n2036), .C(n1579), .D(b[17]), .Y(n2002) );
  oa21d1_hd U1236 ( .A(n2003), .B(n1576), .C(n2002), .Y(n433) );
  ao22d1_hd U1237 ( .A(b_m[20]), .B(n2036), .C(n1579), .D(b[16]), .Y(n2004) );
  oa21d1_hd U1238 ( .A(n2005), .B(n1576), .C(n2004), .Y(n434) );
  ao22d1_hd U1239 ( .A(b_m[19]), .B(n2036), .C(n1579), .D(b[15]), .Y(n2006) );
  oa21d1_hd U1240 ( .A(n2007), .B(n1576), .C(n2006), .Y(n435) );
  ao22d1_hd U1241 ( .A(b_m[18]), .B(n2036), .C(n1579), .D(b[14]), .Y(n2008) );
  oa21d1_hd U1242 ( .A(n2009), .B(n1576), .C(n2008), .Y(n436) );
  ao22d1_hd U1243 ( .A(b_m[17]), .B(n2036), .C(n1579), .D(b[13]), .Y(n2010) );
  oa21d1_hd U1244 ( .A(n2011), .B(n1576), .C(n2010), .Y(n437) );
  ao22d1_hd U1245 ( .A(b_m[16]), .B(n2036), .C(n1579), .D(b[12]), .Y(n2012) );
  oa21d1_hd U1246 ( .A(n2013), .B(n1576), .C(n2012), .Y(n438) );
  ao22d1_hd U1247 ( .A(b_m[15]), .B(n2036), .C(n1579), .D(b[11]), .Y(n2014) );
  oa21d1_hd U1248 ( .A(n2015), .B(n1576), .C(n2014), .Y(n439) );
  ao22d1_hd U1249 ( .A(b_m[14]), .B(n2036), .C(n1579), .D(b[10]), .Y(n2016) );
  oa21d1_hd U1250 ( .A(n2017), .B(n1576), .C(n2016), .Y(n440) );
  ao22d1_hd U1251 ( .A(b_m[13]), .B(n2036), .C(n1579), .D(b[9]), .Y(n2018) );
  oa21d1_hd U1252 ( .A(n2019), .B(n1576), .C(n2018), .Y(n441) );
  ao22d1_hd U1253 ( .A(b_m[12]), .B(n2036), .C(n1579), .D(b[8]), .Y(n2020) );
  oa21d1_hd U1254 ( .A(n2021), .B(n1576), .C(n2020), .Y(n442) );
  ao22d1_hd U1255 ( .A(b_m[11]), .B(n2036), .C(n1579), .D(b[7]), .Y(n2022) );
  oa21d1_hd U1256 ( .A(n2023), .B(n1576), .C(n2022), .Y(n443) );
  ao22d1_hd U1257 ( .A(b_m[10]), .B(n2036), .C(n1579), .D(b[6]), .Y(n2024) );
  oa21d1_hd U1258 ( .A(n2025), .B(n1576), .C(n2024), .Y(n444) );
  ao22d1_hd U1259 ( .A(b_m[9]), .B(n2036), .C(n1579), .D(b[5]), .Y(n2026) );
  oa21d1_hd U1260 ( .A(n2027), .B(n1576), .C(n2026), .Y(n445) );
  ao22d1_hd U1261 ( .A(b_m[8]), .B(n2036), .C(n1579), .D(b[4]), .Y(n2028) );
  oa21d1_hd U1262 ( .A(n2029), .B(n1576), .C(n2028), .Y(n446) );
  ao22d1_hd U1263 ( .A(b_m[7]), .B(n2036), .C(n1579), .D(b[3]), .Y(n2030) );
  oa21d1_hd U1264 ( .A(n2031), .B(n1576), .C(n2030), .Y(n447) );
  ao22d1_hd U1265 ( .A(b_m[6]), .B(n2036), .C(n1579), .D(b[2]), .Y(n2032) );
  oa21d1_hd U1266 ( .A(n2033), .B(n1576), .C(n2032), .Y(n448) );
  ao22d1_hd U1267 ( .A(b_m[5]), .B(n2036), .C(n1579), .D(b[1]), .Y(n2034) );
  oa21d1_hd U1268 ( .A(n2035), .B(n1576), .C(n2034), .Y(n449) );
  ao22d1_hd U1269 ( .A(b_m[4]), .B(n2036), .C(n1579), .D(b[0]), .Y(n2037) );
  oa21d1_hd U1270 ( .A(n2038), .B(n1576), .C(n2037), .Y(n450) );
  oa22d1_hd U1271 ( .A(n2039), .B(n1576), .C(n2038), .D(n2249), .Y(n451) );
  oa22d1_hd U1272 ( .A(n2040), .B(n1576), .C(n2039), .D(n2249), .Y(n452) );
  oa22d1_hd U1273 ( .A(n1580), .B(n2041), .C(n2040), .D(n2249), .Y(n453) );
  ao22d1_hd U1274 ( .A(a_m[25]), .B(n2084), .C(n1579), .D(a[21]), .Y(n2042) );
  oa21d1_hd U1275 ( .A(n2043), .B(n1574), .C(n2042), .Y(n454) );
  ao22d1_hd U1276 ( .A(a_m[24]), .B(n2084), .C(n1579), .D(a[20]), .Y(n2044) );
  oa21d1_hd U1277 ( .A(n2045), .B(n1574), .C(n2044), .Y(n455) );
  ao22d1_hd U1278 ( .A(a_m[23]), .B(n2084), .C(n1579), .D(a[19]), .Y(n2046) );
  oa21d1_hd U1279 ( .A(n2047), .B(n1574), .C(n2046), .Y(n456) );
  ao22d1_hd U1280 ( .A(a_m[22]), .B(n2084), .C(n1579), .D(a[18]), .Y(n2048) );
  oa21d1_hd U1281 ( .A(n2049), .B(n1574), .C(n2048), .Y(n457) );
  ao22d1_hd U1282 ( .A(a_m[21]), .B(n2084), .C(n1579), .D(a[17]), .Y(n2050) );
  oa21d1_hd U1283 ( .A(n2051), .B(n1574), .C(n2050), .Y(n458) );
  ao22d1_hd U1284 ( .A(a_m[20]), .B(n2084), .C(n1580), .D(a[16]), .Y(n2052) );
  oa21d1_hd U1285 ( .A(n2053), .B(n1574), .C(n2052), .Y(n459) );
  ao22d1_hd U1286 ( .A(a_m[19]), .B(n2084), .C(n1579), .D(a[15]), .Y(n2054) );
  oa21d1_hd U1287 ( .A(n2055), .B(n1574), .C(n2054), .Y(n460) );
  ao22d1_hd U1288 ( .A(a_m[18]), .B(n2084), .C(n1579), .D(a[14]), .Y(n2056) );
  oa21d1_hd U1289 ( .A(n2057), .B(n1574), .C(n2056), .Y(n461) );
  ao22d1_hd U1290 ( .A(a_m[17]), .B(n2084), .C(n1580), .D(a[13]), .Y(n2058) );
  oa21d1_hd U1291 ( .A(n2059), .B(n1574), .C(n2058), .Y(n462) );
  ao22d1_hd U1292 ( .A(a_m[16]), .B(n2084), .C(n1579), .D(a[12]), .Y(n2060) );
  oa21d1_hd U1293 ( .A(n2061), .B(n1574), .C(n2060), .Y(n463) );
  ao22d1_hd U1294 ( .A(a_m[15]), .B(n2084), .C(n1580), .D(a[11]), .Y(n2062) );
  oa21d1_hd U1295 ( .A(n2063), .B(n1574), .C(n2062), .Y(n464) );
  ao22d1_hd U1296 ( .A(a_m[14]), .B(n2084), .C(n1578), .D(a[10]), .Y(n2064) );
  oa21d1_hd U1297 ( .A(n2065), .B(n1574), .C(n2064), .Y(n465) );
  ao22d1_hd U1298 ( .A(a_m[13]), .B(n2084), .C(n1578), .D(a[9]), .Y(n2066) );
  oa21d1_hd U1299 ( .A(n2067), .B(n1574), .C(n2066), .Y(n466) );
  ao22d1_hd U1300 ( .A(a_m[12]), .B(n2084), .C(n1578), .D(a[8]), .Y(n2068) );
  oa21d1_hd U1301 ( .A(n2069), .B(n1574), .C(n2068), .Y(n467) );
  ao22d1_hd U1302 ( .A(a_m[11]), .B(n2084), .C(n1578), .D(a[7]), .Y(n2070) );
  oa21d1_hd U1303 ( .A(n2071), .B(n1574), .C(n2070), .Y(n468) );
  ao22d1_hd U1304 ( .A(a_m[10]), .B(n2084), .C(n1578), .D(a[6]), .Y(n2072) );
  oa21d1_hd U1305 ( .A(n2073), .B(n1574), .C(n2072), .Y(n469) );
  ao22d1_hd U1306 ( .A(a_m[9]), .B(n2084), .C(n1578), .D(a[5]), .Y(n2074) );
  oa21d1_hd U1307 ( .A(n2075), .B(n1574), .C(n2074), .Y(n470) );
  ao22d1_hd U1308 ( .A(a_m[8]), .B(n2084), .C(n1578), .D(a[4]), .Y(n2076) );
  oa21d1_hd U1309 ( .A(n2077), .B(n1574), .C(n2076), .Y(n471) );
  ao22d1_hd U1310 ( .A(a_m[7]), .B(n2084), .C(n1578), .D(a[3]), .Y(n2078) );
  oa21d1_hd U1311 ( .A(n2079), .B(n1574), .C(n2078), .Y(n472) );
  ao22d1_hd U1312 ( .A(a_m[6]), .B(n2084), .C(n1579), .D(a[2]), .Y(n2080) );
  oa21d1_hd U1313 ( .A(n2081), .B(n1574), .C(n2080), .Y(n473) );
  ao22d1_hd U1314 ( .A(a_m[5]), .B(n2084), .C(n1578), .D(a[1]), .Y(n2082) );
  oa21d1_hd U1315 ( .A(n2083), .B(n1574), .C(n2082), .Y(n474) );
  ao22d1_hd U1316 ( .A(a_m[4]), .B(n2084), .C(n1578), .D(a[0]), .Y(n2085) );
  oa21d1_hd U1317 ( .A(n2086), .B(n1574), .C(n2085), .Y(n475) );
  oa22d1_hd U1318 ( .A(n2087), .B(n1574), .C(n2086), .D(n2091), .Y(n476) );
  oa22d1_hd U1319 ( .A(n2088), .B(n1574), .C(n2087), .D(n2091), .Y(n477) );
  oa22d1_hd U1320 ( .A(n1580), .B(n2089), .C(n2088), .D(n2091), .Y(n478) );
  ao22d1_hd U1321 ( .A(a_m[25]), .B(n1575), .C(n1578), .D(a[22]), .Y(n2090) );
  oa21d1_hd U1322 ( .A(n2092), .B(n2091), .C(n2090), .Y(n479) );
  nr2d1_hd U1323 ( .A(n2145), .B(n2144), .Y(n2133) );
  nr2d1_hd U1324 ( .A(n2128), .B(n2127), .Y(n2118) );
  ao21d1_hd U1325 ( .A(n2186), .B(n2096), .C(n2151), .Y(n2117) );
  oa21d1_hd U1326 ( .A(n2097), .B(n2116), .C(n2186), .Y(n2095) );
  ao21d1_hd U1327 ( .A(n2136), .B(n2101), .C(n2103), .Y(n2153) );
  ivd1_hd U1328 ( .A(a[25]), .Y(n2135) );
  nr2d1_hd U1329 ( .A(n2147), .B(n2135), .Y(n2134) );
  ivd1_hd U1330 ( .A(a[27]), .Y(n2120) );
  nr2d1_hd U1331 ( .A(n2130), .B(n2120), .Y(n2119) );
  ivd1_hd U1332 ( .A(a[29]), .Y(n2106) );
  nr2d1_hd U1333 ( .A(n2113), .B(n2106), .Y(n2100) );
  nr2d1_hd U1334 ( .A(n2100), .B(n2268), .Y(n2108) );
  nr2d1_hd U1335 ( .A(n2154), .B(n2096), .Y(n2112) );
  nr2d1_hd U1336 ( .A(n2097), .B(n2111), .Y(n2102) );
  nd3d1_hd U1337 ( .A(a_e[7]), .B(n2102), .C(n2099), .Y(n2098) );
  oa211d1_hd U1338 ( .A(n2153), .B(n2099), .C(n2155), .D(n2098), .Y(n480) );
  ao22d1_hd U1339 ( .A(a_e[7]), .B(n2103), .C(n2102), .D(n2101), .Y(n2104) );
  oa211d1_hd U1340 ( .A(n2268), .B(n2105), .C(n2104), .D(n2155), .Y(n481) );
  oa21d1_hd U1341 ( .A(a_e[5]), .B(n2154), .C(n2117), .Y(n2109) );
  ao22d1_hd U1342 ( .A(a_e[6]), .B(n2109), .C(n2108), .D(n2107), .Y(n2110) );
  oa211d1_hd U1343 ( .A(a_e[6]), .B(n2111), .C(n2110), .D(n2140), .Y(n482) );
  ao21d1_hd U1344 ( .A(n2112), .B(n2116), .C(n2156), .Y(n2115) );
  oa211d1_hd U1345 ( .A(n2119), .B(a[28]), .C(n1580), .D(n2113), .Y(n2114) );
  oa211d1_hd U1346 ( .A(n2117), .B(n2116), .C(n2115), .D(n2114), .Y(n483) );
  ao211d1_hd U1347 ( .A(n2130), .B(n2120), .C(n2119), .D(n2268), .Y(n2123) );
  ao21d1_hd U1348 ( .A(n2186), .B(n2127), .C(n2151), .Y(n2129) );
  ao21d1_hd U1349 ( .A(n2129), .B(n2126), .C(n2121), .Y(n2122) );
  nr2d1_hd U1350 ( .A(n2123), .B(n2122), .Y(n2124) );
  oa211d1_hd U1351 ( .A(a_e[4]), .B(n2125), .C(n2124), .D(n2140), .Y(n484) );
  oa22d1_hd U1352 ( .A(n2129), .B(n2128), .C(n2127), .D(n2126), .Y(n2132) );
  oa211d1_hd U1353 ( .A(n2134), .B(a[26]), .C(n1580), .D(n2130), .Y(n2131) );
  scg13d1_hd U1354 ( .A(n2132), .B(n2156), .C(n2131), .Y(n485) );
  ao211d1_hd U1355 ( .A(n2147), .B(n2135), .C(n2134), .D(n2268), .Y(n2139) );
  nr2d1_hd U1356 ( .A(a_e[0]), .B(n2154), .Y(n2150) );
  nr2d1_hd U1357 ( .A(n2151), .B(n2150), .Y(n2146) );
  ao21d1_hd U1358 ( .A(n2146), .B(n2143), .C(n2137), .Y(n2138) );
  nr2d1_hd U1359 ( .A(n2139), .B(n2138), .Y(n2141) );
  oa211d1_hd U1360 ( .A(a_e[2]), .B(n2142), .C(n2141), .D(n2140), .Y(n486) );
  oa22d1_hd U1361 ( .A(n2146), .B(n2145), .C(n2144), .D(n2143), .Y(n2149) );
  oa211d1_hd U1362 ( .A(a[23]), .B(a[24]), .C(n1580), .D(n2147), .Y(n2148) );
  scg13d1_hd U1363 ( .A(n2149), .B(n2156), .C(n2148), .Y(n487) );
  ao21d1_hd U1364 ( .A(n2151), .B(a_e[0]), .C(n2150), .Y(n2152) );
  oa21d1_hd U1365 ( .A(a[23]), .B(n2268), .C(n2152), .Y(n488) );
  oa21d1_hd U1366 ( .A(a_e[8]), .B(n2154), .C(n2153), .Y(n2157) );
  scg17d1_hd U1367 ( .A(a_e[9]), .B(n2157), .C(n2156), .D(n2155), .Y(n489) );
  nr2d1_hd U1368 ( .A(n2212), .B(n2211), .Y(n2201) );
  nr2d1_hd U1369 ( .A(n2161), .B(n2195), .Y(n2191) );
  ao21d1_hd U1370 ( .A(n2162), .B(n2186), .C(n2218), .Y(n2185) );
  oa21d1_hd U1371 ( .A(n2164), .B(n2184), .C(n2186), .Y(n2163) );
  ao21d1_hd U1372 ( .A(n2202), .B(n2168), .C(n2170), .Y(n2251) );
  ivd1_hd U1373 ( .A(b[25]), .Y(n2204) );
  nr2d1_hd U1374 ( .A(n2214), .B(n2204), .Y(n2203) );
  ivd1_hd U1375 ( .A(b[27]), .Y(n2188) );
  nr2d1_hd U1376 ( .A(n2198), .B(n2188), .Y(n2187) );
  ivd1_hd U1377 ( .A(b[29]), .Y(n2174) );
  nr2d1_hd U1378 ( .A(n2181), .B(n2174), .Y(n2167) );
  nr2d1_hd U1379 ( .A(n2167), .B(n2268), .Y(n2177) );
  nr2bd1_hd U1380 ( .AN(n2191), .B(n2194), .Y(n2180) );
  nr2d1_hd U1381 ( .A(n2164), .B(n2179), .Y(n2169) );
  nd3d1_hd U1382 ( .A(b_e[7]), .B(n2169), .C(n2166), .Y(n2165) );
  oa211d1_hd U1383 ( .A(n2251), .B(n2166), .C(n2253), .D(n2165), .Y(n490) );
  ao22d1_hd U1384 ( .A(b_e[7]), .B(n2170), .C(n2169), .D(n2168), .Y(n2171) );
  oa211d1_hd U1385 ( .A(n2173), .B(n2172), .C(n2171), .D(n2253), .Y(n491) );
  oa21d1_hd U1386 ( .A(b_e[5]), .B(n2252), .C(n2185), .Y(n2175) );
  ao22d1_hd U1387 ( .A(n2177), .B(n2176), .C(b_e[6]), .D(n2175), .Y(n2178) );
  oa211d1_hd U1388 ( .A(b_e[6]), .B(n2179), .C(n2178), .D(n2207), .Y(n492) );
  ao21d1_hd U1389 ( .A(n2180), .B(n2184), .C(n2254), .Y(n2183) );
  oa211d1_hd U1390 ( .A(n2187), .B(b[28]), .C(n1580), .D(n2181), .Y(n2182) );
  oa211d1_hd U1391 ( .A(n2185), .B(n2184), .C(n2183), .D(n2182), .Y(n493) );
  scg6d1_hd U1392 ( .A(n2195), .B(n2186), .C(n2218), .Y(n2197) );
  ao211d1_hd U1393 ( .A(n2198), .B(n2188), .C(n2187), .D(n2268), .Y(n2189) );
  ao211d1_hd U1394 ( .A(b_e[4]), .B(n2197), .C(n2254), .D(n2189), .Y(n2193) );
  nd3d1_hd U1395 ( .A(n2202), .B(n2191), .C(n2190), .Y(n2192) );
  oa211d1_hd U1396 ( .A(b_e[3]), .B(n2194), .C(n2193), .D(n2192), .Y(n494) );
  nr3d1_hd U1397 ( .A(b_e[3]), .B(n2252), .C(n2195), .Y(n2196) );
  ao211d1_hd U1398 ( .A(b_e[3]), .B(n2197), .C(n2254), .D(n2196), .Y(n2200) );
  oa211d1_hd U1399 ( .A(n2203), .B(b[26]), .C(n1580), .D(n2198), .Y(n2199) );
  nr2d1_hd U1400 ( .A(b_e[0]), .B(n2252), .Y(n2217) );
  nr2d1_hd U1401 ( .A(n2218), .B(n2217), .Y(n2213) );
  ao211d1_hd U1402 ( .A(n2214), .B(n2204), .C(n2203), .D(n2268), .Y(n2205) );
  ao21d1_hd U1403 ( .A(n2206), .B(b_e[2]), .C(n2205), .Y(n2208) );
  oa211d1_hd U1404 ( .A(b_e[2]), .B(n2209), .C(n2208), .D(n2207), .Y(n496) );
  oa22d1_hd U1405 ( .A(n2213), .B(n2212), .C(n2211), .D(n2210), .Y(n2216) );
  oa211d1_hd U1406 ( .A(b[23]), .B(b[24]), .C(n1580), .D(n2214), .Y(n2215) );
  scg13d1_hd U1407 ( .A(n2216), .B(n2254), .C(n2215), .Y(n497) );
  ao21d1_hd U1408 ( .A(n2218), .B(b_e[0]), .C(n2217), .Y(n2219) );
  oa21d1_hd U1409 ( .A(b[23]), .B(n2268), .C(n2219), .Y(n498) );
  scg21d1_hd U1410 ( .A(n2220), .B(o_AB_ACK), .C(i_RST), .D(n1571), .Y(n499)
         );
  oa211d1_hd U1411 ( .A(state[3]), .B(n2225), .C(n2224), .D(n2223), .Y(n2239)
         );
  nd3d1_hd U1412 ( .A(n1581), .B(o_Z_STB), .C(i_Z_ACK), .Y(n2263) );
  nd4d1_hd U1413 ( .A(N41), .B(n2258), .C(n2263), .D(n2269), .Y(n2226) );
  nr3d1_hd U1414 ( .A(n27), .B(n2239), .C(n2226), .Y(n2231) );
  ao22d1_hd U1415 ( .A(n2229), .B(n2228), .C(n2266), .D(n2227), .Y(n2230) );
  oa211d1_hd U1416 ( .A(n2233), .B(n2232), .C(n2231), .D(n2230), .Y(n2259) );
  ivd1_hd U1417 ( .A(n2259), .Y(n2236) );
  nr2d1_hd U1418 ( .A(n2234), .B(n2244), .Y(n2235) );
  ao22d1_hd U1419 ( .A(state[2]), .B(n2236), .C(N41), .D(n2235), .Y(n2237) );
  oa21d1_hd U1420 ( .A(n2238), .B(n2261), .C(n2237), .Y(n500) );
  nr2d1_hd U1421 ( .A(n2266), .B(n2239), .Y(n2241) );
  oa22d1_hd U1422 ( .A(n2241), .B(n2261), .C(n2240), .D(n2259), .Y(n501) );
  oa211d1_hd U1423 ( .A(n2244), .B(state[0]), .C(n2243), .D(n2242), .Y(n2245)
         );
  ivd1_hd U1424 ( .A(n2245), .Y(n2247) );
  oa22d1_hd U1425 ( .A(n2247), .B(n2261), .C(n2246), .D(n2259), .Y(n502) );
  ao22d1_hd U1426 ( .A(b_m[25]), .B(n2158), .C(n1578), .D(b[22]), .Y(n2248) );
  oa21d1_hd U1427 ( .A(n2250), .B(n2249), .C(n2248), .Y(n503) );
  oa21d1_hd U1428 ( .A(b_e[8]), .B(n2252), .C(n2251), .Y(n2255) );
  scg17d1_hd U1429 ( .A(b_e[9]), .B(n2255), .C(n2254), .D(n2253), .Y(n504) );
  oa22d1_hd U1430 ( .A(n2262), .B(n2261), .C(n2260), .D(n2259), .Y(n505) );
  ivd1_hd U1431 ( .A(n2263), .Y(n2264) );
  scg21d1_hd U1432 ( .A(n1581), .B(o_Z_STB), .C(i_RST), .D(n2264), .Y(n506) );
endmodule


module iir_hpf ( i_X_DATA, i_X_DATA_VALID, o_X_DATA_READY, o_Y_DATA, 
        o_Y_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN );
  input [31:0] i_X_DATA;
  output [31:0] o_Y_DATA;
  input i_X_DATA_VALID, i_Y_ACK, i_CLK, i_RSTN;
  output o_X_DATA_READY, o_Y_DATA_VALID;
  wire   r_add_AB_STB, w_add_AB_ACK, w_add_Z_STB, r_add_Z_ACK, r_mult_AB_STB,
         w_mult_AB_ACK, w_mult_Z_STB, r_mult_Z_ACK, n_1_net_, N17, r_pstate_0_,
         N553, N559, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n221, n223, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n447, n448, n450, n594, n595, n597, n598,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n694, n695, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n731, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n801, n803, n804, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n825, n826, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n215, n216, n217,
         n218, n219, n220, n222, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n445, n446, n449, n451;
  wire   [31:0] r_add_A;
  wire   [31:0] r_add_B;
  wire   [31:0] w_add_Z;
  wire   [31:0] r_mult_A;
  wire   [31:0] r_mult_B;
  wire   [31:0] w_mult_Z;
  wire   [63:0] r_x_data;
  wire   [31:0] r_y_data;

  float_adder_2 add ( .i_A(r_add_A), .i_B(r_add_B), .i_AB_STB(r_add_AB_STB), 
        .o_AB_ACK(w_add_AB_ACK), .o_Z(w_add_Z), .o_Z_STB(w_add_Z_STB), 
        .i_Z_ACK(r_add_Z_ACK), .i_CLK(i_CLK), .i_RST(N17) );
  float_multiplier mult ( .i_A(r_mult_A), .i_B(r_mult_B), .i_AB_STB(
        r_mult_AB_STB), .o_AB_ACK(w_mult_AB_ACK), .o_Z(w_mult_Z), .o_Z_STB(
        w_mult_Z_STB), .i_Z_ACK(r_mult_Z_ACK), .i_CLK(i_CLK), .i_RST(n_1_net_)
         );
  ivd1_hd I_5 ( .A(i_RSTN), .Y(n_1_net_) );
  fd3qd1_hd r_pstate_reg_1_ ( .D(n212), .CK(i_CLK), .SN(i_RSTN), .Q(n213) );
  fd3qd1_hd r_counter_reg_1_ ( .D(n211), .CK(i_CLK), .SN(i_RSTN), .Q(n221) );
  fd3qd1_hd r_counter_reg_0_ ( .D(n210), .CK(i_CLK), .SN(i_RSTN), .Q(n223) );
  ivd1_hd U456 ( .A(i_RSTN), .Y(N17) );
  fd2qd1_hd r_mult_A_reg_2_ ( .D(n78), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[2]) );
  fd2qd1_hd r_mult_A_reg_3_ ( .D(n77), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[3]) );
  fd2qd1_hd r_mult_A_reg_4_ ( .D(n76), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[4]) );
  fd2qd1_hd r_mult_A_reg_10_ ( .D(n70), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[10]) );
  fd2qd1_hd r_mult_A_reg_12_ ( .D(n68), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[12]) );
  fd2qd1_hd r_mult_A_reg_15_ ( .D(n65), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[15]) );
  fd2qd1_hd r_mult_A_reg_18_ ( .D(n62), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[18]) );
  fd2qd1_hd r_mult_A_reg_19_ ( .D(n61), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[19]) );
  fd2qd1_hd r_mult_A_reg_20_ ( .D(n60), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[20]) );
  fd2qd1_hd r_mult_A_reg_23_ ( .D(n57), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[23]) );
  fd2qd1_hd r_mult_A_reg_30_ ( .D(n50), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[30]) );
  fd2qd1_hd r_mult_A_reg_31_ ( .D(n49), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[31]) );
  fd2qd1_hd r_mult_AB_STB_reg ( .D(n145), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_AB_STB) );
  fd2qd1_hd r_mult_B_reg_31_ ( .D(n214), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[31]) );
  fd2qd1_hd r_mult_B_reg_0_ ( .D(n111), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[0]) );
  fd2qd1_hd r_mult_B_reg_1_ ( .D(n110), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[1]) );
  fd2qd1_hd r_mult_B_reg_2_ ( .D(n109), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[2]) );
  fd2qd1_hd r_mult_B_reg_3_ ( .D(n108), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[3]) );
  fd2qd1_hd r_mult_B_reg_4_ ( .D(n107), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[4]) );
  fd2qd1_hd r_mult_B_reg_5_ ( .D(n106), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[5]) );
  fd2qd1_hd r_mult_B_reg_6_ ( .D(n105), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[6]) );
  fd2qd1_hd r_mult_B_reg_7_ ( .D(n104), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[7]) );
  fd2qd1_hd r_mult_B_reg_8_ ( .D(n103), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[8]) );
  fd2qd1_hd r_mult_B_reg_9_ ( .D(n102), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[9]) );
  fd2qd1_hd r_mult_B_reg_10_ ( .D(n101), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[10]) );
  fd2qd1_hd r_mult_B_reg_11_ ( .D(n100), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[11]) );
  fd2qd1_hd r_mult_B_reg_12_ ( .D(n99), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[12]) );
  fd2qd1_hd r_mult_B_reg_13_ ( .D(n98), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[13]) );
  fd2qd1_hd r_mult_B_reg_14_ ( .D(n97), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[14]) );
  fd2qd1_hd r_mult_B_reg_15_ ( .D(n96), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[15]) );
  fd2qd1_hd r_mult_B_reg_16_ ( .D(n95), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[16]) );
  fd2qd1_hd r_mult_B_reg_17_ ( .D(n94), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[17]) );
  fd2qd1_hd r_mult_B_reg_18_ ( .D(n93), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[18]) );
  fd2qd1_hd r_mult_B_reg_19_ ( .D(n92), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[19]) );
  fd2qd1_hd r_mult_B_reg_20_ ( .D(n91), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[20]) );
  fd2qd1_hd r_mult_B_reg_21_ ( .D(n90), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[21]) );
  fd2qd1_hd r_mult_B_reg_22_ ( .D(n89), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[22]) );
  fd2qd1_hd r_mult_B_reg_23_ ( .D(n88), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[23]) );
  fd2qd1_hd r_mult_B_reg_24_ ( .D(n87), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[24]) );
  fd2qd1_hd r_mult_B_reg_25_ ( .D(n86), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[25]) );
  fd2qd1_hd r_mult_B_reg_26_ ( .D(n85), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[26]) );
  fd2qd1_hd r_mult_B_reg_27_ ( .D(n84), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[27]) );
  fd2qd1_hd r_mult_B_reg_28_ ( .D(n83), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[28]) );
  fd2qd1_hd r_mult_B_reg_29_ ( .D(n82), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[29]) );
  fd2qd1_hd r_mult_B_reg_30_ ( .D(n81), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_B[30]) );
  fd2qd1_hd r_mult_A_reg_0_ ( .D(n80), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[0]) );
  fd2qd1_hd r_mult_A_reg_1_ ( .D(n79), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[1]) );
  fd2qd1_hd r_mult_A_reg_5_ ( .D(n75), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[5]) );
  fd2qd1_hd r_mult_A_reg_6_ ( .D(n74), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[6]) );
  fd2qd1_hd r_mult_A_reg_7_ ( .D(n73), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[7]) );
  fd2qd1_hd r_mult_A_reg_8_ ( .D(n72), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[8]) );
  fd2qd1_hd r_mult_A_reg_9_ ( .D(n71), .CK(i_CLK), .RN(i_RSTN), .Q(r_mult_A[9]) );
  fd2qd1_hd r_mult_A_reg_11_ ( .D(n69), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[11]) );
  fd2qd1_hd r_mult_A_reg_13_ ( .D(n67), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[13]) );
  fd2qd1_hd r_mult_A_reg_14_ ( .D(n66), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[14]) );
  fd2qd1_hd r_mult_A_reg_16_ ( .D(n64), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[16]) );
  fd2qd1_hd r_mult_A_reg_17_ ( .D(n63), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[17]) );
  fd2qd1_hd r_mult_A_reg_21_ ( .D(n59), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[21]) );
  fd2qd1_hd r_mult_A_reg_22_ ( .D(n58), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[22]) );
  fd2qd1_hd r_mult_A_reg_24_ ( .D(n56), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[24]) );
  fd2qd1_hd r_mult_A_reg_25_ ( .D(n55), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[25]) );
  fd2qd1_hd r_mult_A_reg_26_ ( .D(n54), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[26]) );
  fd2qd1_hd r_mult_A_reg_27_ ( .D(n53), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[27]) );
  fd2qd1_hd r_mult_A_reg_28_ ( .D(n52), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[28]) );
  fd2qd1_hd r_mult_A_reg_29_ ( .D(n51), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_A[29]) );
  fd2qd1_hd r_mult_Z_ACK_reg ( .D(n144), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_mult_Z_ACK) );
  fd2qd1_hd r_add_A_reg_30_ ( .D(n413), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[30]) );
  fd2qd1_hd r_add_A_reg_29_ ( .D(n414), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[29]) );
  fd2qd1_hd r_add_A_reg_28_ ( .D(n415), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[28]) );
  fd2qd1_hd r_add_A_reg_27_ ( .D(n416), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[27]) );
  fd2qd1_hd r_add_A_reg_26_ ( .D(n417), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[26]) );
  fd2qd1_hd r_add_A_reg_25_ ( .D(n418), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[25]) );
  fd2qd1_hd r_add_A_reg_24_ ( .D(n419), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[24]) );
  fd2qd1_hd r_add_A_reg_23_ ( .D(n420), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[23]) );
  fd2qd1_hd r_add_A_reg_22_ ( .D(n421), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[22]) );
  fd2qd1_hd r_add_A_reg_21_ ( .D(n422), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[21]) );
  fd2qd1_hd r_add_A_reg_20_ ( .D(n423), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[20]) );
  fd2qd1_hd r_add_A_reg_19_ ( .D(n424), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[19]) );
  fd2qd1_hd r_add_A_reg_18_ ( .D(n425), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[18]) );
  fd2qd1_hd r_add_A_reg_17_ ( .D(n426), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[17]) );
  fd2qd1_hd r_add_A_reg_16_ ( .D(n427), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[16]) );
  fd2qd1_hd r_add_A_reg_15_ ( .D(n428), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[15]) );
  fd2qd1_hd r_add_A_reg_14_ ( .D(n429), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[14]) );
  fd2qd1_hd r_add_A_reg_13_ ( .D(n430), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[13]) );
  fd2qd1_hd r_add_A_reg_12_ ( .D(n431), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[12]) );
  fd2qd1_hd r_add_A_reg_11_ ( .D(n432), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[11]) );
  fd2qd1_hd r_add_A_reg_10_ ( .D(n433), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[10]) );
  fd2qd1_hd r_add_A_reg_9_ ( .D(n434), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[9])
         );
  fd2qd1_hd r_add_A_reg_8_ ( .D(n435), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[8])
         );
  fd2qd1_hd r_add_A_reg_7_ ( .D(n436), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[7])
         );
  fd2qd1_hd r_add_A_reg_6_ ( .D(n437), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[6])
         );
  fd2qd1_hd r_add_A_reg_5_ ( .D(n438), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[5])
         );
  fd2qd1_hd r_add_A_reg_4_ ( .D(n439), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[4])
         );
  fd2qd1_hd r_add_A_reg_3_ ( .D(n440), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[3])
         );
  fd2qd1_hd r_add_A_reg_2_ ( .D(n441), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[2])
         );
  fd2qd1_hd r_add_A_reg_1_ ( .D(n442), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[1])
         );
  fd2qd1_hd r_add_A_reg_31_ ( .D(n447), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_A[31]) );
  fd2qd1_hd r_add_A_reg_0_ ( .D(n448), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_A[0])
         );
  fd2qd1_hd r_y_data_reg_0_ ( .D(n143), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[0]) );
  fd2qd1_hd r_y_data_reg_1_ ( .D(n142), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[1]) );
  fd2qd1_hd r_y_data_reg_2_ ( .D(n141), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[2]) );
  fd2qd1_hd r_y_data_reg_3_ ( .D(n140), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[3]) );
  fd2qd1_hd r_y_data_reg_4_ ( .D(n139), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[4]) );
  fd2qd1_hd r_y_data_reg_5_ ( .D(n138), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[5]) );
  fd2qd1_hd r_y_data_reg_6_ ( .D(n137), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[6]) );
  fd2qd1_hd r_y_data_reg_7_ ( .D(n136), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[7]) );
  fd2qd1_hd r_y_data_reg_8_ ( .D(n135), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[8]) );
  fd2qd1_hd r_y_data_reg_9_ ( .D(n134), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[9]) );
  fd2qd1_hd r_y_data_reg_10_ ( .D(n133), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[10]) );
  fd2qd1_hd r_y_data_reg_11_ ( .D(n132), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[11]) );
  fd2qd1_hd r_y_data_reg_12_ ( .D(n131), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[12]) );
  fd2qd1_hd r_y_data_reg_13_ ( .D(n130), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[13]) );
  fd2qd1_hd r_y_data_reg_14_ ( .D(n129), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[14]) );
  fd2qd1_hd r_y_data_reg_15_ ( .D(n128), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[15]) );
  fd2qd1_hd r_y_data_reg_16_ ( .D(n127), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[16]) );
  fd2qd1_hd r_y_data_reg_17_ ( .D(n126), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[17]) );
  fd2qd1_hd r_y_data_reg_18_ ( .D(n125), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[18]) );
  fd2qd1_hd r_y_data_reg_19_ ( .D(n124), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[19]) );
  fd2qd1_hd r_y_data_reg_20_ ( .D(n123), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[20]) );
  fd2qd1_hd r_y_data_reg_21_ ( .D(n122), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[21]) );
  fd2qd1_hd r_y_data_reg_22_ ( .D(n121), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[22]) );
  fd2qd1_hd r_y_data_reg_23_ ( .D(n120), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[23]) );
  fd2qd1_hd r_y_data_reg_24_ ( .D(n119), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[24]) );
  fd2qd1_hd r_y_data_reg_25_ ( .D(n118), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[25]) );
  fd2qd1_hd r_y_data_reg_26_ ( .D(n117), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[26]) );
  fd2qd1_hd r_y_data_reg_27_ ( .D(n116), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[27]) );
  fd2qd1_hd r_y_data_reg_28_ ( .D(n115), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[28]) );
  fd2qd1_hd r_y_data_reg_29_ ( .D(n114), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[29]) );
  fd2qd1_hd r_y_data_reg_30_ ( .D(n113), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[30]) );
  fd2qd1_hd r_y_data_reg_31_ ( .D(n112), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_y_data[31]) );
  fd2qd1_hd r_add_B_reg_31_ ( .D(n348), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[31]) );
  fd2qd1_hd r_add_B_reg_30_ ( .D(n349), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[30]) );
  fd2qd1_hd r_add_B_reg_29_ ( .D(n350), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[29]) );
  fd2qd1_hd r_add_B_reg_28_ ( .D(n351), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[28]) );
  fd2qd1_hd r_add_B_reg_27_ ( .D(n352), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[27]) );
  fd2qd1_hd r_add_B_reg_26_ ( .D(n353), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[26]) );
  fd2qd1_hd r_add_B_reg_25_ ( .D(n354), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[25]) );
  fd2qd1_hd r_add_B_reg_24_ ( .D(n355), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[24]) );
  fd2qd1_hd r_add_B_reg_23_ ( .D(n356), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[23]) );
  fd2qd1_hd r_add_B_reg_22_ ( .D(n357), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[22]) );
  fd2qd1_hd r_add_B_reg_21_ ( .D(n358), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[21]) );
  fd2qd1_hd r_add_B_reg_20_ ( .D(n359), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[20]) );
  fd2qd1_hd r_add_B_reg_19_ ( .D(n360), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[19]) );
  fd2qd1_hd r_add_B_reg_18_ ( .D(n361), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[18]) );
  fd2qd1_hd r_add_B_reg_17_ ( .D(n362), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[17]) );
  fd2qd1_hd r_add_B_reg_16_ ( .D(n363), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[16]) );
  fd2qd1_hd r_add_B_reg_15_ ( .D(n364), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[15]) );
  fd2qd1_hd r_add_B_reg_14_ ( .D(n365), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[14]) );
  fd2qd1_hd r_add_B_reg_13_ ( .D(n366), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[13]) );
  fd2qd1_hd r_add_B_reg_12_ ( .D(n367), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[12]) );
  fd2qd1_hd r_add_B_reg_11_ ( .D(n368), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[11]) );
  fd2qd1_hd r_add_B_reg_10_ ( .D(n369), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_B[10]) );
  fd2qd1_hd r_add_B_reg_9_ ( .D(n370), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[9])
         );
  fd2qd1_hd r_add_B_reg_8_ ( .D(n371), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[8])
         );
  fd2qd1_hd r_add_B_reg_7_ ( .D(n372), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[7])
         );
  fd2qd1_hd r_add_B_reg_6_ ( .D(n373), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[6])
         );
  fd2qd1_hd r_add_B_reg_5_ ( .D(n374), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[5])
         );
  fd2qd1_hd r_add_B_reg_4_ ( .D(n375), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[4])
         );
  fd2qd1_hd r_add_B_reg_3_ ( .D(n376), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[3])
         );
  fd2qd1_hd r_add_B_reg_2_ ( .D(n377), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[2])
         );
  fd2qd1_hd r_add_B_reg_1_ ( .D(n378), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[1])
         );
  fd2qd1_hd r_add_B_reg_0_ ( .D(n379), .CK(i_CLK), .RN(i_RSTN), .Q(r_add_B[0])
         );
  fd2qd1_hd r_x_data_reg_32_ ( .D(n177), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[32]) );
  fd2qd1_hd r_x_data_reg_33_ ( .D(n176), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[33]) );
  fd2qd1_hd r_x_data_reg_34_ ( .D(n175), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[34]) );
  fd2qd1_hd r_x_data_reg_35_ ( .D(n174), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[35]) );
  fd2qd1_hd r_x_data_reg_36_ ( .D(n173), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[36]) );
  fd2qd1_hd r_x_data_reg_37_ ( .D(n172), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[37]) );
  fd2qd1_hd r_x_data_reg_38_ ( .D(n171), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[38]) );
  fd2qd1_hd r_x_data_reg_39_ ( .D(n170), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[39]) );
  fd2qd1_hd r_x_data_reg_40_ ( .D(n169), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[40]) );
  fd2qd1_hd r_x_data_reg_41_ ( .D(n168), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[41]) );
  fd2qd1_hd r_x_data_reg_42_ ( .D(n167), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[42]) );
  fd2qd1_hd r_x_data_reg_43_ ( .D(n166), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[43]) );
  fd2qd1_hd r_x_data_reg_44_ ( .D(n165), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[44]) );
  fd2qd1_hd r_x_data_reg_45_ ( .D(n164), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[45]) );
  fd2qd1_hd r_x_data_reg_46_ ( .D(n163), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[46]) );
  fd2qd1_hd r_x_data_reg_47_ ( .D(n162), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[47]) );
  fd2qd1_hd r_x_data_reg_48_ ( .D(n161), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[48]) );
  fd2qd1_hd r_x_data_reg_49_ ( .D(n160), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[49]) );
  fd2qd1_hd r_x_data_reg_50_ ( .D(n159), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[50]) );
  fd2qd1_hd r_x_data_reg_51_ ( .D(n158), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[51]) );
  fd2qd1_hd r_x_data_reg_52_ ( .D(n157), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[52]) );
  fd2qd1_hd r_x_data_reg_53_ ( .D(n156), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[53]) );
  fd2qd1_hd r_x_data_reg_54_ ( .D(n155), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[54]) );
  fd2qd1_hd r_x_data_reg_55_ ( .D(n154), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[55]) );
  fd2qd1_hd r_x_data_reg_56_ ( .D(n153), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[56]) );
  fd2qd1_hd r_x_data_reg_57_ ( .D(n152), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[57]) );
  fd2qd1_hd r_x_data_reg_58_ ( .D(n151), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[58]) );
  fd2qd1_hd r_x_data_reg_59_ ( .D(n150), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[59]) );
  fd2qd1_hd r_x_data_reg_60_ ( .D(n149), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[60]) );
  fd2qd1_hd r_x_data_reg_61_ ( .D(n148), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[61]) );
  fd2qd1_hd r_x_data_reg_62_ ( .D(n147), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[62]) );
  fd2qd1_hd r_x_data_reg_63_ ( .D(n146), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[63]) );
  fd2qd1_hd o_Y_DATA_reg_0_ ( .D(n411), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[0]) );
  fd2qd1_hd o_Y_DATA_reg_1_ ( .D(n410), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[1]) );
  fd2qd1_hd o_Y_DATA_reg_2_ ( .D(n409), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[2]) );
  fd2qd1_hd o_Y_DATA_reg_3_ ( .D(n408), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[3]) );
  fd2qd1_hd o_Y_DATA_reg_4_ ( .D(n407), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[4]) );
  fd2qd1_hd o_Y_DATA_reg_5_ ( .D(n406), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[5]) );
  fd2qd1_hd o_Y_DATA_reg_6_ ( .D(n405), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[6]) );
  fd2qd1_hd o_Y_DATA_reg_7_ ( .D(n404), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[7]) );
  fd2qd1_hd o_Y_DATA_reg_8_ ( .D(n403), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[8]) );
  fd2qd1_hd o_Y_DATA_reg_9_ ( .D(n402), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[9]) );
  fd2qd1_hd o_Y_DATA_reg_10_ ( .D(n401), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[10]) );
  fd2qd1_hd o_Y_DATA_reg_11_ ( .D(n400), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[11]) );
  fd2qd1_hd o_Y_DATA_reg_12_ ( .D(n399), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[12]) );
  fd2qd1_hd o_Y_DATA_reg_13_ ( .D(n398), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[13]) );
  fd2qd1_hd o_Y_DATA_reg_14_ ( .D(n397), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[14]) );
  fd2qd1_hd o_Y_DATA_reg_15_ ( .D(n396), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[15]) );
  fd2qd1_hd o_Y_DATA_reg_16_ ( .D(n395), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[16]) );
  fd2qd1_hd o_Y_DATA_reg_17_ ( .D(n394), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[17]) );
  fd2qd1_hd o_Y_DATA_reg_18_ ( .D(n393), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[18]) );
  fd2qd1_hd o_Y_DATA_reg_19_ ( .D(n392), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[19]) );
  fd2qd1_hd o_Y_DATA_reg_20_ ( .D(n391), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[20]) );
  fd2qd1_hd o_Y_DATA_reg_21_ ( .D(n390), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[21]) );
  fd2qd1_hd o_Y_DATA_reg_22_ ( .D(n389), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[22]) );
  fd2qd1_hd o_Y_DATA_reg_23_ ( .D(n388), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[23]) );
  fd2qd1_hd o_Y_DATA_reg_24_ ( .D(n387), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[24]) );
  fd2qd1_hd o_Y_DATA_reg_25_ ( .D(n386), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[25]) );
  fd2qd1_hd o_Y_DATA_reg_26_ ( .D(n385), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[26]) );
  fd2qd1_hd o_Y_DATA_reg_27_ ( .D(n384), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[27]) );
  fd2qd1_hd o_Y_DATA_reg_28_ ( .D(n383), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[28]) );
  fd2qd1_hd o_Y_DATA_reg_29_ ( .D(n382), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[29]) );
  fd2qd1_hd o_Y_DATA_reg_30_ ( .D(n381), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[30]) );
  fd2qd1_hd r_x_data_reg_0_ ( .D(n209), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[0]) );
  fd2qd1_hd r_x_data_reg_1_ ( .D(n208), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[1]) );
  fd2qd1_hd r_x_data_reg_2_ ( .D(n207), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[2]) );
  fd2qd1_hd r_x_data_reg_3_ ( .D(n206), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[3]) );
  fd2qd1_hd r_x_data_reg_4_ ( .D(n205), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[4]) );
  fd2qd1_hd r_x_data_reg_5_ ( .D(n204), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[5]) );
  fd2qd1_hd r_x_data_reg_6_ ( .D(n203), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[6]) );
  fd2qd1_hd r_x_data_reg_7_ ( .D(n202), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[7]) );
  fd2qd1_hd r_x_data_reg_8_ ( .D(n201), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[8]) );
  fd2qd1_hd r_x_data_reg_9_ ( .D(n200), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[9]) );
  fd2qd1_hd r_x_data_reg_10_ ( .D(n199), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[10]) );
  fd2qd1_hd r_x_data_reg_11_ ( .D(n198), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[11]) );
  fd2qd1_hd r_x_data_reg_12_ ( .D(n197), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[12]) );
  fd2qd1_hd r_x_data_reg_13_ ( .D(n196), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[13]) );
  fd2qd1_hd r_x_data_reg_14_ ( .D(n195), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[14]) );
  fd2qd1_hd r_x_data_reg_15_ ( .D(n194), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[15]) );
  fd2qd1_hd r_x_data_reg_16_ ( .D(n193), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[16]) );
  fd2qd1_hd r_x_data_reg_17_ ( .D(n192), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[17]) );
  fd2qd1_hd r_x_data_reg_18_ ( .D(n191), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[18]) );
  fd2qd1_hd r_x_data_reg_19_ ( .D(n190), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[19]) );
  fd2qd1_hd r_x_data_reg_20_ ( .D(n189), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[20]) );
  fd2qd1_hd r_x_data_reg_21_ ( .D(n188), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[21]) );
  fd2qd1_hd r_x_data_reg_22_ ( .D(n187), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[22]) );
  fd2qd1_hd r_x_data_reg_23_ ( .D(n186), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[23]) );
  fd2qd1_hd r_x_data_reg_24_ ( .D(n185), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[24]) );
  fd2qd1_hd r_x_data_reg_25_ ( .D(n184), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[25]) );
  fd2qd1_hd r_x_data_reg_26_ ( .D(n183), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[26]) );
  fd2qd1_hd r_x_data_reg_27_ ( .D(n182), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[27]) );
  fd2qd1_hd r_x_data_reg_28_ ( .D(n181), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[28]) );
  fd2qd1_hd r_x_data_reg_29_ ( .D(n180), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[29]) );
  fd2qd1_hd r_x_data_reg_30_ ( .D(n179), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[30]) );
  fd2qd1_hd r_x_data_reg_31_ ( .D(n178), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_x_data[31]) );
  fd2qd1_hd o_Y_DATA_reg_31_ ( .D(n380), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA[31]) );
  fd1eqd1_hd o_X_DATA_READY_reg ( .D(n450), .E(N559), .CK(i_CLK), .Q(
        o_X_DATA_READY) );
  fd2qd1_hd r_add_Z_ACK_reg ( .D(n443), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_Z_ACK) );
  fd2qd1_hd o_Y_DATA_VALID_reg ( .D(n444), .CK(i_CLK), .RN(i_RSTN), .Q(
        o_Y_DATA_VALID) );
  fd2qd1_hd r_add_AB_STB_reg ( .D(n412), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_add_AB_STB) );
  fd2qd1_hd r_pstate_reg_0_ ( .D(N553), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_pstate_0_) );
  ao22d1_hd U533 ( .A(w_add_Z[12]), .B(n6), .C(r_mult_B[12]), .D(n668), .Y(
        n666) );
  ao22d1_hd U535 ( .A(w_add_Z[13]), .B(n6), .C(r_mult_B[13]), .D(n5), .Y(n669)
         );
  ao22d1_hd U537 ( .A(w_add_Z[14]), .B(n6), .C(r_mult_B[14]), .D(n5), .Y(n670)
         );
  ao22d1_hd U539 ( .A(w_add_Z[15]), .B(n667), .C(r_mult_B[15]), .D(n668), .Y(
        n671) );
  ao22d1_hd U541 ( .A(w_add_Z[16]), .B(n667), .C(r_mult_B[16]), .D(n668), .Y(
        n672) );
  ao22d1_hd U543 ( .A(w_add_Z[17]), .B(n667), .C(r_mult_B[17]), .D(n668), .Y(
        n673) );
  ao22d1_hd U545 ( .A(w_add_Z[18]), .B(n667), .C(r_mult_B[18]), .D(n668), .Y(
        n674) );
  ao22d1_hd U547 ( .A(w_add_Z[19]), .B(n667), .C(r_mult_B[19]), .D(n668), .Y(
        n675) );
  ao22d1_hd U549 ( .A(w_add_Z[20]), .B(n667), .C(r_mult_B[20]), .D(n5), .Y(
        n676) );
  ao22d1_hd U551 ( .A(w_add_Z[21]), .B(n6), .C(r_mult_B[21]), .D(n5), .Y(n677)
         );
  ao22d1_hd U553 ( .A(w_add_Z[22]), .B(n6), .C(r_mult_B[22]), .D(n5), .Y(n678)
         );
  ao22d1_hd U555 ( .A(w_add_Z[23]), .B(n6), .C(r_mult_B[23]), .D(n5), .Y(n679)
         );
  ao22d1_hd U557 ( .A(w_add_Z[24]), .B(n6), .C(r_mult_B[24]), .D(n668), .Y(
        n680) );
  ao22d1_hd U559 ( .A(w_add_Z[25]), .B(n6), .C(r_mult_B[25]), .D(n5), .Y(n681)
         );
  ao22d1_hd U561 ( .A(w_add_Z[26]), .B(n6), .C(r_mult_B[26]), .D(n668), .Y(
        n682) );
  ao22d1_hd U563 ( .A(w_add_Z[27]), .B(n6), .C(r_mult_B[27]), .D(n5), .Y(n683)
         );
  ao22d1_hd U565 ( .A(w_add_Z[28]), .B(n6), .C(r_mult_B[28]), .D(n5), .Y(n684)
         );
  ao22d1_hd U567 ( .A(w_add_Z[29]), .B(n6), .C(r_mult_B[29]), .D(n5), .Y(n685)
         );
  ao22d1_hd U569 ( .A(w_add_Z[30]), .B(n6), .C(r_mult_B[30]), .D(n5), .Y(n686)
         );
  nd2bd1_hd U570 ( .AN(r_mult_A[0]), .B(n687), .Y(n80) );
  nd2bd1_hd U571 ( .AN(r_mult_A[1]), .B(n687), .Y(n79) );
  ad2d1_hd U572 ( .A(r_mult_A[2]), .B(n5), .Y(n78) );
  ad2d1_hd U573 ( .A(r_mult_A[3]), .B(n5), .Y(n77) );
  ad2d1_hd U574 ( .A(r_mult_A[4]), .B(n5), .Y(n76) );
  nd2bd1_hd U575 ( .AN(r_mult_A[5]), .B(n687), .Y(n75) );
  nd2bd1_hd U576 ( .AN(r_mult_A[6]), .B(n687), .Y(n74) );
  nd2bd1_hd U577 ( .AN(r_mult_A[7]), .B(n687), .Y(n73) );
  nd2bd1_hd U578 ( .AN(r_mult_A[8]), .B(n687), .Y(n72) );
  nd2bd1_hd U579 ( .AN(r_mult_A[9]), .B(n687), .Y(n71) );
  ad2d1_hd U580 ( .A(r_mult_A[10]), .B(n5), .Y(n70) );
  nd2bd1_hd U581 ( .AN(r_mult_A[11]), .B(n687), .Y(n69) );
  ad2d1_hd U582 ( .A(r_mult_A[12]), .B(n5), .Y(n68) );
  nd2bd1_hd U583 ( .AN(r_mult_A[13]), .B(n687), .Y(n67) );
  nd2bd1_hd U584 ( .AN(r_mult_A[14]), .B(n687), .Y(n66) );
  ad2d1_hd U585 ( .A(r_mult_A[15]), .B(n5), .Y(n65) );
  nd2bd1_hd U586 ( .AN(r_mult_A[16]), .B(n687), .Y(n64) );
  nd2bd1_hd U587 ( .AN(r_mult_A[17]), .B(n687), .Y(n63) );
  ad2d1_hd U588 ( .A(r_mult_A[18]), .B(n5), .Y(n62) );
  ad2d1_hd U589 ( .A(r_mult_A[19]), .B(n5), .Y(n61) );
  ad2d1_hd U590 ( .A(r_mult_A[20]), .B(n5), .Y(n60) );
  nd2bd1_hd U591 ( .AN(r_mult_A[21]), .B(n687), .Y(n59) );
  nd2bd1_hd U592 ( .AN(r_mult_A[22]), .B(n687), .Y(n58) );
  ad2d1_hd U593 ( .A(r_mult_A[23]), .B(n5), .Y(n57) );
  nd2bd1_hd U594 ( .AN(r_mult_A[24]), .B(n687), .Y(n56) );
  nd2bd1_hd U595 ( .AN(r_mult_A[25]), .B(n687), .Y(n55) );
  nd2bd1_hd U596 ( .AN(r_mult_A[26]), .B(n687), .Y(n54) );
  nd2bd1_hd U597 ( .AN(r_mult_A[27]), .B(n687), .Y(n53) );
  nd2bd1_hd U598 ( .AN(r_mult_A[28]), .B(n687), .Y(n52) );
  nd2bd1_hd U599 ( .AN(r_mult_A[29]), .B(n687), .Y(n51) );
  ad2d1_hd U601 ( .A(r_mult_A[30]), .B(n5), .Y(n50) );
  ad2d1_hd U602 ( .A(r_mult_A[31]), .B(n5), .Y(n49) );
  ao22d1_hd U604 ( .A(w_mult_Z[0]), .B(n4), .C(r_add_A[0]), .D(n3), .Y(n688)
         );
  ao22d1_hd U606 ( .A(w_mult_Z[31]), .B(n4), .C(r_add_A[31]), .D(n3), .Y(n691)
         );
  ao22d1_hd U612 ( .A(w_mult_Z[1]), .B(n4), .C(r_add_A[1]), .D(n3), .Y(n699)
         );
  ao22d1_hd U614 ( .A(w_mult_Z[2]), .B(n4), .C(r_add_A[2]), .D(n3), .Y(n700)
         );
  ao22d1_hd U616 ( .A(w_mult_Z[3]), .B(n4), .C(r_add_A[3]), .D(n3), .Y(n701)
         );
  ao22d1_hd U618 ( .A(w_mult_Z[4]), .B(n4), .C(r_add_A[4]), .D(n3), .Y(n702)
         );
  ao22d1_hd U620 ( .A(w_mult_Z[5]), .B(n4), .C(r_add_A[5]), .D(n3), .Y(n703)
         );
  ao22d1_hd U622 ( .A(w_mult_Z[6]), .B(n4), .C(r_add_A[6]), .D(n3), .Y(n704)
         );
  ao22d1_hd U624 ( .A(w_mult_Z[7]), .B(n4), .C(r_add_A[7]), .D(n3), .Y(n705)
         );
  ao22d1_hd U626 ( .A(w_mult_Z[8]), .B(n4), .C(r_add_A[8]), .D(n3), .Y(n706)
         );
  ao22d1_hd U628 ( .A(w_mult_Z[9]), .B(n4), .C(r_add_A[9]), .D(n3), .Y(n707)
         );
  ao22d1_hd U630 ( .A(w_mult_Z[10]), .B(n4), .C(r_add_A[10]), .D(n3), .Y(n708)
         );
  ao22d1_hd U632 ( .A(w_mult_Z[11]), .B(n4), .C(r_add_A[11]), .D(n3), .Y(n709)
         );
  ao22d1_hd U634 ( .A(w_mult_Z[12]), .B(n4), .C(r_add_A[12]), .D(n3), .Y(n710)
         );
  ao22d1_hd U636 ( .A(w_mult_Z[13]), .B(n4), .C(r_add_A[13]), .D(n3), .Y(n711)
         );
  ao22d1_hd U638 ( .A(w_mult_Z[14]), .B(n4), .C(r_add_A[14]), .D(n3), .Y(n712)
         );
  ao22d1_hd U640 ( .A(w_mult_Z[15]), .B(n4), .C(r_add_A[15]), .D(n3), .Y(n713)
         );
  ao22d1_hd U642 ( .A(w_mult_Z[16]), .B(n4), .C(r_add_A[16]), .D(n3), .Y(n714)
         );
  ao22d1_hd U644 ( .A(w_mult_Z[17]), .B(n4), .C(r_add_A[17]), .D(n3), .Y(n715)
         );
  ao22d1_hd U646 ( .A(w_mult_Z[18]), .B(n4), .C(r_add_A[18]), .D(n3), .Y(n716)
         );
  ao22d1_hd U648 ( .A(w_mult_Z[19]), .B(n4), .C(r_add_A[19]), .D(n3), .Y(n717)
         );
  ao22d1_hd U650 ( .A(w_mult_Z[20]), .B(n4), .C(r_add_A[20]), .D(n3), .Y(n718)
         );
  ao22d1_hd U652 ( .A(w_mult_Z[21]), .B(n4), .C(r_add_A[21]), .D(n3), .Y(n719)
         );
  ao22d1_hd U654 ( .A(w_mult_Z[22]), .B(n4), .C(r_add_A[22]), .D(n3), .Y(n720)
         );
  ao22d1_hd U656 ( .A(w_mult_Z[23]), .B(n4), .C(r_add_A[23]), .D(n3), .Y(n721)
         );
  ao22d1_hd U658 ( .A(w_mult_Z[24]), .B(n4), .C(r_add_A[24]), .D(n3), .Y(n722)
         );
  ao22d1_hd U660 ( .A(w_mult_Z[25]), .B(n4), .C(r_add_A[25]), .D(n3), .Y(n723)
         );
  ao22d1_hd U662 ( .A(w_mult_Z[26]), .B(n4), .C(r_add_A[26]), .D(n3), .Y(n724)
         );
  ao22d1_hd U664 ( .A(w_mult_Z[27]), .B(n4), .C(r_add_A[27]), .D(n3), .Y(n725)
         );
  ao22d1_hd U666 ( .A(w_mult_Z[28]), .B(n4), .C(r_add_A[28]), .D(n3), .Y(n726)
         );
  ao22d1_hd U668 ( .A(w_mult_Z[29]), .B(n4), .C(r_add_A[29]), .D(n3), .Y(n727)
         );
  ao22d1_hd U670 ( .A(w_mult_Z[30]), .B(n4), .C(r_add_A[30]), .D(n3), .Y(n728)
         );
  ao22d1_hd U674 ( .A(n734), .B(w_mult_Z[0]), .C(n735), .D(w_add_Z[0]), .Y(
        n733) );
  ao22d1_hd U676 ( .A(n734), .B(w_mult_Z[1]), .C(n735), .D(w_add_Z[1]), .Y(
        n736) );
  ao22d1_hd U678 ( .A(n734), .B(w_mult_Z[2]), .C(n735), .D(w_add_Z[2]), .Y(
        n737) );
  ao22d1_hd U680 ( .A(n734), .B(w_mult_Z[3]), .C(n735), .D(w_add_Z[3]), .Y(
        n738) );
  ao22d1_hd U682 ( .A(n734), .B(w_mult_Z[4]), .C(n735), .D(w_add_Z[4]), .Y(
        n739) );
  ao22d1_hd U684 ( .A(n734), .B(w_mult_Z[5]), .C(n735), .D(w_add_Z[5]), .Y(
        n740) );
  ao22d1_hd U686 ( .A(n734), .B(w_mult_Z[6]), .C(n735), .D(w_add_Z[6]), .Y(
        n741) );
  ao22d1_hd U688 ( .A(n734), .B(w_mult_Z[7]), .C(n735), .D(w_add_Z[7]), .Y(
        n742) );
  ao22d1_hd U690 ( .A(n734), .B(w_mult_Z[8]), .C(n735), .D(w_add_Z[8]), .Y(
        n743) );
  ao22d1_hd U692 ( .A(n734), .B(w_mult_Z[9]), .C(n735), .D(w_add_Z[9]), .Y(
        n744) );
  ao22d1_hd U694 ( .A(n734), .B(w_mult_Z[10]), .C(n735), .D(w_add_Z[10]), .Y(
        n745) );
  ao22d1_hd U696 ( .A(n734), .B(w_mult_Z[11]), .C(n735), .D(w_add_Z[11]), .Y(
        n746) );
  ao22d1_hd U698 ( .A(n734), .B(w_mult_Z[12]), .C(n735), .D(w_add_Z[12]), .Y(
        n747) );
  ao22d1_hd U700 ( .A(n734), .B(w_mult_Z[13]), .C(n735), .D(w_add_Z[13]), .Y(
        n748) );
  ao22d1_hd U702 ( .A(n734), .B(w_mult_Z[14]), .C(n735), .D(w_add_Z[14]), .Y(
        n749) );
  ao22d1_hd U704 ( .A(n734), .B(w_mult_Z[15]), .C(n735), .D(w_add_Z[15]), .Y(
        n750) );
  ao22d1_hd U706 ( .A(n734), .B(w_mult_Z[16]), .C(n735), .D(w_add_Z[16]), .Y(
        n751) );
  ao22d1_hd U708 ( .A(n734), .B(w_mult_Z[17]), .C(n735), .D(w_add_Z[17]), .Y(
        n752) );
  ao22d1_hd U710 ( .A(n734), .B(w_mult_Z[18]), .C(n735), .D(w_add_Z[18]), .Y(
        n753) );
  ao22d1_hd U712 ( .A(n734), .B(w_mult_Z[19]), .C(n735), .D(w_add_Z[19]), .Y(
        n754) );
  ao22d1_hd U714 ( .A(n734), .B(w_mult_Z[20]), .C(n735), .D(w_add_Z[20]), .Y(
        n755) );
  ao22d1_hd U716 ( .A(n734), .B(w_mult_Z[21]), .C(n735), .D(w_add_Z[21]), .Y(
        n756) );
  ao22d1_hd U718 ( .A(n734), .B(w_mult_Z[22]), .C(n735), .D(w_add_Z[22]), .Y(
        n757) );
  ao22d1_hd U720 ( .A(n734), .B(w_mult_Z[23]), .C(n735), .D(w_add_Z[23]), .Y(
        n758) );
  ao22d1_hd U722 ( .A(n734), .B(w_mult_Z[24]), .C(n735), .D(w_add_Z[24]), .Y(
        n759) );
  ao22d1_hd U724 ( .A(n734), .B(w_mult_Z[25]), .C(n735), .D(w_add_Z[25]), .Y(
        n760) );
  ao22d1_hd U726 ( .A(n734), .B(w_mult_Z[26]), .C(n735), .D(w_add_Z[26]), .Y(
        n761) );
  ao22d1_hd U728 ( .A(n734), .B(w_mult_Z[27]), .C(n735), .D(w_add_Z[27]), .Y(
        n762) );
  ao22d1_hd U730 ( .A(n734), .B(w_mult_Z[28]), .C(n735), .D(w_add_Z[28]), .Y(
        n763) );
  ao22d1_hd U732 ( .A(n734), .B(w_mult_Z[29]), .C(n735), .D(w_add_Z[29]), .Y(
        n764) );
  ao22d1_hd U734 ( .A(n734), .B(w_mult_Z[30]), .C(n735), .D(w_add_Z[30]), .Y(
        n765) );
  ao22d1_hd U736 ( .A(w_mult_Z[31]), .B(n734), .C(n735), .D(w_add_Z[31]), .Y(
        n766) );
  ao22d1_hd U807 ( .A(w_add_Z[31]), .B(n6), .C(r_mult_B[31]), .D(n668), .Y(
        n801) );
  ao22d1_hd U883 ( .A(n695), .B(n804), .C(r_mult_Z_ACK), .D(n595), .Y(n810) );
  ao22d1_hd U917 ( .A(w_add_Z[0]), .B(n6), .C(r_mult_B[0]), .D(n668), .Y(n811)
         );
  ao22d1_hd U919 ( .A(w_add_Z[1]), .B(n6), .C(r_mult_B[1]), .D(n5), .Y(n812)
         );
  ao22d1_hd U921 ( .A(w_add_Z[2]), .B(n6), .C(r_mult_B[2]), .D(n668), .Y(n813)
         );
  ao22d1_hd U923 ( .A(w_add_Z[3]), .B(n6), .C(r_mult_B[3]), .D(n5), .Y(n814)
         );
  ao22d1_hd U925 ( .A(w_add_Z[4]), .B(n6), .C(r_mult_B[4]), .D(n5), .Y(n815)
         );
  ao22d1_hd U927 ( .A(w_add_Z[5]), .B(n6), .C(r_mult_B[5]), .D(n5), .Y(n816)
         );
  ao22d1_hd U929 ( .A(w_add_Z[6]), .B(n6), .C(r_mult_B[6]), .D(n668), .Y(n817)
         );
  ao22d1_hd U931 ( .A(w_add_Z[7]), .B(n6), .C(r_mult_B[7]), .D(n5), .Y(n818)
         );
  ao22d1_hd U933 ( .A(w_add_Z[8]), .B(n6), .C(r_mult_B[8]), .D(n5), .Y(n819)
         );
  ao22d1_hd U935 ( .A(w_add_Z[9]), .B(n6), .C(r_mult_B[9]), .D(n5), .Y(n820)
         );
  ao22d1_hd U937 ( .A(w_add_Z[10]), .B(n6), .C(r_mult_B[10]), .D(n5), .Y(n821)
         );
  ao22d1_hd U939 ( .A(w_add_Z[11]), .B(n6), .C(r_mult_B[11]), .D(n5), .Y(n822)
         );
  nd4d1_hd U942 ( .A(n221), .B(n223), .C(w_mult_AB_ACK), .D(w_add_AB_ACK), .Y(
        n823) );
  oa211d1_hd U954 ( .A(w_mult_Z_STB), .B(n597), .C(n223), .D(w_add_Z_STB), .Y(
        n826) );
  scg14d1_hd U956 ( .A(w_mult_AB_ACK), .B(w_add_AB_ACK), .C(n694), .Y(n825) );
  nd3d1_hd U955 ( .A(n221), .B(w_mult_Z_STB), .C(n598), .Y(n803) );
  scg12d1_hd U945 ( .A(w_mult_Z_STB), .B(w_add_Z_STB), .C(n597), .Y(n804) );
  oa211d1_hd U740 ( .A(w_mult_Z_STB), .B(n597), .C(w_add_Z_STB), .D(n698), .Y(
        n767) );
  nd3d1_hd U949 ( .A(n694), .B(w_mult_AB_ACK), .C(w_add_AB_ACK), .Y(n731) );
  ivd6_hd U457 ( .A(n450), .Y(n1) );
  clknd2d1_hd U458 ( .A(n213), .B(n220), .Y(n8) );
  clknd2d1_hd U459 ( .A(r_pstate_0_), .B(n213), .Y(n595) );
  nid2_hd U460 ( .A(n667), .Y(n6) );
  clknd2d1_hd U461 ( .A(n221), .B(n226), .Y(n294) );
  clknd2d1_hd U462 ( .A(r_add_AB_STB), .B(n294), .Y(n295) );
  nd2d4_hd U463 ( .A(i_X_DATA_VALID), .B(o_X_DATA_READY), .Y(n450) );
  clknd2d1_hd U464 ( .A(n1), .B(i_X_DATA[31]), .Y(n22) );
  clknd2d1_hd U465 ( .A(n1), .B(i_X_DATA[30]), .Y(n23) );
  clknd2d1_hd U466 ( .A(n1), .B(i_X_DATA[29]), .Y(n24) );
  clknd2d1_hd U467 ( .A(n1), .B(i_X_DATA[28]), .Y(n25) );
  clknd2d1_hd U468 ( .A(n1), .B(i_X_DATA[27]), .Y(n26) );
  clknd2d1_hd U469 ( .A(n1), .B(i_X_DATA[26]), .Y(n27) );
  clknd2d1_hd U470 ( .A(n1), .B(i_X_DATA[25]), .Y(n28) );
  clknd2d1_hd U471 ( .A(n1), .B(i_X_DATA[24]), .Y(n29) );
  clknd2d1_hd U472 ( .A(n1), .B(i_X_DATA[23]), .Y(n30) );
  clknd2d1_hd U473 ( .A(n1), .B(i_X_DATA[22]), .Y(n31) );
  clknd2d1_hd U474 ( .A(n1), .B(i_X_DATA[21]), .Y(n32) );
  clknd2d1_hd U475 ( .A(n1), .B(i_X_DATA[20]), .Y(n33) );
  clknd2d1_hd U476 ( .A(n1), .B(i_X_DATA[19]), .Y(n34) );
  clknd2d1_hd U477 ( .A(n1), .B(i_X_DATA[18]), .Y(n35) );
  clknd2d1_hd U478 ( .A(n1), .B(i_X_DATA[17]), .Y(n36) );
  clknd2d1_hd U479 ( .A(n1), .B(i_X_DATA[16]), .Y(n37) );
  clknd2d1_hd U480 ( .A(n1), .B(i_X_DATA[15]), .Y(n38) );
  clknd2d1_hd U481 ( .A(n1), .B(i_X_DATA[14]), .Y(n39) );
  clknd2d1_hd U482 ( .A(n1), .B(i_X_DATA[13]), .Y(n40) );
  clknd2d1_hd U483 ( .A(n1), .B(i_X_DATA[12]), .Y(n41) );
  clknd2d1_hd U484 ( .A(n1), .B(i_X_DATA[11]), .Y(n42) );
  clknd2d1_hd U485 ( .A(n1), .B(i_X_DATA[10]), .Y(n43) );
  clknd2d1_hd U486 ( .A(n1), .B(i_X_DATA[9]), .Y(n44) );
  clknd2d1_hd U487 ( .A(n1), .B(i_X_DATA[8]), .Y(n45) );
  clknd2d1_hd U488 ( .A(n1), .B(i_X_DATA[7]), .Y(n46) );
  clknd2d1_hd U489 ( .A(n1), .B(i_X_DATA[6]), .Y(n47) );
  clknd2d1_hd U490 ( .A(n1), .B(i_X_DATA[5]), .Y(n48) );
  clknd2d1_hd U491 ( .A(n1), .B(i_X_DATA[4]), .Y(n215) );
  clknd2d1_hd U492 ( .A(n1), .B(i_X_DATA[3]), .Y(n216) );
  clknd2d1_hd U493 ( .A(n1), .B(i_X_DATA[2]), .Y(n217) );
  clknd2d1_hd U494 ( .A(n1), .B(i_X_DATA[1]), .Y(n218) );
  clknd2d1_hd U495 ( .A(n1), .B(i_X_DATA[0]), .Y(n219) );
  clknd2d1_hd U496 ( .A(n810), .B(n689), .Y(n144) );
  clknd2d1_hd U497 ( .A(r_mult_AB_STB), .B(n594), .Y(n809) );
  nr2d4_hd U498 ( .A(n598), .B(n294), .Y(n332) );
  ivd3_hd U499 ( .A(n689), .Y(n4) );
  ivd6_hd U500 ( .A(n332), .Y(n2) );
  nr2d4_hd U501 ( .A(n221), .B(n767), .Y(n735) );
  scg10d1_hd U502 ( .A(n450), .B(r_x_data[31]), .C(r_x_data[63]), .D(n1), .Y(
        n146) );
  scg10d1_hd U503 ( .A(n450), .B(r_x_data[30]), .C(r_x_data[62]), .D(n1), .Y(
        n147) );
  scg10d1_hd U504 ( .A(n450), .B(r_x_data[29]), .C(r_x_data[61]), .D(n1), .Y(
        n148) );
  scg10d1_hd U505 ( .A(n450), .B(r_x_data[28]), .C(r_x_data[60]), .D(n1), .Y(
        n149) );
  scg10d1_hd U506 ( .A(n450), .B(r_x_data[27]), .C(r_x_data[59]), .D(n1), .Y(
        n150) );
  scg10d1_hd U507 ( .A(n450), .B(r_x_data[26]), .C(r_x_data[58]), .D(n1), .Y(
        n151) );
  scg10d1_hd U508 ( .A(n450), .B(r_x_data[25]), .C(r_x_data[57]), .D(n1), .Y(
        n152) );
  scg10d1_hd U509 ( .A(n450), .B(r_x_data[24]), .C(r_x_data[56]), .D(n1), .Y(
        n153) );
  scg10d1_hd U510 ( .A(n450), .B(r_x_data[23]), .C(r_x_data[55]), .D(n1), .Y(
        n154) );
  scg10d1_hd U511 ( .A(n450), .B(r_x_data[22]), .C(r_x_data[54]), .D(n1), .Y(
        n155) );
  scg10d1_hd U512 ( .A(n450), .B(r_x_data[20]), .C(r_x_data[52]), .D(n1), .Y(
        n157) );
  scg10d1_hd U513 ( .A(n450), .B(r_x_data[19]), .C(r_x_data[51]), .D(n1), .Y(
        n158) );
  scg10d1_hd U514 ( .A(n450), .B(r_x_data[18]), .C(r_x_data[50]), .D(n1), .Y(
        n159) );
  scg10d1_hd U515 ( .A(n450), .B(r_x_data[17]), .C(r_x_data[49]), .D(n1), .Y(
        n160) );
  scg10d1_hd U516 ( .A(n450), .B(r_x_data[16]), .C(r_x_data[48]), .D(n1), .Y(
        n161) );
  scg10d1_hd U517 ( .A(n450), .B(r_x_data[15]), .C(r_x_data[47]), .D(n1), .Y(
        n162) );
  scg10d1_hd U518 ( .A(n450), .B(r_x_data[14]), .C(r_x_data[46]), .D(n1), .Y(
        n163) );
  scg10d1_hd U519 ( .A(n450), .B(r_x_data[13]), .C(r_x_data[45]), .D(n1), .Y(
        n164) );
  scg10d1_hd U520 ( .A(n450), .B(r_x_data[12]), .C(r_x_data[44]), .D(n1), .Y(
        n165) );
  scg10d1_hd U521 ( .A(n450), .B(r_x_data[11]), .C(r_x_data[43]), .D(n1), .Y(
        n166) );
  scg10d1_hd U522 ( .A(n450), .B(r_x_data[10]), .C(r_x_data[42]), .D(n1), .Y(
        n167) );
  scg10d1_hd U523 ( .A(n450), .B(r_x_data[9]), .C(r_x_data[41]), .D(n1), .Y(
        n168) );
  scg10d1_hd U524 ( .A(n450), .B(r_x_data[6]), .C(r_x_data[38]), .D(n1), .Y(
        n171) );
  or2d4_hd U525 ( .A(n803), .B(n594), .Y(n689) );
  ad3d2_hd U526 ( .A(n292), .B(n698), .C(n221), .Y(n734) );
  clknd2d4_hd U527 ( .A(n767), .B(n2), .Y(n292) );
  scg10d1_hd U528 ( .A(n450), .B(r_x_data[7]), .C(r_x_data[39]), .D(n1), .Y(
        n170) );
  scg10d1_hd U529 ( .A(n450), .B(r_x_data[4]), .C(r_x_data[36]), .D(n1), .Y(
        n173) );
  scg10d1_hd U530 ( .A(n450), .B(r_x_data[3]), .C(r_x_data[35]), .D(n1), .Y(
        n174) );
  scg10d1_hd U531 ( .A(n450), .B(r_x_data[8]), .C(r_x_data[40]), .D(n1), .Y(
        n169) );
  scg10d1_hd U532 ( .A(n450), .B(r_x_data[21]), .C(r_x_data[53]), .D(n1), .Y(
        n156) );
  scg10d1_hd U534 ( .A(n450), .B(r_x_data[0]), .C(r_x_data[32]), .D(n1), .Y(
        n177) );
  scg10d1_hd U536 ( .A(n450), .B(r_x_data[5]), .C(r_x_data[37]), .D(n1), .Y(
        n172) );
  scg10d1_hd U538 ( .A(n450), .B(r_x_data[2]), .C(r_x_data[34]), .D(n1), .Y(
        n175) );
  scg10d1_hd U540 ( .A(n450), .B(r_x_data[1]), .C(r_x_data[33]), .D(n1), .Y(
        n176) );
  nr2d4_hd U542 ( .A(n6), .B(n332), .Y(n687) );
  ivd1_hd U544 ( .A(n595), .Y(n694) );
  ivd1_hd U546 ( .A(n695), .Y(n594) );
  ivd1_hd U548 ( .A(n731), .Y(n226) );
  nr2bd1_hd U550 ( .AN(n222), .B(n597), .Y(n225) );
  nid2_hd U552 ( .A(n668), .Y(n5) );
  scg6d1_hd U554 ( .A(n694), .B(n823), .C(n327), .Y(n668) );
  nr2d1_hd U556 ( .A(n327), .B(n594), .Y(n667) );
  nid4_hd U558 ( .A(n690), .Y(n3) );
  scg20d1_hd U560 ( .A(n823), .B(n595), .C(n4), .Y(n690) );
  nr2d1_hd U562 ( .A(n594), .B(n598), .Y(n698) );
  ivd1_hd U564 ( .A(n223), .Y(n598) );
  ivd1_hd U566 ( .A(r_y_data[24]), .Y(n339) );
  ivd1_hd U568 ( .A(r_y_data[20]), .Y(n343) );
  ivd1_hd U600 ( .A(r_y_data[26]), .Y(n337) );
  ivd1_hd U603 ( .A(r_y_data[25]), .Y(n338) );
  ivd1_hd U605 ( .A(r_y_data[14]), .Y(n446) );
  ivd1_hd U607 ( .A(r_y_data[27]), .Y(n336) );
  ivd1_hd U608 ( .A(r_y_data[15]), .Y(n445) );
  ivd1_hd U609 ( .A(r_y_data[19]), .Y(n344) );
  ivd1_hd U610 ( .A(r_y_data[29]), .Y(n334) );
  ivd1_hd U611 ( .A(r_y_data[21]), .Y(n342) );
  ivd1_hd U613 ( .A(r_y_data[13]), .Y(n449) );
  ivd1_hd U615 ( .A(r_y_data[18]), .Y(n345) );
  ivd1_hd U617 ( .A(r_y_data[28]), .Y(n335) );
  ivd1_hd U619 ( .A(r_y_data[22]), .Y(n341) );
  ivd1_hd U621 ( .A(r_y_data[17]), .Y(n346) );
  ivd1_hd U623 ( .A(r_y_data[16]), .Y(n347) );
  ivd1_hd U625 ( .A(r_y_data[30]), .Y(n333) );
  ivd1_hd U627 ( .A(r_y_data[11]), .Y(n9) );
  ao21d1_hd U629 ( .A(n698), .B(n804), .C(n694), .Y(n327) );
  ivd1_hd U631 ( .A(r_x_data[2]), .Y(n324) );
  ivd1_hd U633 ( .A(r_x_data[16]), .Y(n310) );
  ivd1_hd U635 ( .A(r_x_data[15]), .Y(n311) );
  ivd1_hd U637 ( .A(r_x_data[4]), .Y(n322) );
  ivd1_hd U639 ( .A(r_x_data[3]), .Y(n323) );
  ivd1_hd U641 ( .A(r_x_data[0]), .Y(n331) );
  ivd1_hd U643 ( .A(r_x_data[1]), .Y(n325) );
  ivd1_hd U645 ( .A(r_x_data[31]), .Y(n330) );
  ivd1_hd U647 ( .A(r_y_data[31]), .Y(n228) );
  ivd1_hd U649 ( .A(r_y_data[2]), .Y(n18) );
  ivd1_hd U651 ( .A(r_y_data[10]), .Y(n10) );
  ivd1_hd U653 ( .A(r_y_data[6]), .Y(n14) );
  ivd1_hd U655 ( .A(r_x_data[24]), .Y(n302) );
  ivd1_hd U657 ( .A(r_y_data[1]), .Y(n19) );
  ivd1_hd U659 ( .A(r_y_data[7]), .Y(n13) );
  ivd1_hd U661 ( .A(r_y_data[0]), .Y(n20) );
  ivd1_hd U663 ( .A(r_y_data[23]), .Y(n340) );
  ivd1_hd U665 ( .A(r_y_data[5]), .Y(n15) );
  ivd1_hd U667 ( .A(r_y_data[8]), .Y(n12) );
  ivd1_hd U669 ( .A(r_x_data[30]), .Y(n296) );
  ivd1_hd U671 ( .A(r_y_data[4]), .Y(n16) );
  ivd1_hd U672 ( .A(r_x_data[20]), .Y(n306) );
  ivd1_hd U673 ( .A(r_x_data[22]), .Y(n304) );
  ivd1_hd U675 ( .A(r_y_data[3]), .Y(n17) );
  ivd1_hd U677 ( .A(r_x_data[27]), .Y(n299) );
  ivd1_hd U679 ( .A(r_x_data[17]), .Y(n309) );
  ivd1_hd U681 ( .A(r_x_data[25]), .Y(n301) );
  ivd1_hd U683 ( .A(r_x_data[19]), .Y(n307) );
  ivd1_hd U685 ( .A(r_x_data[9]), .Y(n317) );
  ivd1_hd U687 ( .A(r_x_data[10]), .Y(n316) );
  ivd1_hd U689 ( .A(r_x_data[7]), .Y(n319) );
  ivd1_hd U691 ( .A(r_x_data[29]), .Y(n297) );
  ivd1_hd U693 ( .A(r_x_data[14]), .Y(n312) );
  ivd1_hd U695 ( .A(r_x_data[5]), .Y(n321) );
  ivd1_hd U697 ( .A(r_x_data[18]), .Y(n308) );
  ivd1_hd U699 ( .A(r_x_data[23]), .Y(n303) );
  ivd1_hd U701 ( .A(r_x_data[13]), .Y(n313) );
  ivd1_hd U703 ( .A(r_x_data[28]), .Y(n298) );
  ivd1_hd U705 ( .A(r_y_data[12]), .Y(n451) );
  ivd1_hd U707 ( .A(r_x_data[21]), .Y(n305) );
  ivd1_hd U709 ( .A(r_x_data[8]), .Y(n318) );
  ivd1_hd U711 ( .A(r_x_data[6]), .Y(n320) );
  ivd1_hd U713 ( .A(r_x_data[11]), .Y(n315) );
  ivd1_hd U715 ( .A(r_x_data[12]), .Y(n314) );
  ivd1_hd U717 ( .A(r_x_data[26]), .Y(n300) );
  ivd1_hd U719 ( .A(r_y_data[9]), .Y(n11) );
  ivd1_hd U721 ( .A(o_Y_DATA[31]), .Y(n261) );
  ivd1_hd U723 ( .A(o_Y_DATA[24]), .Y(n268) );
  ivd1_hd U725 ( .A(o_Y_DATA[23]), .Y(n269) );
  ivd1_hd U727 ( .A(o_Y_DATA[21]), .Y(n271) );
  ivd1_hd U729 ( .A(o_Y_DATA[22]), .Y(n270) );
  ivd1_hd U731 ( .A(o_Y_DATA[20]), .Y(n272) );
  ivd1_hd U733 ( .A(o_Y_DATA[5]), .Y(n287) );
  ivd1_hd U735 ( .A(o_Y_DATA[7]), .Y(n285) );
  ivd1_hd U737 ( .A(o_Y_DATA[4]), .Y(n288) );
  ivd1_hd U738 ( .A(o_Y_DATA[6]), .Y(n286) );
  ivd1_hd U739 ( .A(o_Y_DATA[3]), .Y(n289) );
  ivd1_hd U741 ( .A(o_Y_DATA[2]), .Y(n290) );
  ivd1_hd U742 ( .A(o_Y_DATA[28]), .Y(n264) );
  ivd1_hd U743 ( .A(o_Y_DATA[27]), .Y(n265) );
  ivd1_hd U744 ( .A(o_Y_DATA[26]), .Y(n266) );
  ivd1_hd U745 ( .A(o_Y_DATA[30]), .Y(n262) );
  ivd1_hd U746 ( .A(o_Y_DATA[29]), .Y(n263) );
  ivd1_hd U747 ( .A(o_Y_DATA[18]), .Y(n274) );
  ivd1_hd U748 ( .A(o_Y_DATA[9]), .Y(n283) );
  ivd1_hd U749 ( .A(o_Y_DATA[10]), .Y(n282) );
  ivd1_hd U750 ( .A(o_Y_DATA[25]), .Y(n267) );
  ivd1_hd U751 ( .A(o_Y_DATA[19]), .Y(n273) );
  ivd1_hd U752 ( .A(o_Y_DATA[11]), .Y(n281) );
  ivd1_hd U753 ( .A(o_Y_DATA[0]), .Y(n293) );
  ivd1_hd U754 ( .A(o_Y_DATA[8]), .Y(n284) );
  ivd1_hd U755 ( .A(o_Y_DATA[1]), .Y(n291) );
  ivd1_hd U756 ( .A(o_Y_DATA[14]), .Y(n278) );
  ivd1_hd U757 ( .A(o_Y_DATA[12]), .Y(n280) );
  ivd1_hd U758 ( .A(o_Y_DATA[13]), .Y(n279) );
  ivd1_hd U759 ( .A(o_Y_DATA[15]), .Y(n277) );
  ivd1_hd U760 ( .A(o_Y_DATA[17]), .Y(n275) );
  nr2d1_hd U761 ( .A(r_pstate_0_), .B(n213), .Y(n695) );
  ivd1_hd U762 ( .A(n221), .Y(n597) );
  ivd1_hd U763 ( .A(o_Y_DATA[16]), .Y(n276) );
  ivd1_hd U764 ( .A(r_pstate_0_), .Y(n220) );
  ao21d1_hd U765 ( .A(n803), .B(n826), .C(n594), .Y(n222) );
  ao211d1_hd U766 ( .A(o_Y_DATA_VALID), .B(i_Y_ACK), .C(n213), .D(n220), .Y(
        n329) );
  nr2d1_hd U767 ( .A(n222), .B(n329), .Y(n7) );
  oa211d1_hd U768 ( .A(n450), .B(n8), .C(n825), .D(n7), .Y(N553) );
  nr2d1_hd U769 ( .A(N17), .B(n8), .Y(N559) );
  oa21d1_hd U770 ( .A(n2), .B(n9), .C(n822), .Y(n100) );
  oa21d1_hd U771 ( .A(n2), .B(n10), .C(n821), .Y(n101) );
  oa21d1_hd U772 ( .A(n2), .B(n11), .C(n820), .Y(n102) );
  oa21d1_hd U773 ( .A(n2), .B(n12), .C(n819), .Y(n103) );
  oa21d1_hd U774 ( .A(n2), .B(n13), .C(n818), .Y(n104) );
  oa21d1_hd U775 ( .A(n2), .B(n14), .C(n817), .Y(n105) );
  oa21d1_hd U776 ( .A(n2), .B(n15), .C(n816), .Y(n106) );
  oa21d1_hd U777 ( .A(n2), .B(n16), .C(n815), .Y(n107) );
  oa21d1_hd U778 ( .A(n2), .B(n17), .C(n814), .Y(n108) );
  oa21d1_hd U779 ( .A(n2), .B(n18), .C(n813), .Y(n109) );
  oa21d1_hd U780 ( .A(n2), .B(n19), .C(n812), .Y(n110) );
  oa21d1_hd U781 ( .A(n2), .B(n20), .C(n811), .Y(n111) );
  ao22d1_hd U782 ( .A(n1), .B(n261), .C(n228), .D(n450), .Y(n112) );
  ao22d1_hd U783 ( .A(n1), .B(n262), .C(n333), .D(n450), .Y(n113) );
  ao22d1_hd U784 ( .A(n1), .B(n263), .C(n334), .D(n450), .Y(n114) );
  ao22d1_hd U785 ( .A(n1), .B(n264), .C(n335), .D(n450), .Y(n115) );
  ao22d1_hd U786 ( .A(n1), .B(n265), .C(n336), .D(n450), .Y(n116) );
  ao22d1_hd U787 ( .A(n1), .B(n266), .C(n337), .D(n450), .Y(n117) );
  ao22d1_hd U788 ( .A(n1), .B(n267), .C(n338), .D(n450), .Y(n118) );
  ao22d1_hd U789 ( .A(n1), .B(n268), .C(n339), .D(n450), .Y(n119) );
  ao22d1_hd U790 ( .A(n1), .B(n269), .C(n340), .D(n450), .Y(n120) );
  ao22d1_hd U791 ( .A(n1), .B(n270), .C(n341), .D(n450), .Y(n121) );
  ao22d1_hd U792 ( .A(n1), .B(n271), .C(n342), .D(n450), .Y(n122) );
  ao22d1_hd U793 ( .A(n1), .B(n272), .C(n343), .D(n450), .Y(n123) );
  ao22d1_hd U794 ( .A(n1), .B(n273), .C(n344), .D(n450), .Y(n124) );
  ao22d1_hd U795 ( .A(n1), .B(n274), .C(n345), .D(n450), .Y(n125) );
  ao22d1_hd U796 ( .A(n1), .B(n275), .C(n346), .D(n450), .Y(n126) );
  ao22d1_hd U797 ( .A(n1), .B(n276), .C(n347), .D(n450), .Y(n127) );
  ao22d1_hd U798 ( .A(n1), .B(n277), .C(n445), .D(n450), .Y(n128) );
  ao22d1_hd U799 ( .A(n1), .B(n278), .C(n446), .D(n450), .Y(n129) );
  ao22d1_hd U800 ( .A(n1), .B(n279), .C(n449), .D(n450), .Y(n130) );
  ao22d1_hd U801 ( .A(n1), .B(n280), .C(n451), .D(n450), .Y(n131) );
  ao22d1_hd U802 ( .A(n1), .B(n281), .C(n9), .D(n450), .Y(n132) );
  ao22d1_hd U803 ( .A(n1), .B(n282), .C(n10), .D(n450), .Y(n133) );
  ao22d1_hd U804 ( .A(n1), .B(n283), .C(n11), .D(n450), .Y(n134) );
  ao22d1_hd U805 ( .A(n1), .B(n284), .C(n12), .D(n450), .Y(n135) );
  ao22d1_hd U806 ( .A(n1), .B(n285), .C(n13), .D(n450), .Y(n136) );
  ao22d1_hd U808 ( .A(n1), .B(n286), .C(n14), .D(n450), .Y(n137) );
  ao22d1_hd U809 ( .A(n1), .B(n287), .C(n15), .D(n450), .Y(n138) );
  ao22d1_hd U810 ( .A(n1), .B(n288), .C(n16), .D(n450), .Y(n139) );
  ao22d1_hd U811 ( .A(n1), .B(n289), .C(n17), .D(n450), .Y(n140) );
  ao22d1_hd U812 ( .A(n1), .B(n290), .C(n18), .D(n450), .Y(n141) );
  ao22d1_hd U813 ( .A(n1), .B(n291), .C(n19), .D(n450), .Y(n142) );
  ao22d1_hd U814 ( .A(n1), .B(n293), .C(n20), .D(n450), .Y(n143) );
  nr2d1_hd U815 ( .A(n731), .B(n598), .Y(n21) );
  oa21d1_hd U816 ( .A(n21), .B(n809), .C(n294), .Y(n145) );
  oa21d1_hd U817 ( .A(n330), .B(n1), .C(n22), .Y(n178) );
  oa21d1_hd U818 ( .A(n296), .B(n1), .C(n23), .Y(n179) );
  oa21d1_hd U819 ( .A(n297), .B(n1), .C(n24), .Y(n180) );
  oa21d1_hd U820 ( .A(n298), .B(n1), .C(n25), .Y(n181) );
  oa21d1_hd U821 ( .A(n299), .B(n1), .C(n26), .Y(n182) );
  oa21d1_hd U822 ( .A(n300), .B(n1), .C(n27), .Y(n183) );
  oa21d1_hd U823 ( .A(n301), .B(n1), .C(n28), .Y(n184) );
  oa21d1_hd U824 ( .A(n302), .B(n1), .C(n29), .Y(n185) );
  oa21d1_hd U825 ( .A(n303), .B(n1), .C(n30), .Y(n186) );
  oa21d1_hd U826 ( .A(n304), .B(n1), .C(n31), .Y(n187) );
  oa21d1_hd U827 ( .A(n305), .B(n1), .C(n32), .Y(n188) );
  oa21d1_hd U828 ( .A(n306), .B(n1), .C(n33), .Y(n189) );
  oa21d1_hd U829 ( .A(n307), .B(n1), .C(n34), .Y(n190) );
  oa21d1_hd U830 ( .A(n308), .B(n1), .C(n35), .Y(n191) );
  oa21d1_hd U831 ( .A(n309), .B(n1), .C(n36), .Y(n192) );
  oa21d1_hd U832 ( .A(n310), .B(n1), .C(n37), .Y(n193) );
  oa21d1_hd U833 ( .A(n311), .B(n1), .C(n38), .Y(n194) );
  oa21d1_hd U834 ( .A(n312), .B(n1), .C(n39), .Y(n195) );
  oa21d1_hd U835 ( .A(n313), .B(n1), .C(n40), .Y(n196) );
  oa21d1_hd U836 ( .A(n314), .B(n1), .C(n41), .Y(n197) );
  oa21d1_hd U837 ( .A(n315), .B(n1), .C(n42), .Y(n198) );
  oa21d1_hd U838 ( .A(n316), .B(n1), .C(n43), .Y(n199) );
  oa21d1_hd U839 ( .A(n317), .B(n1), .C(n44), .Y(n200) );
  oa21d1_hd U840 ( .A(n318), .B(n1), .C(n45), .Y(n201) );
  oa21d1_hd U841 ( .A(n319), .B(n1), .C(n46), .Y(n202) );
  oa21d1_hd U842 ( .A(n320), .B(n1), .C(n47), .Y(n203) );
  oa21d1_hd U843 ( .A(n321), .B(n1), .C(n48), .Y(n204) );
  oa21d1_hd U844 ( .A(n322), .B(n1), .C(n215), .Y(n205) );
  oa21d1_hd U845 ( .A(n323), .B(n1), .C(n216), .Y(n206) );
  oa21d1_hd U846 ( .A(n324), .B(n1), .C(n217), .Y(n207) );
  oa21d1_hd U847 ( .A(n325), .B(n1), .C(n218), .Y(n208) );
  oa21d1_hd U848 ( .A(n331), .B(n1), .C(n219), .Y(n209) );
  oa21d1_hd U849 ( .A(n213), .B(n222), .C(n220), .Y(n224) );
  ao22d1_hd U850 ( .A(n223), .B(n225), .C(n224), .D(n598), .Y(n210) );
  ao22d1_hd U851 ( .A(n225), .B(n598), .C(n597), .D(n224), .Y(n211) );
  nr2d1_hd U852 ( .A(n804), .B(n594), .Y(n227) );
  ao211d1_hd U853 ( .A(n803), .B(n227), .C(n329), .D(n226), .Y(n212) );
  oa21d1_hd U854 ( .A(n2), .B(n228), .C(n801), .Y(n214) );
  ao22d1_hd U855 ( .A(n4), .B(o_Y_DATA[31]), .C(n3), .D(r_add_B[31]), .Y(n229)
         );
  oa21d1_hd U856 ( .A(r_x_data[63]), .B(n2), .C(n229), .Y(n348) );
  ao22d1_hd U857 ( .A(n332), .B(r_x_data[62]), .C(n3), .D(r_add_B[30]), .Y(
        n230) );
  oa21d1_hd U858 ( .A(n689), .B(n262), .C(n230), .Y(n349) );
  ao22d1_hd U859 ( .A(n332), .B(r_x_data[61]), .C(n3), .D(r_add_B[29]), .Y(
        n231) );
  oa21d1_hd U860 ( .A(n689), .B(n263), .C(n231), .Y(n350) );
  ao22d1_hd U861 ( .A(n332), .B(r_x_data[60]), .C(n3), .D(r_add_B[28]), .Y(
        n232) );
  oa21d1_hd U862 ( .A(n689), .B(n264), .C(n232), .Y(n351) );
  ao22d1_hd U863 ( .A(n332), .B(r_x_data[59]), .C(n3), .D(r_add_B[27]), .Y(
        n233) );
  oa21d1_hd U864 ( .A(n689), .B(n265), .C(n233), .Y(n352) );
  ao22d1_hd U865 ( .A(n332), .B(r_x_data[58]), .C(n3), .D(r_add_B[26]), .Y(
        n234) );
  oa21d1_hd U866 ( .A(n689), .B(n266), .C(n234), .Y(n353) );
  ao22d1_hd U867 ( .A(n332), .B(r_x_data[57]), .C(n3), .D(r_add_B[25]), .Y(
        n235) );
  oa21d1_hd U868 ( .A(n689), .B(n267), .C(n235), .Y(n354) );
  ao22d1_hd U869 ( .A(n332), .B(r_x_data[56]), .C(n3), .D(r_add_B[24]), .Y(
        n236) );
  oa21d1_hd U870 ( .A(n689), .B(n268), .C(n236), .Y(n355) );
  ao22d1_hd U871 ( .A(n332), .B(r_x_data[55]), .C(n3), .D(r_add_B[23]), .Y(
        n237) );
  oa21d1_hd U872 ( .A(n689), .B(n269), .C(n237), .Y(n356) );
  ao22d1_hd U873 ( .A(n332), .B(r_x_data[54]), .C(n3), .D(r_add_B[22]), .Y(
        n238) );
  oa21d1_hd U874 ( .A(n689), .B(n270), .C(n238), .Y(n357) );
  ao22d1_hd U875 ( .A(n332), .B(r_x_data[53]), .C(n3), .D(r_add_B[21]), .Y(
        n239) );
  oa21d1_hd U876 ( .A(n689), .B(n271), .C(n239), .Y(n358) );
  ao22d1_hd U877 ( .A(n332), .B(r_x_data[52]), .C(n3), .D(r_add_B[20]), .Y(
        n240) );
  oa21d1_hd U878 ( .A(n689), .B(n272), .C(n240), .Y(n359) );
  ao22d1_hd U879 ( .A(n332), .B(r_x_data[51]), .C(n3), .D(r_add_B[19]), .Y(
        n241) );
  oa21d1_hd U880 ( .A(n689), .B(n273), .C(n241), .Y(n360) );
  ao22d1_hd U881 ( .A(n332), .B(r_x_data[50]), .C(n3), .D(r_add_B[18]), .Y(
        n242) );
  oa21d1_hd U882 ( .A(n689), .B(n274), .C(n242), .Y(n361) );
  ao22d1_hd U884 ( .A(n332), .B(r_x_data[49]), .C(n3), .D(r_add_B[17]), .Y(
        n243) );
  oa21d1_hd U885 ( .A(n689), .B(n275), .C(n243), .Y(n362) );
  ao22d1_hd U886 ( .A(n332), .B(r_x_data[48]), .C(n3), .D(r_add_B[16]), .Y(
        n244) );
  oa21d1_hd U887 ( .A(n689), .B(n276), .C(n244), .Y(n363) );
  ao22d1_hd U888 ( .A(n332), .B(r_x_data[47]), .C(n3), .D(r_add_B[15]), .Y(
        n245) );
  oa21d1_hd U889 ( .A(n689), .B(n277), .C(n245), .Y(n364) );
  ao22d1_hd U890 ( .A(n332), .B(r_x_data[46]), .C(n3), .D(r_add_B[14]), .Y(
        n246) );
  oa21d1_hd U891 ( .A(n689), .B(n278), .C(n246), .Y(n365) );
  ao22d1_hd U892 ( .A(n332), .B(r_x_data[45]), .C(n3), .D(r_add_B[13]), .Y(
        n247) );
  oa21d1_hd U893 ( .A(n689), .B(n279), .C(n247), .Y(n366) );
  ao22d1_hd U894 ( .A(n332), .B(r_x_data[44]), .C(n3), .D(r_add_B[12]), .Y(
        n248) );
  oa21d1_hd U895 ( .A(n689), .B(n280), .C(n248), .Y(n367) );
  ao22d1_hd U896 ( .A(n332), .B(r_x_data[43]), .C(n3), .D(r_add_B[11]), .Y(
        n249) );
  oa21d1_hd U897 ( .A(n689), .B(n281), .C(n249), .Y(n368) );
  ao22d1_hd U898 ( .A(n332), .B(r_x_data[42]), .C(n3), .D(r_add_B[10]), .Y(
        n250) );
  oa21d1_hd U899 ( .A(n689), .B(n282), .C(n250), .Y(n369) );
  ao22d1_hd U900 ( .A(n332), .B(r_x_data[41]), .C(n3), .D(r_add_B[9]), .Y(n251) );
  oa21d1_hd U901 ( .A(n689), .B(n283), .C(n251), .Y(n370) );
  ao22d1_hd U902 ( .A(n332), .B(r_x_data[40]), .C(n3), .D(r_add_B[8]), .Y(n252) );
  oa21d1_hd U903 ( .A(n689), .B(n284), .C(n252), .Y(n371) );
  ao22d1_hd U904 ( .A(n332), .B(r_x_data[39]), .C(n3), .D(r_add_B[7]), .Y(n253) );
  oa21d1_hd U905 ( .A(n689), .B(n285), .C(n253), .Y(n372) );
  ao22d1_hd U906 ( .A(n332), .B(r_x_data[38]), .C(n3), .D(r_add_B[6]), .Y(n254) );
  oa21d1_hd U907 ( .A(n689), .B(n286), .C(n254), .Y(n373) );
  ao22d1_hd U908 ( .A(n332), .B(r_x_data[37]), .C(n3), .D(r_add_B[5]), .Y(n255) );
  oa21d1_hd U909 ( .A(n689), .B(n287), .C(n255), .Y(n374) );
  ao22d1_hd U910 ( .A(n332), .B(r_x_data[36]), .C(n3), .D(r_add_B[4]), .Y(n256) );
  oa21d1_hd U911 ( .A(n689), .B(n288), .C(n256), .Y(n375) );
  ao22d1_hd U912 ( .A(n332), .B(r_x_data[35]), .C(n3), .D(r_add_B[3]), .Y(n257) );
  oa21d1_hd U913 ( .A(n689), .B(n289), .C(n257), .Y(n376) );
  ao22d1_hd U914 ( .A(n332), .B(r_x_data[34]), .C(n3), .D(r_add_B[2]), .Y(n258) );
  oa21d1_hd U915 ( .A(n689), .B(n290), .C(n258), .Y(n377) );
  ao22d1_hd U916 ( .A(n332), .B(r_x_data[33]), .C(n3), .D(r_add_B[1]), .Y(n259) );
  oa21d1_hd U918 ( .A(n689), .B(n291), .C(n259), .Y(n378) );
  ao22d1_hd U920 ( .A(n332), .B(r_x_data[32]), .C(n3), .D(r_add_B[0]), .Y(n260) );
  oa21d1_hd U922 ( .A(n689), .B(n293), .C(n260), .Y(n379) );
  oa21d1_hd U924 ( .A(n261), .B(n292), .C(n766), .Y(n380) );
  oa21d1_hd U926 ( .A(n262), .B(n292), .C(n765), .Y(n381) );
  oa21d1_hd U928 ( .A(n263), .B(n292), .C(n764), .Y(n382) );
  oa21d1_hd U930 ( .A(n264), .B(n292), .C(n763), .Y(n383) );
  oa21d1_hd U932 ( .A(n265), .B(n292), .C(n762), .Y(n384) );
  oa21d1_hd U934 ( .A(n266), .B(n292), .C(n761), .Y(n385) );
  oa21d1_hd U936 ( .A(n267), .B(n292), .C(n760), .Y(n386) );
  oa21d1_hd U938 ( .A(n268), .B(n292), .C(n759), .Y(n387) );
  oa21d1_hd U940 ( .A(n269), .B(n292), .C(n758), .Y(n388) );
  oa21d1_hd U941 ( .A(n270), .B(n292), .C(n757), .Y(n389) );
  oa21d1_hd U943 ( .A(n271), .B(n292), .C(n756), .Y(n390) );
  oa21d1_hd U944 ( .A(n272), .B(n292), .C(n755), .Y(n391) );
  oa21d1_hd U946 ( .A(n273), .B(n292), .C(n754), .Y(n392) );
  oa21d1_hd U947 ( .A(n274), .B(n292), .C(n753), .Y(n393) );
  oa21d1_hd U948 ( .A(n275), .B(n292), .C(n752), .Y(n394) );
  oa21d1_hd U950 ( .A(n276), .B(n292), .C(n751), .Y(n395) );
  oa21d1_hd U951 ( .A(n277), .B(n292), .C(n750), .Y(n396) );
  oa21d1_hd U952 ( .A(n278), .B(n292), .C(n749), .Y(n397) );
  oa21d1_hd U953 ( .A(n279), .B(n292), .C(n748), .Y(n398) );
  oa21d1_hd U957 ( .A(n280), .B(n292), .C(n747), .Y(n399) );
  oa21d1_hd U958 ( .A(n281), .B(n292), .C(n746), .Y(n400) );
  oa21d1_hd U959 ( .A(n282), .B(n292), .C(n745), .Y(n401) );
  oa21d1_hd U960 ( .A(n283), .B(n292), .C(n744), .Y(n402) );
  oa21d1_hd U961 ( .A(n284), .B(n292), .C(n743), .Y(n403) );
  oa21d1_hd U962 ( .A(n285), .B(n292), .C(n742), .Y(n404) );
  oa21d1_hd U963 ( .A(n286), .B(n292), .C(n741), .Y(n405) );
  oa21d1_hd U964 ( .A(n287), .B(n292), .C(n740), .Y(n406) );
  oa21d1_hd U965 ( .A(n288), .B(n292), .C(n739), .Y(n407) );
  oa21d1_hd U966 ( .A(n289), .B(n292), .C(n738), .Y(n408) );
  oa21d1_hd U967 ( .A(n290), .B(n292), .C(n737), .Y(n409) );
  oa21d1_hd U968 ( .A(n291), .B(n292), .C(n736), .Y(n410) );
  oa21d1_hd U969 ( .A(n293), .B(n292), .C(n733), .Y(n411) );
  oa22d1_hd U970 ( .A(n695), .B(n295), .C(n731), .D(n598), .Y(n412) );
  oa21d1_hd U971 ( .A(n2), .B(n296), .C(n728), .Y(n413) );
  oa21d1_hd U972 ( .A(n2), .B(n297), .C(n727), .Y(n414) );
  oa21d1_hd U973 ( .A(n2), .B(n298), .C(n726), .Y(n415) );
  oa21d1_hd U974 ( .A(n2), .B(n299), .C(n725), .Y(n416) );
  oa21d1_hd U975 ( .A(n2), .B(n300), .C(n724), .Y(n417) );
  oa21d1_hd U976 ( .A(n2), .B(n301), .C(n723), .Y(n418) );
  oa21d1_hd U977 ( .A(n2), .B(n302), .C(n722), .Y(n419) );
  oa21d1_hd U978 ( .A(n2), .B(n303), .C(n721), .Y(n420) );
  oa21d1_hd U979 ( .A(n2), .B(n304), .C(n720), .Y(n421) );
  oa21d1_hd U980 ( .A(n2), .B(n305), .C(n719), .Y(n422) );
  oa21d1_hd U981 ( .A(n2), .B(n306), .C(n718), .Y(n423) );
  oa21d1_hd U982 ( .A(n2), .B(n307), .C(n717), .Y(n424) );
  oa21d1_hd U983 ( .A(n2), .B(n308), .C(n716), .Y(n425) );
  oa21d1_hd U984 ( .A(n2), .B(n309), .C(n715), .Y(n426) );
  oa21d1_hd U985 ( .A(n2), .B(n310), .C(n714), .Y(n427) );
  oa21d1_hd U986 ( .A(n2), .B(n311), .C(n713), .Y(n428) );
  oa21d1_hd U987 ( .A(n2), .B(n312), .C(n712), .Y(n429) );
  oa21d1_hd U988 ( .A(n2), .B(n313), .C(n711), .Y(n430) );
  oa21d1_hd U989 ( .A(n2), .B(n314), .C(n710), .Y(n431) );
  oa21d1_hd U990 ( .A(n2), .B(n315), .C(n709), .Y(n432) );
  oa21d1_hd U991 ( .A(n2), .B(n316), .C(n708), .Y(n433) );
  oa21d1_hd U992 ( .A(n2), .B(n317), .C(n707), .Y(n434) );
  oa21d1_hd U993 ( .A(n2), .B(n318), .C(n706), .Y(n435) );
  oa21d1_hd U994 ( .A(n2), .B(n319), .C(n705), .Y(n436) );
  oa21d1_hd U995 ( .A(n2), .B(n320), .C(n704), .Y(n437) );
  oa21d1_hd U996 ( .A(n2), .B(n321), .C(n703), .Y(n438) );
  oa21d1_hd U997 ( .A(n2), .B(n322), .C(n702), .Y(n439) );
  oa21d1_hd U998 ( .A(n2), .B(n323), .C(n701), .Y(n440) );
  oa21d1_hd U999 ( .A(n2), .B(n324), .C(n700), .Y(n441) );
  oa21d1_hd U1000 ( .A(n2), .B(n325), .C(n699), .Y(n442) );
  nd3d1_hd U1001 ( .A(n698), .B(w_add_Z_STB), .C(n597), .Y(n326) );
  scg17d1_hd U1002 ( .A(n327), .B(r_add_Z_ACK), .C(n6), .D(n326), .Y(n443) );
  oa21d1_hd U1003 ( .A(n694), .B(n695), .C(o_Y_DATA_VALID), .Y(n328) );
  nd2bd1_hd U1004 ( .AN(n329), .B(n328), .Y(n444) );
  oa21d1_hd U1005 ( .A(n2), .B(n330), .C(n691), .Y(n447) );
  oa21d1_hd U1006 ( .A(n2), .B(n331), .C(n688), .Y(n448) );
  oa21d1_hd U1007 ( .A(n2), .B(n333), .C(n686), .Y(n81) );
  oa21d1_hd U1008 ( .A(n2), .B(n334), .C(n685), .Y(n82) );
  oa21d1_hd U1009 ( .A(n2), .B(n335), .C(n684), .Y(n83) );
  oa21d1_hd U1010 ( .A(n2), .B(n336), .C(n683), .Y(n84) );
  oa21d1_hd U1011 ( .A(n2), .B(n337), .C(n682), .Y(n85) );
  oa21d1_hd U1012 ( .A(n2), .B(n338), .C(n681), .Y(n86) );
  oa21d1_hd U1013 ( .A(n2), .B(n339), .C(n680), .Y(n87) );
  oa21d1_hd U1014 ( .A(n2), .B(n340), .C(n679), .Y(n88) );
  oa21d1_hd U1015 ( .A(n2), .B(n341), .C(n678), .Y(n89) );
  oa21d1_hd U1016 ( .A(n2), .B(n342), .C(n677), .Y(n90) );
  oa21d1_hd U1017 ( .A(n2), .B(n343), .C(n676), .Y(n91) );
  oa21d1_hd U1018 ( .A(n2), .B(n344), .C(n675), .Y(n92) );
  oa21d1_hd U1019 ( .A(n2), .B(n345), .C(n674), .Y(n93) );
  oa21d1_hd U1020 ( .A(n2), .B(n346), .C(n673), .Y(n94) );
  oa21d1_hd U1021 ( .A(n2), .B(n347), .C(n672), .Y(n95) );
  oa21d1_hd U1022 ( .A(n2), .B(n445), .C(n671), .Y(n96) );
  oa21d1_hd U1023 ( .A(n2), .B(n446), .C(n670), .Y(n97) );
  oa21d1_hd U1024 ( .A(n2), .B(n449), .C(n669), .Y(n98) );
  oa21d1_hd U1025 ( .A(n2), .B(n451), .C(n666), .Y(n99) );
endmodule


module converter_f2i ( i_A, i_A_STB, o_A_ACK, o_Z, o_Z_STB, i_Z_ACK, i_CLK, 
        i_RST );
  input [31:0] i_A;
  output [31:0] o_Z;
  input i_A_STB, i_Z_ACK, i_CLK, i_RST;
  output o_A_ACK, o_Z_STB;
  wire   a_s, N65, N174, N175, N176, N177, N178, N179, N180, N181, N182, n1,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n427, n473, n475, n731, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n165, n166, n167, n168, n169, n170, n171,
         n172, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263;
  wire   [2:0] state;
  wire   [31:0] a;
  wire   [8:0] a_e;
  wire   [31:1] a_m;
  wire   [31:8] z;

  fd1qd1_hd z_reg_30_ ( .D(n142), .CK(i_CLK), .Q(z[30]) );
  fd1qd1_hd z_reg_29_ ( .D(n143), .CK(i_CLK), .Q(z[29]) );
  fd1qd1_hd z_reg_28_ ( .D(n144), .CK(i_CLK), .Q(z[28]) );
  fd1qd1_hd z_reg_27_ ( .D(n145), .CK(i_CLK), .Q(z[27]) );
  fd1qd1_hd z_reg_26_ ( .D(n146), .CK(i_CLK), .Q(z[26]) );
  fd1qd1_hd z_reg_25_ ( .D(n147), .CK(i_CLK), .Q(z[25]) );
  fd1qd1_hd z_reg_24_ ( .D(n148), .CK(i_CLK), .Q(z[24]) );
  fd1qd1_hd z_reg_23_ ( .D(n149), .CK(i_CLK), .Q(z[23]) );
  fd1qd1_hd z_reg_22_ ( .D(n150), .CK(i_CLK), .Q(z[22]) );
  fd1qd1_hd z_reg_21_ ( .D(n151), .CK(i_CLK), .Q(z[21]) );
  fd1qd1_hd z_reg_20_ ( .D(n152), .CK(i_CLK), .Q(z[20]) );
  fd1qd1_hd z_reg_19_ ( .D(n153), .CK(i_CLK), .Q(z[19]) );
  fd1qd1_hd z_reg_18_ ( .D(n154), .CK(i_CLK), .Q(z[18]) );
  fd1qd1_hd z_reg_17_ ( .D(n155), .CK(i_CLK), .Q(z[17]) );
  fd1qd1_hd z_reg_16_ ( .D(n156), .CK(i_CLK), .Q(z[16]) );
  fd1qd1_hd z_reg_15_ ( .D(n157), .CK(i_CLK), .Q(z[15]) );
  fd1qd1_hd z_reg_14_ ( .D(n158), .CK(i_CLK), .Q(z[14]) );
  fd1qd1_hd z_reg_13_ ( .D(n159), .CK(i_CLK), .Q(z[13]) );
  fd1qd1_hd z_reg_12_ ( .D(n160), .CK(i_CLK), .Q(z[12]) );
  fd1qd1_hd z_reg_11_ ( .D(n161), .CK(i_CLK), .Q(z[11]) );
  fd1qd1_hd z_reg_10_ ( .D(n162), .CK(i_CLK), .Q(z[10]) );
  fd1qd1_hd z_reg_9_ ( .D(n163), .CK(i_CLK), .Q(z[9]) );
  fd1qd1_hd z_reg_8_ ( .D(n164), .CK(i_CLK), .Q(z[8]) );
  fd1qd1_hd z_reg_31_ ( .D(n141), .CK(i_CLK), .Q(z[31]) );
  fd1qd1_hd o_A_ACK_reg ( .D(n208), .CK(i_CLK), .Q(o_A_ACK) );
  fd1qd1_hd a_m_reg_31_ ( .D(n204), .CK(i_CLK), .Q(a_m[31]) );
  fd1qd1_hd a_m_reg_30_ ( .D(n173), .CK(i_CLK), .Q(a_m[30]) );
  fd1eqd1_hd a_e_reg_3_ ( .D(N177), .E(n475), .CK(i_CLK), .Q(a_e[3]) );
  fd1eqd1_hd a_e_reg_8_ ( .D(N182), .E(n475), .CK(i_CLK), .Q(a_e[8]) );
  fd1qd1_hd state_reg_0_ ( .D(n206), .CK(i_CLK), .Q(state[0]) );
  fd1qd1_hd state_reg_2_ ( .D(n207), .CK(i_CLK), .Q(state[2]) );
  fd1qd1_hd state_reg_1_ ( .D(n205), .CK(i_CLK), .Q(state[1]) );
  fd1eqd1_hd a_e_reg_6_ ( .D(N180), .E(n475), .CK(i_CLK), .Q(a_e[6]) );
  fd1qd1_hd a_m_reg_28_ ( .D(n175), .CK(i_CLK), .Q(a_m[28]) );
  fd1qd1_hd a_m_reg_26_ ( .D(n177), .CK(i_CLK), .Q(a_m[26]) );
  fd1eqd1_hd a_e_reg_0_ ( .D(N174), .E(n475), .CK(i_CLK), .Q(a_e[0]) );
  fd1eqd1_hd a_e_reg_4_ ( .D(N178), .E(n475), .CK(i_CLK), .Q(a_e[4]) );
  fd1eqd1_hd a_e_reg_2_ ( .D(N176), .E(n475), .CK(i_CLK), .Q(a_e[2]) );
  fd1eqd1_hd a_e_reg_1_ ( .D(N175), .E(n475), .CK(i_CLK), .Q(a_e[1]) );
  fd1qd1_hd a_m_reg_29_ ( .D(n174), .CK(i_CLK), .Q(a_m[29]) );
  fd1qd1_hd a_m_reg_27_ ( .D(n176), .CK(i_CLK), .Q(a_m[27]) );
  fd1eqd1_hd a_e_reg_5_ ( .D(N179), .E(n475), .CK(i_CLK), .Q(a_e[5]) );
  fd1eqd1_hd a_e_reg_7_ ( .D(N181), .E(n475), .CK(i_CLK), .Q(a_e[7]) );
  fd1qd1_hd a_m_reg_24_ ( .D(n179), .CK(i_CLK), .Q(a_m[24]) );
  fd1qd1_hd a_m_reg_22_ ( .D(n181), .CK(i_CLK), .Q(a_m[22]) );
  fd1qd1_hd a_m_reg_20_ ( .D(n183), .CK(i_CLK), .Q(a_m[20]) );
  fd1qd1_hd a_m_reg_25_ ( .D(n178), .CK(i_CLK), .Q(a_m[25]) );
  fd1qd1_hd a_m_reg_23_ ( .D(n180), .CK(i_CLK), .Q(a_m[23]) );
  fd1qd1_hd a_m_reg_21_ ( .D(n182), .CK(i_CLK), .Q(a_m[21]) );
  fd1qd1_hd a_m_reg_18_ ( .D(n185), .CK(i_CLK), .Q(a_m[18]) );
  fd1qd1_hd a_m_reg_16_ ( .D(n187), .CK(i_CLK), .Q(a_m[16]) );
  fd1qd1_hd a_m_reg_19_ ( .D(n184), .CK(i_CLK), .Q(a_m[19]) );
  fd1qd1_hd a_m_reg_17_ ( .D(n186), .CK(i_CLK), .Q(a_m[17]) );
  fd1qd1_hd a_m_reg_14_ ( .D(n189), .CK(i_CLK), .Q(a_m[14]) );
  fd1qd1_hd a_m_reg_12_ ( .D(n191), .CK(i_CLK), .Q(a_m[12]) );
  fd1qd1_hd a_m_reg_10_ ( .D(n193), .CK(i_CLK), .Q(a_m[10]) );
  fd1qd1_hd a_m_reg_15_ ( .D(n188), .CK(i_CLK), .Q(a_m[15]) );
  fd1qd1_hd a_m_reg_13_ ( .D(n190), .CK(i_CLK), .Q(a_m[13]) );
  fd1qd1_hd a_m_reg_11_ ( .D(n192), .CK(i_CLK), .Q(a_m[11]) );
  fd1qd1_hd a_m_reg_6_ ( .D(n197), .CK(i_CLK), .Q(a_m[6]) );
  fd1qd1_hd a_m_reg_8_ ( .D(n195), .CK(i_CLK), .Q(a_m[8]) );
  fd1qd1_hd a_m_reg_7_ ( .D(n196), .CK(i_CLK), .Q(a_m[7]) );
  fd1qd1_hd a_m_reg_9_ ( .D(n194), .CK(i_CLK), .Q(a_m[9]) );
  fd1qd1_hd a_m_reg_4_ ( .D(n199), .CK(i_CLK), .Q(a_m[4]) );
  fd1qd1_hd a_m_reg_2_ ( .D(n201), .CK(i_CLK), .Q(a_m[2]) );
  fd1qd1_hd a_m_reg_1_ ( .D(n202), .CK(i_CLK), .Q(a_m[1]) );
  fd1qd1_hd a_m_reg_5_ ( .D(n198), .CK(i_CLK), .Q(a_m[5]) );
  fd1qd1_hd a_m_reg_3_ ( .D(n200), .CK(i_CLK), .Q(a_m[3]) );
  fd1qd1_hd a_m_reg_0_ ( .D(n203), .CK(i_CLK), .Q(N65) );
  fd1eqd1_hd o_Z_reg_23_ ( .D(z[23]), .E(n1), .CK(i_CLK), .Q(o_Z[23]) );
  fd1eqd1_hd o_Z_reg_22_ ( .D(z[22]), .E(n1), .CK(i_CLK), .Q(o_Z[22]) );
  fd1eqd1_hd o_Z_reg_21_ ( .D(z[21]), .E(n1), .CK(i_CLK), .Q(o_Z[21]) );
  fd1eqd1_hd o_Z_reg_20_ ( .D(z[20]), .E(n1), .CK(i_CLK), .Q(o_Z[20]) );
  fd1eqd1_hd o_Z_reg_19_ ( .D(z[19]), .E(n1), .CK(i_CLK), .Q(o_Z[19]) );
  fd1eqd1_hd o_Z_reg_18_ ( .D(z[18]), .E(n1), .CK(i_CLK), .Q(o_Z[18]) );
  fd1eqd1_hd a_reg_31_ ( .D(i_A[31]), .E(n4), .CK(i_CLK), .Q(a[31]) );
  fd1eqd1_hd a_reg_30_ ( .D(i_A[30]), .E(n4), .CK(i_CLK), .Q(a[30]) );
  fd1eqd1_hd a_reg_29_ ( .D(i_A[29]), .E(n4), .CK(i_CLK), .Q(a[29]) );
  fd1eqd1_hd a_reg_28_ ( .D(i_A[28]), .E(n4), .CK(i_CLK), .Q(a[28]) );
  fd1eqd1_hd a_reg_27_ ( .D(i_A[27]), .E(n4), .CK(i_CLK), .Q(a[27]) );
  fd1eqd1_hd a_reg_26_ ( .D(i_A[26]), .E(n4), .CK(i_CLK), .Q(a[26]) );
  fd1eqd1_hd a_reg_25_ ( .D(i_A[25]), .E(n473), .CK(i_CLK), .Q(a[25]) );
  fd1eqd1_hd a_reg_24_ ( .D(i_A[24]), .E(n473), .CK(i_CLK), .Q(a[24]) );
  fd1eqd1_hd a_reg_23_ ( .D(i_A[23]), .E(n4), .CK(i_CLK), .Q(a[23]) );
  fd1eqd1_hd a_reg_22_ ( .D(i_A[22]), .E(n4), .CK(i_CLK), .Q(a[22]) );
  fd1eqd1_hd a_reg_21_ ( .D(i_A[21]), .E(n4), .CK(i_CLK), .Q(a[21]) );
  fd1eqd1_hd a_reg_20_ ( .D(i_A[20]), .E(n4), .CK(i_CLK), .Q(a[20]) );
  fd1eqd1_hd a_reg_19_ ( .D(i_A[19]), .E(n4), .CK(i_CLK), .Q(a[19]) );
  fd1eqd1_hd a_reg_5_ ( .D(i_A[5]), .E(n4), .CK(i_CLK), .Q(a[5]) );
  fd1eqd1_hd a_reg_4_ ( .D(i_A[4]), .E(n4), .CK(i_CLK), .Q(a[4]) );
  fd1eqd1_hd a_reg_3_ ( .D(i_A[3]), .E(n4), .CK(i_CLK), .Q(a[3]) );
  fd1eqd1_hd a_reg_2_ ( .D(i_A[2]), .E(n4), .CK(i_CLK), .Q(a[2]) );
  fd1eqd1_hd a_reg_18_ ( .D(i_A[18]), .E(n4), .CK(i_CLK), .Q(a[18]) );
  fd1eqd1_hd a_reg_17_ ( .D(i_A[17]), .E(n4), .CK(i_CLK), .Q(a[17]) );
  fd1eqd1_hd a_reg_16_ ( .D(i_A[16]), .E(n4), .CK(i_CLK), .Q(a[16]) );
  fd1eqd1_hd a_reg_15_ ( .D(i_A[15]), .E(n4), .CK(i_CLK), .Q(a[15]) );
  fd1eqd1_hd a_reg_14_ ( .D(i_A[14]), .E(n4), .CK(i_CLK), .Q(a[14]) );
  fd1eqd1_hd a_reg_13_ ( .D(i_A[13]), .E(n4), .CK(i_CLK), .Q(a[13]) );
  fd1eqd1_hd a_reg_12_ ( .D(i_A[12]), .E(n4), .CK(i_CLK), .Q(a[12]) );
  fd1eqd1_hd a_reg_11_ ( .D(i_A[11]), .E(n4), .CK(i_CLK), .Q(a[11]) );
  fd1eqd1_hd a_reg_10_ ( .D(i_A[10]), .E(n4), .CK(i_CLK), .Q(a[10]) );
  fd1eqd1_hd a_reg_9_ ( .D(i_A[9]), .E(n4), .CK(i_CLK), .Q(a[9]) );
  fd1eqd1_hd a_reg_8_ ( .D(i_A[8]), .E(n473), .CK(i_CLK), .Q(a[8]) );
  fd1eqd1_hd a_reg_7_ ( .D(i_A[7]), .E(n473), .CK(i_CLK), .Q(a[7]) );
  fd1eqd1_hd a_reg_6_ ( .D(i_A[6]), .E(n473), .CK(i_CLK), .Q(a[6]) );
  fd1eqd1_hd a_reg_1_ ( .D(i_A[1]), .E(n473), .CK(i_CLK), .Q(a[1]) );
  fd1eqd1_hd a_reg_0_ ( .D(i_A[0]), .E(n473), .CK(i_CLK), .Q(a[0]) );
  fd1eqd1_hd o_Z_reg_31_ ( .D(z[31]), .E(n1), .CK(i_CLK), .Q(o_Z[31]) );
  fd1eqd1_hd o_Z_reg_30_ ( .D(z[30]), .E(n1), .CK(i_CLK), .Q(o_Z[30]) );
  fd1eqd1_hd o_Z_reg_29_ ( .D(z[29]), .E(n1), .CK(i_CLK), .Q(o_Z[29]) );
  fd1eqd1_hd o_Z_reg_28_ ( .D(z[28]), .E(n1), .CK(i_CLK), .Q(o_Z[28]) );
  fd1eqd1_hd o_Z_reg_27_ ( .D(z[27]), .E(n1), .CK(i_CLK), .Q(o_Z[27]) );
  fd1eqd1_hd o_Z_reg_26_ ( .D(z[26]), .E(n1), .CK(i_CLK), .Q(o_Z[26]) );
  fd1eqd1_hd o_Z_reg_25_ ( .D(z[25]), .E(n1), .CK(i_CLK), .Q(o_Z[25]) );
  fd1eqd1_hd o_Z_reg_24_ ( .D(z[24]), .E(n1), .CK(i_CLK), .Q(o_Z[24]) );
  fd1eqd1_hd o_Z_reg_17_ ( .D(z[17]), .E(n1), .CK(i_CLK), .Q(o_Z[17]) );
  fd1eqd1_hd o_Z_reg_16_ ( .D(z[16]), .E(n1), .CK(i_CLK), .Q(o_Z[16]) );
  fd1eqd1_hd o_Z_reg_15_ ( .D(z[15]), .E(n1), .CK(i_CLK), .Q(o_Z[15]) );
  fd1eqd1_hd o_Z_reg_14_ ( .D(z[14]), .E(n1), .CK(i_CLK), .Q(o_Z[14]) );
  fd1eqd1_hd o_Z_reg_13_ ( .D(z[13]), .E(n1), .CK(i_CLK), .Q(o_Z[13]) );
  fd1eqd1_hd o_Z_reg_12_ ( .D(z[12]), .E(n1), .CK(i_CLK), .Q(o_Z[12]) );
  fd1eqd1_hd o_Z_reg_11_ ( .D(z[11]), .E(n1), .CK(i_CLK), .Q(o_Z[11]) );
  fd1eqd1_hd o_Z_reg_10_ ( .D(z[10]), .E(n1), .CK(i_CLK), .Q(o_Z[10]) );
  fd1eqd1_hd o_Z_reg_9_ ( .D(z[9]), .E(n1), .CK(i_CLK), .Q(o_Z[9]) );
  fd1eqd1_hd o_Z_reg_8_ ( .D(z[8]), .E(n1), .CK(i_CLK), .Q(o_Z[8]) );
  ivd1_hd U406 ( .A(i_RST), .Y(n427) );
  fd1d1_hd o_Z_STB_reg ( .D(n263), .CK(i_CLK), .QN(o_Z_STB) );
  fd1eqd1_hd a_s_reg ( .D(a[31]), .E(n3), .CK(i_CLK), .Q(a_s) );
  clknd2d1_hd U223 ( .A(a_e[0]), .B(n5), .Y(n44) );
  clknd2d1_hd U224 ( .A(a_e[1]), .B(a_e[0]), .Y(n11) );
  clknd2d1_hd U225 ( .A(a[23]), .B(a[24]), .Y(n10) );
  clknd2d1_hd U226 ( .A(a_e[5]), .B(n25), .Y(n30) );
  clknd2d1_hd U227 ( .A(n26), .B(a[28]), .Y(n29) );
  clknd2d1_hd U228 ( .A(n246), .B(n262), .Y(n255) );
  clknd2d1_hd U229 ( .A(n427), .B(n255), .Y(n257) );
  clknd2d1_hd U230 ( .A(a_e[7]), .B(n35), .Y(n40) );
  clknd2d1_hd U231 ( .A(n49), .B(n48), .Y(n50) );
  clknd2d1_hd U232 ( .A(n256), .B(state[1]), .Y(n167) );
  clknd2d1_hd U233 ( .A(a_e[3]), .B(n15), .Y(n21) );
  clknd2d1_hd U234 ( .A(n16), .B(a[26]), .Y(n20) );
  clknd2d1_hd U235 ( .A(n244), .B(n256), .Y(n261) );
  clknd2d1_hd U236 ( .A(n47), .B(n46), .Y(n138) );
  clknd2d1_hd U237 ( .A(n133), .B(n240), .Y(n129) );
  clknd2d1_hd U238 ( .A(n125), .B(n236), .Y(n122) );
  clknd2d1_hd U239 ( .A(n118), .B(n233), .Y(n115) );
  clknd2d1_hd U240 ( .A(n111), .B(n230), .Y(n108) );
  clknd2d1_hd U241 ( .A(n104), .B(n227), .Y(n101) );
  clknd2d1_hd U242 ( .A(n97), .B(n224), .Y(n94) );
  clknd2d1_hd U243 ( .A(n90), .B(n221), .Y(n87) );
  clknd2d1_hd U244 ( .A(n83), .B(n218), .Y(n80) );
  clknd2d1_hd U245 ( .A(n76), .B(n215), .Y(n73) );
  clknd2d1_hd U246 ( .A(n69), .B(n212), .Y(n66) );
  clknd2d1_hd U247 ( .A(n62), .B(n209), .Y(n59) );
  clknd2d1_hd U248 ( .A(a[30]), .B(n34), .Y(n38) );
  clknd2d1_hd U249 ( .A(n8), .B(n7), .Y(N175) );
  clknd2d1_hd U250 ( .A(n253), .B(n6), .Y(n8) );
  clknd2d1_hd U251 ( .A(n14), .B(n13), .Y(N176) );
  clknd2d1_hd U252 ( .A(n24), .B(n23), .Y(N178) );
  clknd2d1_hd U253 ( .A(n29), .B(n28), .Y(n33) );
  clknd2d1_hd U254 ( .A(state[1]), .B(n250), .Y(n249) );
  clknd2d1_hd U255 ( .A(n252), .B(n251), .Y(n206) );
  clknd2d1_hd U256 ( .A(n42), .B(n41), .Y(N182) );
  clknd2d1_hd U257 ( .A(n51), .B(n40), .Y(n39) );
  clknd2d1_hd U258 ( .A(n18), .B(n17), .Y(N177) );
  clknd2d1_hd U259 ( .A(n2), .B(z[31]), .Y(n56) );
  clknd2d1_hd U260 ( .A(a_s), .B(n138), .Y(n139) );
  clknd2d1_hd U261 ( .A(a_m[9]), .B(n136), .Y(n134) );
  clknd2d1_hd U262 ( .A(a_s), .B(n129), .Y(n130) );
  clknd2d1_hd U263 ( .A(a_m[11]), .B(n127), .Y(n126) );
  clknd2d1_hd U264 ( .A(a_s), .B(n122), .Y(n123) );
  clknd2d1_hd U265 ( .A(a_m[13]), .B(n120), .Y(n119) );
  clknd2d1_hd U266 ( .A(a_s), .B(n115), .Y(n116) );
  clknd2d1_hd U267 ( .A(a_m[15]), .B(n113), .Y(n112) );
  clknd2d1_hd U268 ( .A(a_s), .B(n108), .Y(n109) );
  clknd2d1_hd U269 ( .A(a_m[17]), .B(n106), .Y(n105) );
  clknd2d1_hd U270 ( .A(a_s), .B(n101), .Y(n102) );
  clknd2d1_hd U271 ( .A(a_m[19]), .B(n99), .Y(n98) );
  clknd2d1_hd U272 ( .A(a_s), .B(n94), .Y(n95) );
  clknd2d1_hd U273 ( .A(a_m[21]), .B(n92), .Y(n91) );
  clknd2d1_hd U274 ( .A(a_s), .B(n87), .Y(n88) );
  clknd2d1_hd U275 ( .A(a_m[23]), .B(n85), .Y(n84) );
  clknd2d1_hd U276 ( .A(a_s), .B(n80), .Y(n81) );
  clknd2d1_hd U277 ( .A(a_m[25]), .B(n78), .Y(n77) );
  clknd2d1_hd U278 ( .A(a_s), .B(n73), .Y(n74) );
  clknd2d1_hd U279 ( .A(a_m[27]), .B(n71), .Y(n70) );
  clknd2d1_hd U280 ( .A(a_s), .B(n66), .Y(n67) );
  clknd2d1_hd U281 ( .A(a_m[29]), .B(n64), .Y(n63) );
  clknd2d1_hd U282 ( .A(a_s), .B(n59), .Y(n60) );
  xo2d1_hd U283 ( .A(a_m[14]), .B(n116), .Y(n117) );
  xo2d1_hd U284 ( .A(a_m[12]), .B(n123), .Y(n124) );
  xo2d1_hd U285 ( .A(a_m[10]), .B(n130), .Y(n131) );
  xo2d1_hd U286 ( .A(a_m[8]), .B(n139), .Y(n165) );
  scg2d1_hd U287 ( .A(a_m[5]), .B(n242), .C(a_m[4]), .D(n241), .Y(n199) );
  scg2d1_hd U288 ( .A(a_m[5]), .B(n241), .C(a_m[6]), .D(n242), .Y(n198) );
  scg2d1_hd U289 ( .A(a_m[7]), .B(n242), .C(a_m[6]), .D(n241), .Y(n197) );
  scg2d1_hd U290 ( .A(a_m[1]), .B(n242), .C(N65), .D(n241), .Y(n203) );
  scg2d1_hd U291 ( .A(a_m[8]), .B(n242), .C(a_m[7]), .D(n241), .Y(n196) );
  scg2d1_hd U292 ( .A(a_m[3]), .B(n241), .C(a_m[4]), .D(n242), .Y(n200) );
  scg2d1_hd U293 ( .A(a_m[3]), .B(n242), .C(a_m[2]), .D(n241), .Y(n201) );
  scg2d1_hd U294 ( .A(a_m[1]), .B(n241), .C(a_m[2]), .D(n242), .Y(n202) );
  xo2d1_hd U295 ( .A(a_m[30]), .B(n60), .Y(n61) );
  xo2d1_hd U296 ( .A(a_m[28]), .B(n67), .Y(n68) );
  xo2d1_hd U297 ( .A(a_m[26]), .B(n74), .Y(n75) );
  xo2d1_hd U298 ( .A(a_m[24]), .B(n81), .Y(n82) );
  xo2d1_hd U299 ( .A(a_m[22]), .B(n88), .Y(n89) );
  xo2d1_hd U300 ( .A(a_m[20]), .B(n95), .Y(n96) );
  xo2d1_hd U301 ( .A(a_m[18]), .B(n102), .Y(n103) );
  xo2d1_hd U302 ( .A(a_m[16]), .B(n109), .Y(n110) );
  scg10d1_hd U303 ( .A(n243), .B(n54), .C(n53), .D(n52), .Y(n58) );
  or2d1_hd U304 ( .A(state[0]), .B(n167), .Y(n731) );
  or4d1_hd U305 ( .A(a_e[4]), .B(a_e[3]), .C(a_e[2]), .D(n51), .Y(n43) );
  scg20d4_hd U306 ( .A(n169), .B(n168), .C(n167), .Y(n475) );
  nid2_hd U307 ( .A(n140), .Y(n2) );
  ivd1_hd U308 ( .A(n135), .Y(n166) );
  nd2d1_hd U309 ( .A(n253), .B(n475), .Y(n239) );
  nr2d1_hd U310 ( .A(a_m[30]), .B(n59), .Y(n55) );
  nid2_hd U311 ( .A(n473), .Y(n4) );
  ivd2_hd U312 ( .A(n475), .Y(n241) );
  ivd2_hd U313 ( .A(n239), .Y(n242) );
  nr2d1_hd U314 ( .A(n254), .B(n245), .Y(n140) );
  nr2d1_hd U315 ( .A(n168), .B(n54), .Y(n245) );
  ivd1_hd U316 ( .A(n253), .Y(n54) );
  nr2d1_hd U317 ( .A(n169), .B(n167), .Y(n253) );
  ao22d1_hd U318 ( .A(n55), .B(n243), .C(n51), .D(n50), .Y(n168) );
  nr2d1_hd U319 ( .A(a_m[28]), .B(n66), .Y(n62) );
  nr2d1_hd U320 ( .A(a_m[26]), .B(n73), .Y(n69) );
  ivd1_hd U321 ( .A(a_m[11]), .Y(n236) );
  ivd1_hd U322 ( .A(a_m[9]), .Y(n240) );
  scg12d1_hd U323 ( .A(o_A_ACK), .B(i_A_STB), .C(n261), .Y(n473) );
  ivd1_hd U324 ( .A(a_s), .Y(n132) );
  ivd2_hd U325 ( .A(n731), .Y(n3) );
  nr3d2_hd U326 ( .A(a_m[31]), .B(n140), .C(n54), .Y(n135) );
  ivd1_hd U327 ( .A(state[2]), .Y(n256) );
  nr2d1_hd U328 ( .A(n22), .B(n21), .Y(n25) );
  ivd1_hd U329 ( .A(a_m[31]), .Y(n243) );
  ivd1_hd U330 ( .A(a_m[29]), .Y(n209) );
  ivd1_hd U331 ( .A(a_m[27]), .Y(n212) );
  ivd1_hd U332 ( .A(a_m[25]), .Y(n215) );
  ivd1_hd U333 ( .A(a_m[23]), .Y(n218) );
  ivd1_hd U334 ( .A(a_m[21]), .Y(n221) );
  ivd1_hd U335 ( .A(a_m[19]), .Y(n224) );
  ivd1_hd U336 ( .A(a_m[17]), .Y(n227) );
  ivd1_hd U337 ( .A(n248), .Y(n53) );
  ivd1_hd U338 ( .A(state[0]), .Y(n169) );
  ivd1_hd U339 ( .A(a_e[8]), .Y(n51) );
  scg6d1_hd U340 ( .A(n36), .B(n33), .C(n32), .Y(N180) );
  ivd1_hd U341 ( .A(a[29]), .Y(n28) );
  scg14d1_hd U342 ( .A(n2), .B(z[15]), .C(n114), .Y(n157) );
  scg14d1_hd U343 ( .A(n2), .B(z[27]), .C(n72), .Y(n145) );
  scg14d1_hd U344 ( .A(n2), .B(z[17]), .C(n107), .Y(n155) );
  scg14d1_hd U345 ( .A(n2), .B(z[19]), .C(n100), .Y(n153) );
  scg14d1_hd U346 ( .A(n2), .B(z[9]), .C(n137), .Y(n163) );
  scg14d1_hd U347 ( .A(n2), .B(z[23]), .C(n86), .Y(n149) );
  scg14d1_hd U348 ( .A(n2), .B(z[13]), .C(n121), .Y(n159) );
  scg14d1_hd U349 ( .A(n2), .B(z[25]), .C(n79), .Y(n147) );
  scg14d1_hd U350 ( .A(n2), .B(z[29]), .C(n65), .Y(n143) );
  scg14d1_hd U351 ( .A(n2), .B(z[11]), .C(n128), .Y(n161) );
  scg14d1_hd U352 ( .A(n2), .B(z[21]), .C(n93), .Y(n151) );
  ivd1_hd U353 ( .A(a_e[4]), .Y(n22) );
  ivd1_hd U354 ( .A(a_m[15]), .Y(n230) );
  ivd1_hd U355 ( .A(a_m[13]), .Y(n233) );
  nr2d1_hd U356 ( .A(n247), .B(n53), .Y(n254) );
  nd2bd1_hd U357 ( .AN(a[30]), .B(n36), .Y(n41) );
  nr2d1_hd U358 ( .A(state[1]), .B(state[0]), .Y(n244) );
  nr3d1_hd U359 ( .A(n169), .B(state[2]), .C(state[1]), .Y(n248) );
  nr2d1_hd U360 ( .A(a_e[6]), .B(a_e[7]), .Y(n49) );
  ad2d2_hd U361 ( .A(n244), .B(state[2]), .Y(n1) );
  oa22d1_hd U362 ( .A(a_e[0]), .B(n54), .C(a[23]), .D(n731), .Y(N174) );
  ivd1_hd U363 ( .A(a_e[1]), .Y(n5) );
  oa21d1_hd U364 ( .A(n5), .B(a_e[0]), .C(n44), .Y(n6) );
  oa211d1_hd U365 ( .A(a[23]), .B(a[24]), .C(n3), .D(n10), .Y(n7) );
  ivd1_hd U366 ( .A(a[25]), .Y(n9) );
  nr2d1_hd U367 ( .A(n10), .B(n9), .Y(n16) );
  scg17d1_hd U368 ( .A(n10), .B(n9), .C(n16), .D(n3), .Y(n14) );
  ivd1_hd U369 ( .A(a_e[2]), .Y(n12) );
  nr2d1_hd U370 ( .A(n12), .B(n11), .Y(n15) );
  scg17d1_hd U371 ( .A(n12), .B(n11), .C(n15), .D(n253), .Y(n13) );
  oa211d1_hd U372 ( .A(a_e[3]), .B(n15), .C(n253), .D(n21), .Y(n18) );
  oa211d1_hd U373 ( .A(n16), .B(a[26]), .C(n3), .D(n20), .Y(n17) );
  ivd1_hd U374 ( .A(a[27]), .Y(n19) );
  nr2d1_hd U375 ( .A(n20), .B(n19), .Y(n26) );
  scg17d1_hd U376 ( .A(n20), .B(n19), .C(n26), .D(n3), .Y(n24) );
  scg17d1_hd U377 ( .A(n22), .B(n21), .C(n25), .D(n253), .Y(n23) );
  nr2d1_hd U378 ( .A(a_e[5]), .B(n25), .Y(n48) );
  oa211d1_hd U379 ( .A(n26), .B(a[28]), .C(n3), .D(n29), .Y(n27) );
  scg22d1_hd U380 ( .A(n253), .B(n30), .C(n48), .D(n27), .Y(N179) );
  nr2d1_hd U381 ( .A(n29), .B(n28), .Y(n34) );
  nr2d1_hd U382 ( .A(n34), .B(n731), .Y(n36) );
  ivd1_hd U383 ( .A(a_e[6]), .Y(n31) );
  nr2d1_hd U384 ( .A(n31), .B(n30), .Y(n35) );
  ao211d1_hd U385 ( .A(n31), .B(n30), .C(n35), .D(n54), .Y(n32) );
  oa211d1_hd U386 ( .A(a_e[7]), .B(n35), .C(n253), .D(n40), .Y(n37) );
  oa211d1_hd U387 ( .A(n731), .B(n38), .C(n37), .D(n41), .Y(N181) );
  oa211d1_hd U388 ( .A(n51), .B(n40), .C(n253), .D(n39), .Y(n42) );
  ivd1_hd U389 ( .A(n49), .Y(n45) );
  nr4d1_hd U390 ( .A(a_e[5]), .B(a_e[6]), .C(n44), .D(n43), .Y(n52) );
  oa22d1_hd U391 ( .A(a_e[5]), .B(n45), .C(n52), .D(n51), .Y(n247) );
  nr4d1_hd U392 ( .A(N65), .B(a_m[6]), .C(a_m[4]), .D(a_m[2]), .Y(n47) );
  nr4d1_hd U393 ( .A(a_m[7]), .B(a_m[1]), .C(a_m[5]), .D(a_m[3]), .Y(n46) );
  nr2d1_hd U394 ( .A(a_m[8]), .B(n138), .Y(n133) );
  nr2d1_hd U395 ( .A(a_m[10]), .B(n129), .Y(n125) );
  nr2d1_hd U396 ( .A(a_m[12]), .B(n122), .Y(n118) );
  nr2d1_hd U397 ( .A(a_m[14]), .B(n115), .Y(n111) );
  nr2d1_hd U398 ( .A(a_m[16]), .B(n108), .Y(n104) );
  nr2d1_hd U399 ( .A(a_m[18]), .B(n101), .Y(n97) );
  nr2d1_hd U400 ( .A(a_m[20]), .B(n94), .Y(n90) );
  nr2d1_hd U401 ( .A(a_m[22]), .B(n87), .Y(n83) );
  nr2d1_hd U402 ( .A(a_m[24]), .B(n80), .Y(n76) );
  scg13d1_hd U403 ( .A(n55), .B(n132), .C(n135), .Y(n57) );
  oa211d1_hd U404 ( .A(n2), .B(n58), .C(n57), .D(n56), .Y(n141) );
  oa22ad1_hd U405 ( .A(n166), .B(n61), .C(n2), .D(z[30]), .Y(n142) );
  nr2d1_hd U407 ( .A(n62), .B(n132), .Y(n64) );
  oa211d1_hd U408 ( .A(a_m[29]), .B(n64), .C(n135), .D(n63), .Y(n65) );
  oa22ad1_hd U409 ( .A(n166), .B(n68), .C(n2), .D(z[28]), .Y(n144) );
  nr2d1_hd U410 ( .A(n69), .B(n132), .Y(n71) );
  oa211d1_hd U411 ( .A(a_m[27]), .B(n71), .C(n135), .D(n70), .Y(n72) );
  oa22ad1_hd U412 ( .A(n166), .B(n75), .C(n2), .D(z[26]), .Y(n146) );
  nr2d1_hd U413 ( .A(n76), .B(n132), .Y(n78) );
  oa211d1_hd U414 ( .A(a_m[25]), .B(n78), .C(n135), .D(n77), .Y(n79) );
  oa22ad1_hd U415 ( .A(n166), .B(n82), .C(n2), .D(z[24]), .Y(n148) );
  nr2d1_hd U416 ( .A(n83), .B(n132), .Y(n85) );
  oa211d1_hd U417 ( .A(a_m[23]), .B(n85), .C(n135), .D(n84), .Y(n86) );
  oa22ad1_hd U418 ( .A(n166), .B(n89), .C(n2), .D(z[22]), .Y(n150) );
  nr2d1_hd U419 ( .A(n90), .B(n132), .Y(n92) );
  oa211d1_hd U420 ( .A(a_m[21]), .B(n92), .C(n135), .D(n91), .Y(n93) );
  oa22ad1_hd U421 ( .A(n166), .B(n96), .C(n2), .D(z[20]), .Y(n152) );
  nr2d1_hd U422 ( .A(n97), .B(n132), .Y(n99) );
  oa211d1_hd U423 ( .A(a_m[19]), .B(n99), .C(n135), .D(n98), .Y(n100) );
  oa22ad1_hd U424 ( .A(n166), .B(n103), .C(n2), .D(z[18]), .Y(n154) );
  nr2d1_hd U425 ( .A(n104), .B(n132), .Y(n106) );
  oa211d1_hd U426 ( .A(a_m[17]), .B(n106), .C(n135), .D(n105), .Y(n107) );
  oa22ad1_hd U427 ( .A(n166), .B(n110), .C(n2), .D(z[16]), .Y(n156) );
  nr2d1_hd U428 ( .A(n111), .B(n132), .Y(n113) );
  oa211d1_hd U429 ( .A(a_m[15]), .B(n113), .C(n135), .D(n112), .Y(n114) );
  oa22ad1_hd U430 ( .A(n166), .B(n117), .C(n2), .D(z[14]), .Y(n158) );
  nr2d1_hd U431 ( .A(n118), .B(n132), .Y(n120) );
  oa211d1_hd U432 ( .A(a_m[13]), .B(n120), .C(n135), .D(n119), .Y(n121) );
  oa22ad1_hd U433 ( .A(n166), .B(n124), .C(n2), .D(z[12]), .Y(n160) );
  nr2d1_hd U434 ( .A(n125), .B(n132), .Y(n127) );
  oa211d1_hd U435 ( .A(a_m[11]), .B(n127), .C(n135), .D(n126), .Y(n128) );
  oa22ad1_hd U436 ( .A(n166), .B(n131), .C(n2), .D(z[10]), .Y(n162) );
  nr2d1_hd U437 ( .A(n133), .B(n132), .Y(n136) );
  oa211d1_hd U438 ( .A(a_m[9]), .B(n136), .C(n135), .D(n134), .Y(n137) );
  oa22ad1_hd U439 ( .A(n166), .B(n165), .C(n2), .D(z[8]), .Y(n164) );
  ao22d1_hd U440 ( .A(a_m[30]), .B(n241), .C(n3), .D(a[22]), .Y(n170) );
  oa21d1_hd U441 ( .A(n243), .B(n239), .C(n170), .Y(n173) );
  ao22d1_hd U442 ( .A(a_m[30]), .B(n242), .C(n3), .D(a[21]), .Y(n171) );
  oa21d1_hd U443 ( .A(n475), .B(n209), .C(n171), .Y(n174) );
  ao22d1_hd U444 ( .A(a_m[28]), .B(n241), .C(n3), .D(a[20]), .Y(n172) );
  oa21d1_hd U445 ( .A(n209), .B(n239), .C(n172), .Y(n175) );
  ao22d1_hd U446 ( .A(a_m[28]), .B(n242), .C(n3), .D(a[19]), .Y(n210) );
  oa21d1_hd U447 ( .A(n475), .B(n212), .C(n210), .Y(n176) );
  ao22d1_hd U448 ( .A(a_m[26]), .B(n241), .C(n3), .D(a[18]), .Y(n211) );
  oa21d1_hd U449 ( .A(n212), .B(n239), .C(n211), .Y(n177) );
  ao22d1_hd U450 ( .A(a_m[26]), .B(n242), .C(n3), .D(a[17]), .Y(n213) );
  oa21d1_hd U451 ( .A(n475), .B(n215), .C(n213), .Y(n178) );
  ao22d1_hd U452 ( .A(a_m[24]), .B(n241), .C(n3), .D(a[16]), .Y(n214) );
  oa21d1_hd U453 ( .A(n215), .B(n239), .C(n214), .Y(n179) );
  ao22d1_hd U454 ( .A(a_m[24]), .B(n242), .C(n3), .D(a[15]), .Y(n216) );
  oa21d1_hd U455 ( .A(n475), .B(n218), .C(n216), .Y(n180) );
  ao22d1_hd U456 ( .A(a_m[22]), .B(n241), .C(n3), .D(a[14]), .Y(n217) );
  oa21d1_hd U457 ( .A(n218), .B(n239), .C(n217), .Y(n181) );
  ao22d1_hd U458 ( .A(a_m[22]), .B(n242), .C(n3), .D(a[13]), .Y(n219) );
  oa21d1_hd U459 ( .A(n475), .B(n221), .C(n219), .Y(n182) );
  ao22d1_hd U460 ( .A(a_m[20]), .B(n241), .C(n3), .D(a[12]), .Y(n220) );
  oa21d1_hd U461 ( .A(n221), .B(n239), .C(n220), .Y(n183) );
  ao22d1_hd U462 ( .A(a_m[20]), .B(n242), .C(n3), .D(a[11]), .Y(n222) );
  oa21d1_hd U463 ( .A(n475), .B(n224), .C(n222), .Y(n184) );
  ao22d1_hd U464 ( .A(a_m[18]), .B(n241), .C(n3), .D(a[10]), .Y(n223) );
  oa21d1_hd U465 ( .A(n224), .B(n239), .C(n223), .Y(n185) );
  ao22d1_hd U466 ( .A(a_m[18]), .B(n242), .C(n3), .D(a[9]), .Y(n225) );
  oa21d1_hd U467 ( .A(n475), .B(n227), .C(n225), .Y(n186) );
  ao22d1_hd U468 ( .A(a_m[16]), .B(n241), .C(n3), .D(a[8]), .Y(n226) );
  oa21d1_hd U469 ( .A(n227), .B(n239), .C(n226), .Y(n187) );
  ao22d1_hd U470 ( .A(a_m[16]), .B(n242), .C(n3), .D(a[7]), .Y(n228) );
  oa21d1_hd U471 ( .A(n475), .B(n230), .C(n228), .Y(n188) );
  ao22d1_hd U472 ( .A(a_m[14]), .B(n241), .C(n3), .D(a[6]), .Y(n229) );
  oa21d1_hd U473 ( .A(n230), .B(n239), .C(n229), .Y(n189) );
  ao22d1_hd U474 ( .A(a_m[14]), .B(n242), .C(n3), .D(a[5]), .Y(n231) );
  oa21d1_hd U475 ( .A(n475), .B(n233), .C(n231), .Y(n190) );
  ao22d1_hd U476 ( .A(a_m[12]), .B(n241), .C(n3), .D(a[4]), .Y(n232) );
  oa21d1_hd U477 ( .A(n233), .B(n239), .C(n232), .Y(n191) );
  ao22d1_hd U478 ( .A(a_m[12]), .B(n242), .C(n3), .D(a[3]), .Y(n234) );
  oa21d1_hd U479 ( .A(n475), .B(n236), .C(n234), .Y(n192) );
  ao22d1_hd U480 ( .A(a_m[10]), .B(n241), .C(n3), .D(a[2]), .Y(n235) );
  oa21d1_hd U481 ( .A(n236), .B(n239), .C(n235), .Y(n193) );
  ao22d1_hd U482 ( .A(a_m[10]), .B(n242), .C(n3), .D(a[1]), .Y(n237) );
  oa21d1_hd U483 ( .A(n475), .B(n240), .C(n237), .Y(n194) );
  ao22d1_hd U484 ( .A(a_m[8]), .B(n241), .C(n3), .D(a[0]), .Y(n238) );
  oa21d1_hd U485 ( .A(n240), .B(n239), .C(n238), .Y(n195) );
  oa21d1_hd U486 ( .A(n475), .B(n243), .C(n731), .Y(n204) );
  nd2bd1_hd U487 ( .AN(n4), .B(n427), .Y(n259) );
  nr4d1_hd U488 ( .A(n248), .B(n245), .C(n3), .D(n259), .Y(n246) );
  nd3d1_hd U489 ( .A(n1), .B(i_Z_ACK), .C(o_Z_STB), .Y(n262) );
  nd3bd1_hd U490 ( .AN(i_RST), .B(n248), .C(n247), .Y(n251) );
  ivd1_hd U491 ( .A(n255), .Y(n250) );
  oa211d1_hd U492 ( .A(n261), .B(n257), .C(n251), .D(n249), .Y(n205) );
  ao22d1_hd U493 ( .A(state[0]), .B(n250), .C(n3), .D(n427), .Y(n252) );
  nr2d1_hd U494 ( .A(n254), .B(n253), .Y(n258) );
  oa22d1_hd U495 ( .A(n258), .B(n257), .C(n256), .D(n255), .Y(n207) );
  ivd1_hd U496 ( .A(o_A_ACK), .Y(n260) );
  ao21d1_hd U497 ( .A(n261), .B(n260), .C(n259), .Y(n208) );
  oa211d1_hd U498 ( .A(n1), .B(o_Z_STB), .C(n427), .D(n262), .Y(n263) );
endmodule


module ads1292_filter ( i_ADS1292_DATA_OUT, i_ADS1292_DATA_VALID, 
        o_ADS1292_FILTERED_DATA, o_ADS1292_FILTERED_DATA_VALID, 
        i_ADS1292_FILTERED_DATA_ACK, i_CLK, i_RSTN );
  input [71:0] i_ADS1292_DATA_OUT;
  output [23:0] o_ADS1292_FILTERED_DATA;
  input i_ADS1292_DATA_VALID, i_ADS1292_FILTERED_DATA_ACK, i_CLK, i_RSTN;
  output o_ADS1292_FILTERED_DATA_VALID;
  wire   r_converter_i2f_a_stb, w_converter_i2f_a_ack, w_converter_i2f_z_stb,
         r_converter_i2f_z_ack, r_iir_lpf_x_valid, w_iir_lpf_x_ready,
         w_iir_lpf_y_valid, r_iir_lpf_y_ack, r_iir_notch_x_valid,
         w_iir_notch_x_ready, w_iir_notch_y_valid, r_iir_notch_y_ack,
         r_iir_hpf_x_valid, w_iir_hpf_x_ready, w_iir_hpf_y_valid,
         r_iir_hpf_y_ack, r_converter_f2i_a_stb, w_converter_f2i_a_ack,
         w_converter_f2i_z_stb, r_converter_f2i_z_ack, r_counter_0_, N31, n1,
         n2, n3, n4, n5, n6, n7, n8, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n255, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8;
  wire   [31:7] r_converter_i2f_a;
  wire   [31:0] w_converter_i2f_z;
  wire   [31:0] r_iir_lpf_x;
  wire   [31:0] w_iir_lpf_y;
  wire   [31:0] r_iir_notch_x;
  wire   [31:0] w_iir_notch_y;
  wire   [31:0] r_iir_hpf_x;
  wire   [31:0] w_iir_hpf_y;
  wire   [31:0] r_converter_f2i_a;
  wire   [31:8] w_converter_f2i_z;

  converter_i2f converter_i2f ( .i_A({r_converter_i2f_a[31:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .i_A_STB(r_converter_i2f_a_stb), 
        .o_A_ACK(w_converter_i2f_a_ack), .o_Z(w_converter_i2f_z), .o_Z_STB(
        w_converter_i2f_z_stb), .i_Z_ACK(r_converter_i2f_z_ack), .i_CLK(i_CLK), 
        .i_RST(N31) );
  iir_lpf iir_lpf ( .i_X_DATA(r_iir_lpf_x), .i_X_DATA_VALID(r_iir_lpf_x_valid), 
        .o_X_DATA_READY(w_iir_lpf_x_ready), .o_Y_DATA(w_iir_lpf_y), 
        .o_Y_DATA_VALID(w_iir_lpf_y_valid), .i_Y_ACK(r_iir_lpf_y_ack), .i_CLK(
        i_CLK), .i_RSTN(i_RSTN) );
  iir_notch iir_notch ( .i_X_DATA(r_iir_notch_x), .i_X_DATA_VALID(
        r_iir_notch_x_valid), .o_X_DATA_READY(w_iir_notch_x_ready), .o_Y_DATA(
        w_iir_notch_y), .o_Y_DATA_VALID(w_iir_notch_y_valid), .i_Y_ACK(
        r_iir_notch_y_ack), .i_CLK(i_CLK), .i_RSTN(i_RSTN) );
  iir_hpf iir_hpf ( .i_X_DATA(r_iir_hpf_x), .i_X_DATA_VALID(r_iir_hpf_x_valid), 
        .o_X_DATA_READY(w_iir_hpf_x_ready), .o_Y_DATA(w_iir_hpf_y), 
        .o_Y_DATA_VALID(w_iir_hpf_y_valid), .i_Y_ACK(r_iir_hpf_y_ack), .i_CLK(
        i_CLK), .i_RSTN(i_RSTN) );
  converter_f2i converter_f2i ( .i_A(r_converter_f2i_a), .i_A_STB(
        r_converter_f2i_a_stb), .o_A_ACK(w_converter_f2i_a_ack), .o_Z({
        w_converter_f2i_z, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8}), .o_Z_STB(w_converter_f2i_z_stb), .i_Z_ACK(r_converter_f2i_z_ack), .i_CLK(
        i_CLK), .i_RST(N31) );
  fd3qd1_hd r_pstate_reg_1_ ( .D(n7), .CK(i_CLK), .SN(i_RSTN), .Q(n8) );
  fd3qd1_hd r_pstate_reg_0_ ( .D(n5), .CK(i_CLK), .SN(i_RSTN), .Q(n6) );
  fd3qd1_hd r_counter_reg_2_ ( .D(n3), .CK(i_CLK), .SN(i_RSTN), .Q(n4) );
  fd3qd1_hd r_counter_reg_1_ ( .D(n1), .CK(i_CLK), .SN(i_RSTN), .Q(n2) );
  ivd1_hd U242 ( .A(i_RSTN), .Y(N31) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_0_ ( .D(n112), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[0]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_1_ ( .D(n111), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[1]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_2_ ( .D(n110), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[2]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_3_ ( .D(n109), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[3]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_4_ ( .D(n108), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[4]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_5_ ( .D(n107), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[5]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_6_ ( .D(n106), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[6]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_7_ ( .D(n105), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[7]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_8_ ( .D(n104), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[8]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_9_ ( .D(n103), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[9]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_10_ ( .D(n102), .CK(i_CLK), .RN(i_RSTN), .Q(o_ADS1292_FILTERED_DATA[10]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_11_ ( .D(n101), .CK(i_CLK), .RN(i_RSTN), .Q(o_ADS1292_FILTERED_DATA[11]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_12_ ( .D(n100), .CK(i_CLK), .RN(i_RSTN), .Q(o_ADS1292_FILTERED_DATA[12]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_13_ ( .D(n99), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[13]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_14_ ( .D(n98), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[14]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_15_ ( .D(n97), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[15]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_16_ ( .D(n96), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[16]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_17_ ( .D(n95), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[17]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_18_ ( .D(n94), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[18]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_19_ ( .D(n93), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[19]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_20_ ( .D(n92), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[20]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_21_ ( .D(n91), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[21]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_22_ ( .D(n90), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[22]) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_reg_23_ ( .D(n89), .CK(i_CLK), .RN(i_RSTN), 
        .Q(o_ADS1292_FILTERED_DATA[23]) );
  fd2qd1_hd r_converter_i2f_a_reg_8_ ( .D(n282), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[8]) );
  fd2qd1_hd r_converter_i2f_a_reg_9_ ( .D(n281), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[9]) );
  fd2qd1_hd r_converter_i2f_a_reg_10_ ( .D(n280), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[10]) );
  fd2qd1_hd r_converter_i2f_a_reg_11_ ( .D(n279), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[11]) );
  fd2qd1_hd r_converter_i2f_a_reg_12_ ( .D(n278), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[12]) );
  fd2qd1_hd r_converter_i2f_a_reg_13_ ( .D(n277), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[13]) );
  fd2qd1_hd r_converter_i2f_a_reg_14_ ( .D(n276), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[14]) );
  fd2qd1_hd r_converter_i2f_a_reg_15_ ( .D(n275), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[15]) );
  fd2qd1_hd r_converter_i2f_a_reg_16_ ( .D(n274), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[16]) );
  fd2qd1_hd r_converter_i2f_a_reg_17_ ( .D(n273), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[17]) );
  fd2qd1_hd r_converter_i2f_a_reg_18_ ( .D(n272), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[18]) );
  fd2qd1_hd r_converter_i2f_a_reg_19_ ( .D(n271), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[19]) );
  fd2qd1_hd r_converter_i2f_a_reg_20_ ( .D(n270), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[20]) );
  fd2qd1_hd r_converter_i2f_a_reg_21_ ( .D(n269), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[21]) );
  fd2qd1_hd r_converter_i2f_a_reg_22_ ( .D(n268), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[22]) );
  fd2qd1_hd r_converter_i2f_a_reg_23_ ( .D(n267), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[23]) );
  fd2qd1_hd r_converter_i2f_a_reg_24_ ( .D(n266), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[24]) );
  fd2qd1_hd r_converter_i2f_a_reg_25_ ( .D(n265), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[25]) );
  fd2qd1_hd r_converter_i2f_a_reg_26_ ( .D(n264), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[26]) );
  fd2qd1_hd r_converter_i2f_a_reg_27_ ( .D(n263), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[27]) );
  fd2qd1_hd r_converter_i2f_a_reg_28_ ( .D(n262), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[28]) );
  fd2qd1_hd r_converter_i2f_a_reg_29_ ( .D(n261), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[29]) );
  fd2qd1_hd r_converter_i2f_a_reg_30_ ( .D(n260), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[30]) );
  fd2qd1_hd r_converter_i2f_a_reg_31_ ( .D(n259), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a[31]) );
  fd2qd1_hd r_converter_f2i_a_reg_0_ ( .D(n144), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[0]) );
  fd2qd1_hd r_converter_f2i_a_reg_1_ ( .D(n143), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[1]) );
  fd2qd1_hd r_converter_f2i_a_reg_2_ ( .D(n142), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[2]) );
  fd2qd1_hd r_converter_f2i_a_reg_3_ ( .D(n141), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[3]) );
  fd2qd1_hd r_converter_f2i_a_reg_4_ ( .D(n140), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[4]) );
  fd2qd1_hd r_converter_f2i_a_reg_5_ ( .D(n139), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[5]) );
  fd2qd1_hd r_converter_f2i_a_reg_6_ ( .D(n138), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[6]) );
  fd2qd1_hd r_converter_f2i_a_reg_7_ ( .D(n137), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[7]) );
  fd2qd1_hd r_converter_f2i_a_reg_8_ ( .D(n136), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[8]) );
  fd2qd1_hd r_converter_f2i_a_reg_9_ ( .D(n135), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[9]) );
  fd2qd1_hd r_converter_f2i_a_reg_10_ ( .D(n134), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[10]) );
  fd2qd1_hd r_converter_f2i_a_reg_11_ ( .D(n133), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[11]) );
  fd2qd1_hd r_converter_f2i_a_reg_12_ ( .D(n132), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[12]) );
  fd2qd1_hd r_converter_f2i_a_reg_13_ ( .D(n131), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[13]) );
  fd2qd1_hd r_converter_f2i_a_reg_14_ ( .D(n130), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[14]) );
  fd2qd1_hd r_converter_f2i_a_reg_15_ ( .D(n129), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[15]) );
  fd2qd1_hd r_converter_f2i_a_reg_16_ ( .D(n128), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[16]) );
  fd2qd1_hd r_converter_f2i_a_reg_17_ ( .D(n127), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[17]) );
  fd2qd1_hd r_converter_f2i_a_reg_18_ ( .D(n126), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[18]) );
  fd2qd1_hd r_converter_f2i_a_reg_19_ ( .D(n125), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[19]) );
  fd2qd1_hd r_converter_f2i_a_reg_20_ ( .D(n124), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[20]) );
  fd2qd1_hd r_converter_f2i_a_reg_21_ ( .D(n123), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[21]) );
  fd2qd1_hd r_converter_f2i_a_reg_22_ ( .D(n122), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[22]) );
  fd2qd1_hd r_converter_f2i_a_reg_23_ ( .D(n121), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[23]) );
  fd2qd1_hd r_converter_f2i_a_reg_24_ ( .D(n120), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[24]) );
  fd2qd1_hd r_converter_f2i_a_reg_25_ ( .D(n119), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[25]) );
  fd2qd1_hd r_converter_f2i_a_reg_26_ ( .D(n118), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[26]) );
  fd2qd1_hd r_converter_f2i_a_reg_27_ ( .D(n117), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[27]) );
  fd2qd1_hd r_converter_f2i_a_reg_28_ ( .D(n116), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[28]) );
  fd2qd1_hd r_converter_f2i_a_reg_29_ ( .D(n115), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[29]) );
  fd2qd1_hd r_converter_f2i_a_reg_30_ ( .D(n114), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[30]) );
  fd2qd1_hd r_converter_f2i_a_reg_31_ ( .D(n113), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a[31]) );
  fd2qd1_hd r_iir_lpf_x_reg_28_ ( .D(n219), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[28]) );
  fd2qd1_hd r_iir_lpf_x_reg_29_ ( .D(n218), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[29]) );
  fd2qd1_hd r_iir_lpf_x_reg_30_ ( .D(n217), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[30]) );
  fd2qd1_hd r_iir_lpf_x_reg_31_ ( .D(n216), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[31]) );
  fd2qd1_hd r_iir_lpf_x_reg_0_ ( .D(n247), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[0]) );
  fd2qd1_hd r_iir_lpf_x_reg_1_ ( .D(n246), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[1]) );
  fd2qd1_hd r_iir_lpf_x_reg_2_ ( .D(n245), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[2]) );
  fd2qd1_hd r_iir_lpf_x_reg_3_ ( .D(n244), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[3]) );
  fd2qd1_hd r_iir_lpf_x_reg_4_ ( .D(n243), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[4]) );
  fd2qd1_hd r_iir_lpf_x_reg_5_ ( .D(n242), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[5]) );
  fd2qd1_hd r_iir_lpf_x_reg_6_ ( .D(n241), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[6]) );
  fd2qd1_hd r_iir_lpf_x_reg_7_ ( .D(n240), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[7]) );
  fd2qd1_hd r_iir_lpf_x_reg_8_ ( .D(n239), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[8]) );
  fd2qd1_hd r_iir_lpf_x_reg_9_ ( .D(n238), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[9]) );
  fd2qd1_hd r_iir_lpf_x_reg_10_ ( .D(n237), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[10]) );
  fd2qd1_hd r_iir_lpf_x_reg_11_ ( .D(n236), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[11]) );
  fd2qd1_hd r_iir_lpf_x_reg_12_ ( .D(n235), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[12]) );
  fd2qd1_hd r_iir_lpf_x_reg_13_ ( .D(n234), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[13]) );
  fd2qd1_hd r_iir_lpf_x_reg_14_ ( .D(n233), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[14]) );
  fd2qd1_hd r_iir_lpf_x_reg_15_ ( .D(n232), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[15]) );
  fd2qd1_hd r_iir_lpf_x_reg_16_ ( .D(n231), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[16]) );
  fd2qd1_hd r_iir_lpf_x_reg_17_ ( .D(n230), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[17]) );
  fd2qd1_hd r_iir_lpf_x_reg_18_ ( .D(n229), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[18]) );
  fd2qd1_hd r_iir_lpf_x_reg_19_ ( .D(n228), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[19]) );
  fd2qd1_hd r_iir_lpf_x_reg_20_ ( .D(n227), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[20]) );
  fd2qd1_hd r_iir_lpf_x_reg_21_ ( .D(n226), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[21]) );
  fd2qd1_hd r_iir_lpf_x_reg_22_ ( .D(n225), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[22]) );
  fd2qd1_hd r_iir_lpf_x_reg_23_ ( .D(n224), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[23]) );
  fd2qd1_hd r_iir_lpf_x_reg_24_ ( .D(n223), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[24]) );
  fd2qd1_hd r_iir_lpf_x_reg_25_ ( .D(n222), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[25]) );
  fd2qd1_hd r_iir_lpf_x_reg_26_ ( .D(n221), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[26]) );
  fd2qd1_hd r_iir_lpf_x_reg_27_ ( .D(n220), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x[27]) );
  fd2qd1_hd r_iir_notch_x_reg_0_ ( .D(n213), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[0]) );
  fd2qd1_hd r_iir_notch_x_reg_1_ ( .D(n212), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[1]) );
  fd2qd1_hd r_iir_notch_x_reg_2_ ( .D(n211), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[2]) );
  fd2qd1_hd r_iir_notch_x_reg_3_ ( .D(n210), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[3]) );
  fd2qd1_hd r_iir_notch_x_reg_4_ ( .D(n209), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[4]) );
  fd2qd1_hd r_iir_notch_x_reg_5_ ( .D(n208), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[5]) );
  fd2qd1_hd r_iir_notch_x_reg_6_ ( .D(n207), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[6]) );
  fd2qd1_hd r_iir_notch_x_reg_7_ ( .D(n206), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[7]) );
  fd2qd1_hd r_iir_notch_x_reg_8_ ( .D(n205), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[8]) );
  fd2qd1_hd r_iir_notch_x_reg_9_ ( .D(n204), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[9]) );
  fd2qd1_hd r_iir_notch_x_reg_10_ ( .D(n203), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[10]) );
  fd2qd1_hd r_iir_notch_x_reg_11_ ( .D(n202), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[11]) );
  fd2qd1_hd r_iir_notch_x_reg_12_ ( .D(n201), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[12]) );
  fd2qd1_hd r_iir_notch_x_reg_13_ ( .D(n200), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[13]) );
  fd2qd1_hd r_iir_notch_x_reg_14_ ( .D(n199), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[14]) );
  fd2qd1_hd r_iir_notch_x_reg_15_ ( .D(n198), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[15]) );
  fd2qd1_hd r_iir_notch_x_reg_16_ ( .D(n197), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[16]) );
  fd2qd1_hd r_iir_notch_x_reg_17_ ( .D(n196), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[17]) );
  fd2qd1_hd r_iir_notch_x_reg_18_ ( .D(n195), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[18]) );
  fd2qd1_hd r_iir_notch_x_reg_19_ ( .D(n194), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[19]) );
  fd2qd1_hd r_iir_notch_x_reg_20_ ( .D(n193), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[20]) );
  fd2qd1_hd r_iir_notch_x_reg_21_ ( .D(n192), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[21]) );
  fd2qd1_hd r_iir_notch_x_reg_22_ ( .D(n191), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[22]) );
  fd2qd1_hd r_iir_notch_x_reg_23_ ( .D(n190), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[23]) );
  fd2qd1_hd r_iir_notch_x_reg_24_ ( .D(n189), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[24]) );
  fd2qd1_hd r_iir_notch_x_reg_25_ ( .D(n188), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[25]) );
  fd2qd1_hd r_iir_notch_x_reg_26_ ( .D(n187), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[26]) );
  fd2qd1_hd r_iir_notch_x_reg_27_ ( .D(n186), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[27]) );
  fd2qd1_hd r_iir_notch_x_reg_28_ ( .D(n185), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[28]) );
  fd2qd1_hd r_iir_notch_x_reg_29_ ( .D(n184), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[29]) );
  fd2qd1_hd r_iir_notch_x_reg_30_ ( .D(n183), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[30]) );
  fd2qd1_hd r_iir_notch_x_reg_31_ ( .D(n182), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x[31]) );
  fd2qd1_hd r_iir_hpf_x_reg_0_ ( .D(n180), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[0]) );
  fd2qd1_hd r_iir_hpf_x_reg_1_ ( .D(n179), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[1]) );
  fd2qd1_hd r_iir_hpf_x_reg_2_ ( .D(n178), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[2]) );
  fd2qd1_hd r_iir_hpf_x_reg_3_ ( .D(n177), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[3]) );
  fd2qd1_hd r_iir_hpf_x_reg_4_ ( .D(n176), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[4]) );
  fd2qd1_hd r_iir_hpf_x_reg_5_ ( .D(n175), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[5]) );
  fd2qd1_hd r_iir_hpf_x_reg_6_ ( .D(n174), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[6]) );
  fd2qd1_hd r_iir_hpf_x_reg_7_ ( .D(n173), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[7]) );
  fd2qd1_hd r_iir_hpf_x_reg_8_ ( .D(n172), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[8]) );
  fd2qd1_hd r_iir_hpf_x_reg_9_ ( .D(n171), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[9]) );
  fd2qd1_hd r_iir_hpf_x_reg_10_ ( .D(n170), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[10]) );
  fd2qd1_hd r_iir_hpf_x_reg_11_ ( .D(n169), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[11]) );
  fd2qd1_hd r_iir_hpf_x_reg_12_ ( .D(n168), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[12]) );
  fd2qd1_hd r_iir_hpf_x_reg_13_ ( .D(n167), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[13]) );
  fd2qd1_hd r_iir_hpf_x_reg_14_ ( .D(n166), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[14]) );
  fd2qd1_hd r_iir_hpf_x_reg_15_ ( .D(n165), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[15]) );
  fd2qd1_hd r_iir_hpf_x_reg_16_ ( .D(n164), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[16]) );
  fd2qd1_hd r_iir_hpf_x_reg_17_ ( .D(n163), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[17]) );
  fd2qd1_hd r_iir_hpf_x_reg_18_ ( .D(n162), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[18]) );
  fd2qd1_hd r_iir_hpf_x_reg_19_ ( .D(n161), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[19]) );
  fd2qd1_hd r_iir_hpf_x_reg_20_ ( .D(n160), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[20]) );
  fd2qd1_hd r_iir_hpf_x_reg_21_ ( .D(n159), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[21]) );
  fd2qd1_hd r_iir_hpf_x_reg_22_ ( .D(n158), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[22]) );
  fd2qd1_hd r_iir_hpf_x_reg_23_ ( .D(n157), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[23]) );
  fd2qd1_hd r_iir_hpf_x_reg_24_ ( .D(n156), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[24]) );
  fd2qd1_hd r_iir_hpf_x_reg_25_ ( .D(n155), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[25]) );
  fd2qd1_hd r_iir_hpf_x_reg_26_ ( .D(n154), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[26]) );
  fd2qd1_hd r_iir_hpf_x_reg_27_ ( .D(n153), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[27]) );
  fd2qd1_hd r_iir_hpf_x_reg_28_ ( .D(n152), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[28]) );
  fd2qd1_hd r_iir_hpf_x_reg_29_ ( .D(n151), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[29]) );
  fd2qd1_hd r_iir_hpf_x_reg_30_ ( .D(n150), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[30]) );
  fd2qd1_hd r_iir_hpf_x_reg_31_ ( .D(n149), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x[31]) );
  fd2qd1_hd r_converter_i2f_z_ack_reg ( .D(n248), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_z_ack) );
  fd2qd1_hd r_iir_lpf_y_ack_reg ( .D(n214), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_y_ack) );
  fd2qd1_hd r_converter_i2f_a_stb_reg ( .D(n147), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_i2f_a_stb) );
  fd2qd1_hd r_iir_notch_y_ack_reg ( .D(n181), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_y_ack) );
  fd2qd1_hd r_iir_hpf_y_ack_reg ( .D(n145), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_y_ack) );
  fd2qd1_hd r_converter_f2i_z_ack_reg ( .D(n257), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_z_ack) );
  fd2qd1_hd o_ADS1292_FILTERED_DATA_VALID_reg ( .D(n258), .CK(i_CLK), .RN(
        i_RSTN), .Q(o_ADS1292_FILTERED_DATA_VALID) );
  fd2qd1_hd r_iir_lpf_x_valid_reg ( .D(n215), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_lpf_x_valid) );
  fd2qd1_hd r_iir_hpf_x_valid_reg ( .D(n146), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_hpf_x_valid) );
  fd2qd1_hd r_iir_notch_x_valid_reg ( .D(n148), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_iir_notch_x_valid) );
  fd2qd1_hd r_converter_f2i_a_stb_reg ( .D(n88), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_converter_f2i_a_stb) );
  fd2qd1_hd r_counter_reg_0_ ( .D(n255), .CK(i_CLK), .RN(i_RSTN), .Q(
        r_counter_0_) );
  clknd2d1_hd U293 ( .A(n6), .B(n8), .Y(n293) );
  clknd2d1_hd U294 ( .A(n310), .B(w_iir_hpf_y_valid), .Y(n311) );
  clknd2d1_hd U295 ( .A(n324), .B(w_iir_lpf_y_valid), .Y(n301) );
  clknd2d1_hd U296 ( .A(n322), .B(w_iir_notch_y_valid), .Y(n305) );
  clknd2d1_hd U297 ( .A(n323), .B(w_converter_i2f_z_stb), .Y(n296) );
  clknd2d1_hd U298 ( .A(n4), .B(n2), .Y(n291) );
  clknd2d1_hd U299 ( .A(n341), .B(n293), .Y(n351) );
  clknd2d1_hd U300 ( .A(n4), .B(n348), .Y(n332) );
  clknd2d1_hd U301 ( .A(n334), .B(n327), .Y(n318) );
  clknd2d1_hd U302 ( .A(n322), .B(w_iir_notch_x_ready), .Y(n320) );
  clknd2d1_hd U303 ( .A(n310), .B(w_iir_hpf_x_ready), .Y(n319) );
  clknd2d1_hd U304 ( .A(n317), .B(r_converter_f2i_a_stb), .Y(n316) );
  clknd2d1_hd U305 ( .A(n324), .B(w_iir_lpf_x_ready), .Y(n300) );
  clknd2d1_hd U306 ( .A(n283), .B(n290), .Y(n257) );
  clknd2d1_hd U307 ( .A(i_ADS1292_FILTERED_DATA_ACK), .B(
        o_ADS1292_FILTERED_DATA_VALID), .Y(n289) );
  clknd2d1_hd U308 ( .A(n323), .B(w_converter_i2f_a_ack), .Y(n309) );
  clknd2d1_hd U309 ( .A(n347), .B(n346), .Y(n3) );
  clknd2d1_hd U310 ( .A(n351), .B(n349), .Y(n347) );
  ivd2_hd U311 ( .A(n313), .Y(n314) );
  ivd2_hd U312 ( .A(n303), .Y(n304) );
  ivd2_hd U313 ( .A(n307), .Y(n308) );
  ivd2_hd U314 ( .A(n298), .Y(n299) );
  nr2d4_hd U315 ( .A(r_counter_0_), .B(n287), .Y(n315) );
  scg2d1_hd U316 ( .A(n2), .B(n352), .C(n351), .D(n350), .Y(n1) );
  scg2d1_hd U317 ( .A(n314), .B(w_iir_hpf_y[15]), .C(r_converter_f2i_a[15]), 
        .D(n313), .Y(n129) );
  scg2d1_hd U318 ( .A(n314), .B(w_iir_hpf_y[14]), .C(r_converter_f2i_a[14]), 
        .D(n313), .Y(n130) );
  scg2d1_hd U319 ( .A(n314), .B(w_iir_hpf_y[13]), .C(r_converter_f2i_a[13]), 
        .D(n313), .Y(n131) );
  scg2d1_hd U320 ( .A(n314), .B(w_iir_hpf_y[12]), .C(r_converter_f2i_a[12]), 
        .D(n313), .Y(n132) );
  scg2d1_hd U321 ( .A(n314), .B(w_iir_hpf_y[11]), .C(r_converter_f2i_a[11]), 
        .D(n313), .Y(n133) );
  scg2d1_hd U322 ( .A(n314), .B(w_iir_hpf_y[10]), .C(r_converter_f2i_a[10]), 
        .D(n313), .Y(n134) );
  scg2d1_hd U323 ( .A(n314), .B(w_iir_hpf_y[9]), .C(r_converter_f2i_a[9]), .D(
        n313), .Y(n135) );
  scg2d1_hd U324 ( .A(n314), .B(w_iir_hpf_y[8]), .C(r_converter_f2i_a[8]), .D(
        n313), .Y(n136) );
  scg2d1_hd U325 ( .A(n314), .B(w_iir_hpf_y[7]), .C(r_converter_f2i_a[7]), .D(
        n313), .Y(n137) );
  scg2d1_hd U326 ( .A(n314), .B(w_iir_hpf_y[6]), .C(r_converter_f2i_a[6]), .D(
        n313), .Y(n138) );
  scg2d1_hd U327 ( .A(n314), .B(w_iir_hpf_y[5]), .C(r_converter_f2i_a[5]), .D(
        n313), .Y(n139) );
  scg2d1_hd U328 ( .A(n314), .B(w_iir_hpf_y[4]), .C(r_converter_f2i_a[4]), .D(
        n313), .Y(n140) );
  scg2d1_hd U329 ( .A(n314), .B(w_iir_hpf_y[3]), .C(r_converter_f2i_a[3]), .D(
        n313), .Y(n141) );
  scg2d1_hd U330 ( .A(n314), .B(w_iir_hpf_y[29]), .C(r_converter_f2i_a[29]), 
        .D(n313), .Y(n115) );
  scg2d1_hd U331 ( .A(n314), .B(w_iir_hpf_y[28]), .C(r_converter_f2i_a[28]), 
        .D(n313), .Y(n116) );
  scg2d1_hd U332 ( .A(n314), .B(w_iir_hpf_y[30]), .C(r_converter_f2i_a[30]), 
        .D(n313), .Y(n114) );
  scg2d1_hd U333 ( .A(n314), .B(w_iir_hpf_y[27]), .C(r_converter_f2i_a[27]), 
        .D(n313), .Y(n117) );
  scg2d1_hd U334 ( .A(n314), .B(w_iir_hpf_y[31]), .C(r_converter_f2i_a[31]), 
        .D(n313), .Y(n113) );
  scg2d1_hd U335 ( .A(n314), .B(w_iir_hpf_y[26]), .C(r_converter_f2i_a[26]), 
        .D(n313), .Y(n118) );
  scg2d1_hd U336 ( .A(n314), .B(w_iir_hpf_y[25]), .C(r_converter_f2i_a[25]), 
        .D(n313), .Y(n119) );
  scg2d1_hd U337 ( .A(n314), .B(w_iir_hpf_y[24]), .C(r_converter_f2i_a[24]), 
        .D(n313), .Y(n120) );
  scg2d1_hd U338 ( .A(n314), .B(w_iir_hpf_y[23]), .C(r_converter_f2i_a[23]), 
        .D(n313), .Y(n121) );
  scg2d1_hd U339 ( .A(n314), .B(w_iir_hpf_y[22]), .C(r_converter_f2i_a[22]), 
        .D(n313), .Y(n122) );
  or2d1_hd U340 ( .A(n349), .B(n348), .Y(n350) );
  scg2d1_hd U341 ( .A(n314), .B(w_iir_hpf_y[21]), .C(r_converter_f2i_a[21]), 
        .D(n313), .Y(n123) );
  scg2d1_hd U342 ( .A(n314), .B(w_iir_hpf_y[20]), .C(r_converter_f2i_a[20]), 
        .D(n313), .Y(n124) );
  scg2d1_hd U343 ( .A(n314), .B(w_iir_hpf_y[19]), .C(r_converter_f2i_a[19]), 
        .D(n313), .Y(n125) );
  scg2d1_hd U344 ( .A(n314), .B(w_iir_hpf_y[18]), .C(r_converter_f2i_a[18]), 
        .D(n313), .Y(n126) );
  scg2d1_hd U345 ( .A(n314), .B(w_iir_hpf_y[17]), .C(r_converter_f2i_a[17]), 
        .D(n313), .Y(n127) );
  scg2d1_hd U346 ( .A(n314), .B(w_iir_hpf_y[16]), .C(r_converter_f2i_a[16]), 
        .D(n313), .Y(n128) );
  scg2d1_hd U347 ( .A(n314), .B(w_iir_hpf_y[0]), .C(r_converter_f2i_a[0]), .D(
        n313), .Y(n144) );
  scg2d1_hd U348 ( .A(n314), .B(w_iir_hpf_y[1]), .C(r_converter_f2i_a[1]), .D(
        n313), .Y(n143) );
  scg2d1_hd U349 ( .A(n314), .B(w_iir_hpf_y[2]), .C(r_converter_f2i_a[2]), .D(
        n313), .Y(n142) );
  scg2d1_hd U350 ( .A(n304), .B(w_iir_lpf_y[11]), .C(r_iir_notch_x[11]), .D(
        n303), .Y(n202) );
  scg2d1_hd U351 ( .A(n315), .B(w_converter_f2i_z[22]), .C(
        o_ADS1292_FILTERED_DATA[14]), .D(n283), .Y(n98) );
  scg2d1_hd U352 ( .A(n304), .B(w_iir_lpf_y[12]), .C(r_iir_notch_x[12]), .D(
        n303), .Y(n201) );
  scg2d1_hd U353 ( .A(n308), .B(w_iir_notch_y[5]), .C(r_iir_hpf_x[5]), .D(n307), .Y(n175) );
  scg2d1_hd U354 ( .A(n304), .B(w_iir_lpf_y[13]), .C(r_iir_notch_x[13]), .D(
        n303), .Y(n200) );
  scg2d1_hd U355 ( .A(n308), .B(w_iir_notch_y[14]), .C(r_iir_hpf_x[14]), .D(
        n307), .Y(n166) );
  scg2d1_hd U356 ( .A(n308), .B(w_iir_notch_y[19]), .C(r_iir_hpf_x[19]), .D(
        n307), .Y(n161) );
  scg2d1_hd U357 ( .A(n304), .B(w_iir_lpf_y[14]), .C(r_iir_notch_x[14]), .D(
        n303), .Y(n199) );
  scg2d1_hd U358 ( .A(n315), .B(w_converter_f2i_z[23]), .C(
        o_ADS1292_FILTERED_DATA[15]), .D(n283), .Y(n97) );
  scg2d1_hd U359 ( .A(n308), .B(w_iir_notch_y[22]), .C(r_iir_hpf_x[22]), .D(
        n307), .Y(n158) );
  scg2d1_hd U360 ( .A(n304), .B(w_iir_lpf_y[10]), .C(r_iir_notch_x[10]), .D(
        n303), .Y(n203) );
  scg2d1_hd U361 ( .A(n308), .B(w_iir_notch_y[3]), .C(r_iir_hpf_x[3]), .D(n307), .Y(n177) );
  scg2d1_hd U362 ( .A(n304), .B(w_iir_lpf_y[9]), .C(r_iir_notch_x[9]), .D(n303), .Y(n204) );
  scg2d1_hd U363 ( .A(n308), .B(w_iir_notch_y[16]), .C(r_iir_hpf_x[16]), .D(
        n307), .Y(n164) );
  scg2d1_hd U364 ( .A(n308), .B(w_iir_notch_y[21]), .C(r_iir_hpf_x[21]), .D(
        n307), .Y(n159) );
  scg2d1_hd U365 ( .A(n308), .B(w_iir_notch_y[15]), .C(r_iir_hpf_x[15]), .D(
        n307), .Y(n165) );
  scg2d1_hd U366 ( .A(n308), .B(w_iir_notch_y[2]), .C(r_iir_hpf_x[2]), .D(n307), .Y(n178) );
  scg2d1_hd U367 ( .A(n304), .B(w_iir_lpf_y[8]), .C(r_iir_notch_x[8]), .D(n303), .Y(n205) );
  scg2d1_hd U368 ( .A(n315), .B(w_converter_f2i_z[21]), .C(
        o_ADS1292_FILTERED_DATA[13]), .D(n283), .Y(n99) );
  scg2d1_hd U369 ( .A(n308), .B(w_iir_notch_y[0]), .C(r_iir_hpf_x[0]), .D(n307), .Y(n180) );
  scg2d1_hd U370 ( .A(n308), .B(w_iir_notch_y[20]), .C(r_iir_hpf_x[20]), .D(
        n307), .Y(n160) );
  scg2d1_hd U371 ( .A(n308), .B(w_iir_notch_y[1]), .C(r_iir_hpf_x[1]), .D(n307), .Y(n179) );
  scg2d1_hd U372 ( .A(n308), .B(w_iir_notch_y[24]), .C(r_iir_hpf_x[24]), .D(
        n307), .Y(n156) );
  scg2d1_hd U373 ( .A(n315), .B(w_converter_f2i_z[29]), .C(
        o_ADS1292_FILTERED_DATA[21]), .D(n283), .Y(n91) );
  scg2d1_hd U374 ( .A(n304), .B(w_iir_lpf_y[26]), .C(r_iir_notch_x[26]), .D(
        n303), .Y(n187) );
  scg2d1_hd U375 ( .A(n304), .B(w_iir_lpf_y[25]), .C(r_iir_notch_x[25]), .D(
        n303), .Y(n188) );
  scg2d1_hd U376 ( .A(n304), .B(w_iir_lpf_y[24]), .C(r_iir_notch_x[24]), .D(
        n303), .Y(n189) );
  scg2d1_hd U377 ( .A(n315), .B(w_converter_f2i_z[28]), .C(
        o_ADS1292_FILTERED_DATA[20]), .D(n283), .Y(n92) );
  scg2d1_hd U378 ( .A(n308), .B(w_iir_notch_y[25]), .C(r_iir_hpf_x[25]), .D(
        n307), .Y(n155) );
  scg2d1_hd U379 ( .A(n304), .B(w_iir_lpf_y[27]), .C(r_iir_notch_x[27]), .D(
        n303), .Y(n186) );
  scg2d1_hd U380 ( .A(n315), .B(w_converter_f2i_z[27]), .C(
        o_ADS1292_FILTERED_DATA[19]), .D(n283), .Y(n93) );
  scg2d1_hd U381 ( .A(n315), .B(w_converter_f2i_z[30]), .C(
        o_ADS1292_FILTERED_DATA[22]), .D(n283), .Y(n90) );
  scg2d1_hd U382 ( .A(n308), .B(w_iir_notch_y[18]), .C(r_iir_hpf_x[18]), .D(
        n307), .Y(n162) );
  scg2d1_hd U383 ( .A(n315), .B(w_converter_f2i_z[26]), .C(
        o_ADS1292_FILTERED_DATA[18]), .D(n283), .Y(n94) );
  scg2d1_hd U384 ( .A(n315), .B(w_converter_f2i_z[25]), .C(
        o_ADS1292_FILTERED_DATA[17]), .D(n283), .Y(n95) );
  scg2d1_hd U385 ( .A(n304), .B(w_iir_lpf_y[28]), .C(r_iir_notch_x[28]), .D(
        n303), .Y(n185) );
  scg2d1_hd U386 ( .A(n304), .B(w_iir_lpf_y[23]), .C(r_iir_notch_x[23]), .D(
        n303), .Y(n190) );
  scg2d1_hd U387 ( .A(n308), .B(w_iir_notch_y[6]), .C(r_iir_hpf_x[6]), .D(n307), .Y(n174) );
  scg2d1_hd U388 ( .A(n315), .B(w_converter_f2i_z[24]), .C(
        o_ADS1292_FILTERED_DATA[16]), .D(n283), .Y(n96) );
  scg2d1_hd U389 ( .A(n308), .B(w_iir_notch_y[26]), .C(r_iir_hpf_x[26]), .D(
        n307), .Y(n154) );
  scg2d1_hd U390 ( .A(n304), .B(w_iir_lpf_y[22]), .C(r_iir_notch_x[22]), .D(
        n303), .Y(n191) );
  scg2d1_hd U391 ( .A(n308), .B(w_iir_notch_y[27]), .C(r_iir_hpf_x[27]), .D(
        n307), .Y(n153) );
  scg2d1_hd U392 ( .A(n308), .B(w_iir_notch_y[7]), .C(r_iir_hpf_x[7]), .D(n307), .Y(n173) );
  scg2d1_hd U393 ( .A(n304), .B(w_iir_lpf_y[21]), .C(r_iir_notch_x[21]), .D(
        n303), .Y(n192) );
  scg2d1_hd U394 ( .A(n304), .B(w_iir_lpf_y[29]), .C(r_iir_notch_x[29]), .D(
        n303), .Y(n184) );
  scg2d1_hd U395 ( .A(n315), .B(w_converter_f2i_z[31]), .C(
        o_ADS1292_FILTERED_DATA[23]), .D(n283), .Y(n89) );
  scg2d1_hd U396 ( .A(n308), .B(w_iir_notch_y[8]), .C(r_iir_hpf_x[8]), .D(n307), .Y(n172) );
  scg2d1_hd U397 ( .A(n304), .B(w_iir_lpf_y[20]), .C(r_iir_notch_x[20]), .D(
        n303), .Y(n193) );
  scg2d1_hd U398 ( .A(n308), .B(w_iir_notch_y[28]), .C(r_iir_hpf_x[28]), .D(
        n307), .Y(n152) );
  scg2d1_hd U399 ( .A(n308), .B(w_iir_notch_y[9]), .C(r_iir_hpf_x[9]), .D(n307), .Y(n171) );
  scg2d1_hd U400 ( .A(n304), .B(w_iir_lpf_y[19]), .C(r_iir_notch_x[19]), .D(
        n303), .Y(n194) );
  scg2d1_hd U401 ( .A(n304), .B(w_iir_lpf_y[30]), .C(r_iir_notch_x[30]), .D(
        n303), .Y(n183) );
  scg2d1_hd U402 ( .A(n308), .B(w_iir_notch_y[23]), .C(r_iir_hpf_x[23]), .D(
        n307), .Y(n157) );
  scg2d1_hd U403 ( .A(n308), .B(w_iir_notch_y[10]), .C(r_iir_hpf_x[10]), .D(
        n307), .Y(n170) );
  scg2d1_hd U404 ( .A(n308), .B(w_iir_notch_y[29]), .C(r_iir_hpf_x[29]), .D(
        n307), .Y(n151) );
  scg2d1_hd U405 ( .A(n304), .B(w_iir_lpf_y[18]), .C(r_iir_notch_x[18]), .D(
        n303), .Y(n195) );
  scg2d1_hd U406 ( .A(n308), .B(w_iir_notch_y[30]), .C(r_iir_hpf_x[30]), .D(
        n307), .Y(n150) );
  scg2d1_hd U407 ( .A(n308), .B(w_iir_notch_y[11]), .C(r_iir_hpf_x[11]), .D(
        n307), .Y(n169) );
  scg2d1_hd U408 ( .A(n304), .B(w_iir_lpf_y[17]), .C(r_iir_notch_x[17]), .D(
        n303), .Y(n196) );
  scg2d1_hd U409 ( .A(n308), .B(w_iir_notch_y[12]), .C(r_iir_hpf_x[12]), .D(
        n307), .Y(n168) );
  scg2d1_hd U410 ( .A(n308), .B(w_iir_notch_y[17]), .C(r_iir_hpf_x[17]), .D(
        n307), .Y(n163) );
  scg2d1_hd U411 ( .A(n304), .B(w_iir_lpf_y[16]), .C(r_iir_notch_x[16]), .D(
        n303), .Y(n197) );
  scg2d1_hd U412 ( .A(n308), .B(w_iir_notch_y[4]), .C(r_iir_hpf_x[4]), .D(n307), .Y(n176) );
  scg2d1_hd U413 ( .A(n308), .B(w_iir_notch_y[31]), .C(r_iir_hpf_x[31]), .D(
        n307), .Y(n149) );
  scg2d1_hd U414 ( .A(n308), .B(w_iir_notch_y[13]), .C(r_iir_hpf_x[13]), .D(
        n307), .Y(n167) );
  scg2d1_hd U415 ( .A(n304), .B(w_iir_lpf_y[31]), .C(r_iir_notch_x[31]), .D(
        n303), .Y(n182) );
  scg2d1_hd U416 ( .A(n304), .B(w_iir_lpf_y[15]), .C(r_iir_notch_x[15]), .D(
        n303), .Y(n198) );
  scg2d1_hd U417 ( .A(n299), .B(w_converter_i2f_z[26]), .C(r_iir_lpf_x[26]), 
        .D(n298), .Y(n221) );
  scg2d1_hd U418 ( .A(n315), .B(w_converter_f2i_z[13]), .C(
        o_ADS1292_FILTERED_DATA[5]), .D(n283), .Y(n107) );
  scg2d1_hd U419 ( .A(n304), .B(w_iir_lpf_y[4]), .C(r_iir_notch_x[4]), .D(n303), .Y(n209) );
  scg2d1_hd U420 ( .A(n299), .B(w_converter_i2f_z[27]), .C(r_iir_lpf_x[27]), 
        .D(n298), .Y(n220) );
  scg2d1_hd U421 ( .A(n315), .B(w_converter_f2i_z[14]), .C(
        o_ADS1292_FILTERED_DATA[6]), .D(n283), .Y(n106) );
  scg2d1_hd U422 ( .A(n299), .B(w_converter_i2f_z[28]), .C(r_iir_lpf_x[28]), 
        .D(n298), .Y(n219) );
  scg2d1_hd U423 ( .A(n315), .B(w_converter_f2i_z[15]), .C(
        o_ADS1292_FILTERED_DATA[7]), .D(n283), .Y(n105) );
  scg2d1_hd U424 ( .A(n315), .B(w_converter_f2i_z[16]), .C(
        o_ADS1292_FILTERED_DATA[8]), .D(n283), .Y(n104) );
  scg2d1_hd U425 ( .A(n299), .B(w_converter_i2f_z[0]), .C(r_iir_lpf_x[0]), .D(
        n298), .Y(n247) );
  scg2d1_hd U426 ( .A(n304), .B(w_iir_lpf_y[3]), .C(r_iir_notch_x[3]), .D(n303), .Y(n210) );
  scg2d1_hd U427 ( .A(n299), .B(w_converter_i2f_z[1]), .C(r_iir_lpf_x[1]), .D(
        n298), .Y(n246) );
  scg2d1_hd U428 ( .A(n315), .B(w_converter_f2i_z[17]), .C(
        o_ADS1292_FILTERED_DATA[9]), .D(n283), .Y(n103) );
  scg2d1_hd U429 ( .A(n299), .B(w_converter_i2f_z[14]), .C(r_iir_lpf_x[14]), 
        .D(n298), .Y(n233) );
  scg2d1_hd U430 ( .A(n299), .B(w_converter_i2f_z[2]), .C(r_iir_lpf_x[2]), .D(
        n298), .Y(n245) );
  scg2d1_hd U431 ( .A(n299), .B(w_converter_i2f_z[29]), .C(r_iir_lpf_x[29]), 
        .D(n298), .Y(n218) );
  scg2d1_hd U432 ( .A(n315), .B(w_converter_f2i_z[19]), .C(
        o_ADS1292_FILTERED_DATA[11]), .D(n283), .Y(n101) );
  scg2d1_hd U433 ( .A(n299), .B(w_converter_i2f_z[21]), .C(r_iir_lpf_x[21]), 
        .D(n298), .Y(n226) );
  scg2d1_hd U434 ( .A(n299), .B(w_converter_i2f_z[13]), .C(r_iir_lpf_x[13]), 
        .D(n298), .Y(n234) );
  scg2d1_hd U435 ( .A(n299), .B(w_converter_i2f_z[3]), .C(r_iir_lpf_x[3]), .D(
        n298), .Y(n244) );
  scg2d1_hd U436 ( .A(n299), .B(w_converter_i2f_z[30]), .C(r_iir_lpf_x[30]), 
        .D(n298), .Y(n217) );
  scg2d1_hd U437 ( .A(n299), .B(w_converter_i2f_z[20]), .C(r_iir_lpf_x[20]), 
        .D(n298), .Y(n227) );
  scg2d1_hd U438 ( .A(n299), .B(w_converter_i2f_z[4]), .C(r_iir_lpf_x[4]), .D(
        n298), .Y(n243) );
  scg2d1_hd U439 ( .A(n304), .B(w_iir_lpf_y[2]), .C(r_iir_notch_x[2]), .D(n303), .Y(n211) );
  scg2d1_hd U440 ( .A(n299), .B(w_converter_i2f_z[5]), .C(r_iir_lpf_x[5]), .D(
        n298), .Y(n242) );
  scg2d1_hd U441 ( .A(n315), .B(w_converter_f2i_z[18]), .C(
        o_ADS1292_FILTERED_DATA[10]), .D(n283), .Y(n102) );
  scg2d1_hd U442 ( .A(n299), .B(w_converter_i2f_z[31]), .C(r_iir_lpf_x[31]), 
        .D(n298), .Y(n216) );
  scg2d1_hd U443 ( .A(n299), .B(w_converter_i2f_z[6]), .C(r_iir_lpf_x[6]), .D(
        n298), .Y(n241) );
  scg2d1_hd U444 ( .A(n299), .B(w_converter_i2f_z[7]), .C(r_iir_lpf_x[7]), .D(
        n298), .Y(n240) );
  scg2d1_hd U445 ( .A(n299), .B(w_converter_i2f_z[12]), .C(r_iir_lpf_x[12]), 
        .D(n298), .Y(n235) );
  scg2d1_hd U446 ( .A(n299), .B(w_converter_i2f_z[19]), .C(r_iir_lpf_x[19]), 
        .D(n298), .Y(n228) );
  scg2d1_hd U447 ( .A(n299), .B(w_converter_i2f_z[8]), .C(r_iir_lpf_x[8]), .D(
        n298), .Y(n239) );
  scg2d1_hd U448 ( .A(n299), .B(w_converter_i2f_z[9]), .C(r_iir_lpf_x[9]), .D(
        n298), .Y(n238) );
  scg2d1_hd U449 ( .A(n299), .B(w_converter_i2f_z[18]), .C(r_iir_lpf_x[18]), 
        .D(n298), .Y(n229) );
  scg2d1_hd U450 ( .A(n299), .B(w_converter_i2f_z[10]), .C(r_iir_lpf_x[10]), 
        .D(n298), .Y(n237) );
  scg2d1_hd U451 ( .A(n299), .B(w_converter_i2f_z[11]), .C(r_iir_lpf_x[11]), 
        .D(n298), .Y(n236) );
  scg2d1_hd U452 ( .A(n299), .B(w_converter_i2f_z[17]), .C(r_iir_lpf_x[17]), 
        .D(n298), .Y(n230) );
  scg2d1_hd U453 ( .A(n304), .B(w_iir_lpf_y[1]), .C(r_iir_notch_x[1]), .D(n303), .Y(n212) );
  scg2d1_hd U454 ( .A(n299), .B(w_converter_i2f_z[16]), .C(r_iir_lpf_x[16]), 
        .D(n298), .Y(n231) );
  scg2d1_hd U455 ( .A(n299), .B(w_converter_i2f_z[23]), .C(r_iir_lpf_x[23]), 
        .D(n298), .Y(n224) );
  scg2d1_hd U456 ( .A(n304), .B(w_iir_lpf_y[7]), .C(r_iir_notch_x[7]), .D(n303), .Y(n206) );
  scg2d1_hd U457 ( .A(n315), .B(w_converter_f2i_z[8]), .C(
        o_ADS1292_FILTERED_DATA[0]), .D(n283), .Y(n112) );
  scg2d1_hd U458 ( .A(n315), .B(w_converter_f2i_z[9]), .C(
        o_ADS1292_FILTERED_DATA[1]), .D(n283), .Y(n111) );
  scg2d1_hd U459 ( .A(n304), .B(w_iir_lpf_y[6]), .C(r_iir_notch_x[6]), .D(n303), .Y(n207) );
  scg2d1_hd U460 ( .A(n315), .B(w_converter_f2i_z[10]), .C(
        o_ADS1292_FILTERED_DATA[2]), .D(n283), .Y(n110) );
  scg2d1_hd U461 ( .A(n299), .B(w_converter_i2f_z[24]), .C(r_iir_lpf_x[24]), 
        .D(n298), .Y(n223) );
  scg2d1_hd U462 ( .A(n304), .B(w_iir_lpf_y[5]), .C(r_iir_notch_x[5]), .D(n303), .Y(n208) );
  scg2d1_hd U463 ( .A(n315), .B(w_converter_f2i_z[12]), .C(
        o_ADS1292_FILTERED_DATA[4]), .D(n283), .Y(n108) );
  scg2d1_hd U464 ( .A(n315), .B(w_converter_f2i_z[11]), .C(
        o_ADS1292_FILTERED_DATA[3]), .D(n283), .Y(n109) );
  scg2d1_hd U465 ( .A(n299), .B(w_converter_i2f_z[25]), .C(r_iir_lpf_x[25]), 
        .D(n298), .Y(n222) );
  scg2d1_hd U466 ( .A(n315), .B(w_converter_f2i_z[20]), .C(
        o_ADS1292_FILTERED_DATA[12]), .D(n283), .Y(n100) );
  scg2d1_hd U467 ( .A(n299), .B(w_converter_i2f_z[22]), .C(r_iir_lpf_x[22]), 
        .D(n298), .Y(n225) );
  scg2d1_hd U468 ( .A(n299), .B(w_converter_i2f_z[15]), .C(r_iir_lpf_x[15]), 
        .D(n298), .Y(n232) );
  scg2d1_hd U469 ( .A(n304), .B(w_iir_lpf_y[0]), .C(r_iir_notch_x[0]), .D(n303), .Y(n213) );
  nd2d2_hd U470 ( .A(n342), .B(n312), .Y(n313) );
  nd2d2_hd U471 ( .A(n342), .B(n306), .Y(n307) );
  nd2d2_hd U472 ( .A(n342), .B(n302), .Y(n303) );
  scg2d1_hd U473 ( .A(n284), .B(i_ADS1292_DATA_OUT[12]), .C(
        r_converter_i2f_a[20]), .D(n340), .Y(n270) );
  scg2d1_hd U474 ( .A(n284), .B(i_ADS1292_DATA_OUT[11]), .C(
        r_converter_i2f_a[19]), .D(n340), .Y(n271) );
  scg2d1_hd U475 ( .A(n284), .B(i_ADS1292_DATA_OUT[1]), .C(
        r_converter_i2f_a[9]), .D(n340), .Y(n281) );
  scg2d1_hd U476 ( .A(n284), .B(i_ADS1292_DATA_OUT[0]), .C(
        r_converter_i2f_a[8]), .D(n340), .Y(n282) );
  nd2d2_hd U477 ( .A(n342), .B(n297), .Y(n298) );
  scg2d1_hd U478 ( .A(n284), .B(i_ADS1292_DATA_OUT[13]), .C(
        r_converter_i2f_a[21]), .D(n340), .Y(n269) );
  scg2d1_hd U479 ( .A(n284), .B(i_ADS1292_DATA_OUT[23]), .C(
        r_converter_i2f_a[31]), .D(n340), .Y(n259) );
  scg2d1_hd U480 ( .A(n284), .B(i_ADS1292_DATA_OUT[22]), .C(
        r_converter_i2f_a[30]), .D(n340), .Y(n260) );
  scg2d1_hd U481 ( .A(n284), .B(i_ADS1292_DATA_OUT[21]), .C(
        r_converter_i2f_a[29]), .D(n340), .Y(n261) );
  scg2d1_hd U482 ( .A(n284), .B(i_ADS1292_DATA_OUT[20]), .C(
        r_converter_i2f_a[28]), .D(n340), .Y(n262) );
  scg2d1_hd U483 ( .A(n284), .B(i_ADS1292_DATA_OUT[19]), .C(
        r_converter_i2f_a[27]), .D(n340), .Y(n263) );
  scg2d1_hd U484 ( .A(n284), .B(i_ADS1292_DATA_OUT[18]), .C(
        r_converter_i2f_a[26]), .D(n340), .Y(n264) );
  scg2d1_hd U485 ( .A(n284), .B(i_ADS1292_DATA_OUT[17]), .C(
        r_converter_i2f_a[25]), .D(n340), .Y(n265) );
  scg2d1_hd U486 ( .A(n284), .B(i_ADS1292_DATA_OUT[16]), .C(
        r_converter_i2f_a[24]), .D(n340), .Y(n266) );
  scg2d1_hd U487 ( .A(n284), .B(i_ADS1292_DATA_OUT[15]), .C(
        r_converter_i2f_a[23]), .D(n340), .Y(n267) );
  scg2d1_hd U488 ( .A(n284), .B(i_ADS1292_DATA_OUT[14]), .C(
        r_converter_i2f_a[22]), .D(n340), .Y(n268) );
  scg2d1_hd U489 ( .A(n284), .B(i_ADS1292_DATA_OUT[10]), .C(
        r_converter_i2f_a[18]), .D(n340), .Y(n272) );
  scg2d1_hd U490 ( .A(n284), .B(i_ADS1292_DATA_OUT[4]), .C(
        r_converter_i2f_a[12]), .D(n340), .Y(n278) );
  scg2d1_hd U491 ( .A(n284), .B(i_ADS1292_DATA_OUT[2]), .C(
        r_converter_i2f_a[10]), .D(n340), .Y(n280) );
  scg2d1_hd U492 ( .A(n284), .B(i_ADS1292_DATA_OUT[5]), .C(
        r_converter_i2f_a[13]), .D(n340), .Y(n277) );
  scg2d1_hd U493 ( .A(n284), .B(i_ADS1292_DATA_OUT[6]), .C(
        r_converter_i2f_a[14]), .D(n340), .Y(n276) );
  scg2d1_hd U494 ( .A(n284), .B(i_ADS1292_DATA_OUT[7]), .C(
        r_converter_i2f_a[15]), .D(n340), .Y(n275) );
  scg2d1_hd U495 ( .A(n284), .B(i_ADS1292_DATA_OUT[8]), .C(
        r_converter_i2f_a[16]), .D(n340), .Y(n274) );
  scg2d1_hd U496 ( .A(n284), .B(i_ADS1292_DATA_OUT[9]), .C(
        r_converter_i2f_a[17]), .D(n340), .Y(n273) );
  scg2d1_hd U497 ( .A(n284), .B(i_ADS1292_DATA_OUT[3]), .C(
        r_converter_i2f_a[11]), .D(n340), .Y(n279) );
  ivd2_hd U498 ( .A(n284), .Y(n340) );
  clknd2d2_hd U499 ( .A(n6), .B(n285), .Y(n328) );
  ivd2_hd U500 ( .A(n288), .Y(n342) );
  ivd1_hd U501 ( .A(n332), .Y(n310) );
  ivd1_hd U502 ( .A(n328), .Y(n295) );
  oa21d1_hd U503 ( .A(n328), .B(n296), .C(n342), .Y(n297) );
  oa21d1_hd U504 ( .A(n328), .B(n305), .C(n342), .Y(n306) );
  oa21d1_hd U505 ( .A(n328), .B(n301), .C(n342), .Y(n302) );
  oa21d1_hd U506 ( .A(n328), .B(n311), .C(n342), .Y(n312) );
  ad2bd2_hd U507 ( .B(i_ADS1292_DATA_VALID), .AN(n293), .Y(n284) );
  nr2d1_hd U508 ( .A(n6), .B(n285), .Y(n288) );
  ivd2_hd U509 ( .A(n315), .Y(n283) );
  nr2d1_hd U510 ( .A(n294), .B(n291), .Y(n324) );
  ivd1_hd U511 ( .A(n4), .Y(n327) );
  ivd1_hd U512 ( .A(n8), .Y(n285) );
  nd4d1_hd U513 ( .A(n2), .B(n295), .C(w_converter_f2i_z_stb), .D(n327), .Y(
        n287) );
  ivd1_hd U514 ( .A(r_counter_0_), .Y(n294) );
  nr2d1_hd U515 ( .A(r_counter_0_), .B(n291), .Y(n323) );
  nr2d1_hd U516 ( .A(n294), .B(n2), .Y(n348) );
  nr3d1_hd U517 ( .A(n2), .B(r_counter_0_), .C(n327), .Y(n322) );
  nr3d1_hd U518 ( .A(n325), .B(n327), .C(n326), .Y(n329) );
  nr3d1_hd U519 ( .A(n337), .B(n339), .C(n338), .Y(n343) );
  ao211d1_hd U521 ( .A(i_ADS1292_FILTERED_DATA_ACK), .B(
        o_ADS1292_FILTERED_DATA_VALID), .C(n6), .D(n8), .Y(n345) );
  oa21d1_hd U522 ( .A(n288), .B(n295), .C(o_ADS1292_FILTERED_DATA_VALID), .Y(
        n286) );
  nd2bd1_hd U523 ( .AN(n345), .B(n286), .Y(n258) );
  oa211d1_hd U524 ( .A(n6), .B(n289), .C(r_converter_f2i_z_ack), .D(n342), .Y(
        n290) );
  nd4d1_hd U525 ( .A(n305), .B(n311), .C(n296), .D(n301), .Y(n292) );
  ao21d1_hd U526 ( .A(n295), .B(n292), .C(n315), .Y(n341) );
  nd3d1_hd U527 ( .A(n295), .B(n4), .C(n351), .Y(n349) );
  ao22d1_hd U528 ( .A(r_counter_0_), .B(n351), .C(n349), .D(n294), .Y(n255) );
  ao22ad1_hd U529 ( .A(n328), .B(n297), .C(n297), .D(r_converter_i2f_z_ack), 
        .Y(n248) );
  oa22ad1_hd U530 ( .A(n342), .B(n300), .C(n328), .D(r_iir_lpf_x_valid), .Y(
        n215) );
  ao22ad1_hd U531 ( .A(n328), .B(n302), .C(n302), .D(r_iir_lpf_y_ack), .Y(n214) );
  ao22ad1_hd U532 ( .A(n328), .B(n306), .C(n306), .D(r_iir_notch_y_ack), .Y(
        n181) );
  oa22ad1_hd U533 ( .A(n342), .B(n320), .C(n328), .D(r_iir_notch_x_valid), .Y(
        n148) );
  oa22ad1_hd U534 ( .A(n342), .B(n309), .C(n328), .D(r_converter_i2f_a_stb), 
        .Y(n147) );
  oa22ad1_hd U535 ( .A(n342), .B(n319), .C(n328), .D(r_iir_hpf_x_valid), .Y(
        n146) );
  ao22ad1_hd U536 ( .A(n328), .B(n312), .C(n312), .D(r_iir_hpf_y_ack), .Y(n145) );
  scg12d1_hd U537 ( .A(n2), .B(w_converter_f2i_a_ack), .C(r_counter_0_), .Y(
        n334) );
  scg20d1_hd U538 ( .A(n318), .B(n342), .C(n295), .Y(n317) );
  oa21d1_hd U539 ( .A(n342), .B(n317), .C(n316), .Y(n88) );
  ao22d1_hd U540 ( .A(n323), .B(w_converter_i2f_a_ack), .C(n324), .D(
        w_iir_lpf_x_ready), .Y(n321) );
  nd4d1_hd U541 ( .A(n321), .B(n320), .C(n319), .D(n318), .Y(n331) );
  ivd1_hd U542 ( .A(n322), .Y(n333) );
  ivd1_hd U543 ( .A(n323), .Y(n336) );
  oa22d1_hd U544 ( .A(w_iir_notch_y_valid), .B(n333), .C(w_converter_i2f_z_stb), .D(n336), .Y(n326) );
  ivd1_hd U545 ( .A(n324), .Y(n335) );
  oa22d1_hd U546 ( .A(w_iir_hpf_y_valid), .B(n332), .C(w_iir_lpf_y_valid), .D(
        n335), .Y(n325) );
  nr2d1_hd U547 ( .A(n329), .B(n328), .Y(n330) );
  ao211d1_hd U548 ( .A(n288), .B(n331), .C(n345), .D(n330), .Y(n7) );
  nr2d1_hd U549 ( .A(w_iir_hpf_x_ready), .B(n332), .Y(n339) );
  oa22d1_hd U550 ( .A(n4), .B(n334), .C(w_iir_notch_x_ready), .D(n333), .Y(
        n338) );
  oa22d1_hd U551 ( .A(w_converter_i2f_a_ack), .B(n336), .C(w_iir_lpf_x_ready), 
        .D(n335), .Y(n337) );
  oa211d1_hd U552 ( .A(n343), .B(n342), .C(n341), .D(n340), .Y(n344) );
  nr2d1_hd U553 ( .A(n345), .B(n344), .Y(n5) );
  nd2bd1_hd U554 ( .AN(n349), .B(r_counter_0_), .Y(n352) );
  oa21d1_hd U555 ( .A(n2), .B(n352), .C(n4), .Y(n346) );
endmodule

